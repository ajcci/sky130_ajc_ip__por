* NGSPICE file created from sky130_ajc_ip__por_rcx.ext - technology: sky130A

.subckt sky130_ajc_ip__por_rcx otrip[1] otrip[0] force_ena_rc_osc porb_h porb por
+ force_pdn ibg_200n dcomp startup_timed_out force_dis_rc_osc vbg_1v2 otrip[2] force_short_oneshot
+ itest vin osc_ck por_timed_out isrc_sel avdd avss pwup_filt dvdd dvss
X0 avdd.t207 por_ana_0.comparator_0.vpp.t14 por_ana_0.comparator_0.vpp.t15 avdd.t195 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1 por_ana_0.ibias_gen_0.vn0.t1 por_ana_0.ibias_gen_0.vp0.t12 avdd.t555 avdd.t554 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X2 dvdd.t101 a_39510_31251# por_dig_0._044_ dvdd.t100 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3 por_ana_0.comparator_1.n1.t1 por_ana_0.comparator_1.n0.t5 avdd.t545 avdd.t544 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.6
X4 a_34662_34363# por_dig_0.cnt_por\[6\] a_34580_34110# dvss.t462 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X5 a_38518_21903# a_38150_22885# dvss.t116 dvss.t115 sky130_fd_pr__nfet_01v8 ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X6 a_32980_33287# a_32464_32915# a_32885_33275# dvss.t472 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X7 dvss.t540 a_25863_32638# a_26288_32594# dvss.t539 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X8 a_29802_22973# a_29702_22885# dvss.t491 dvss.t490 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X9 porb.t31 por_ana_0.sky130_fd_sc_hd__inv_4_1.Y dvdd.t303 dvdd.t302 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 vbg_1v2.t1 dvss.t1679 dvss.t1681 dvss.t1680 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X11 dvss.t618 por_dig_0._009_ a_36331_33819# dvss.t617 sky130_fd_pr__nfet_01v8 ad=0.2205 pd=1.89 as=0.066 ps=0.745 w=0.42 l=0.15
X12 dvdd.t501 a_35583_34541# por_dig_0.clknet_1_1__leaf_osc_ck.t31 dvdd.t500 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X13 dvdd.t1524 dvss.t2234 dvdd.t1523 dvdd.t1522 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X14 dvdd.t499 a_35583_34541# por_dig_0.clknet_1_1__leaf_osc_ck.t30 dvdd.t498 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X15 a_34486_33703# por_dig_0.net22.t4 dvdd.t1238 dvdd.t1237 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.1725 ps=1.345 w=1 l=0.15
X16 dvdd.t369 por_dig_0.net24 a_35913_33819# dvdd.t368 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1092 ps=1.36 w=0.42 l=0.15
X17 por_ana_0.rstring_mux_0.vtrip_decoded_b_avdd[3] por_ana_0.rstring_mux_0.vtrip_decoded_avdd[3] avss.t9 avss.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X18 a_35468_30163# a_35293_30189# a_35647_30189# dvss.t383 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X19 a_32610_35603# por_dig_0._047_ dvss.t845 dvss.t844 sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.25675 ps=1.44 w=0.65 l=0.15
X20 por.t15 por_ana_0.sky130_fd_sc_hd__inv_4_4.Y dvss.t1167 dvss.t1166 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X21 dvdd.t978 por_ana_0.sky130_fd_sc_hd__inv_4_4.Y por.t31 dvdd.t977 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X22 a_35552_13935# a_35930_6535# avss.t26 sky130_fd_pr__res_xhigh_po_1p41 l=35
X23 dvdd.t1527 dvss.t2235 dvdd.t1526 dvdd.t1525 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X24 dvdd.t301 por_ana_0.sky130_fd_sc_hd__inv_4_1.Y porb.t30 dvdd.t300 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X25 a_8591_22912# a_8969_15512# avss.t27 sky130_fd_pr__res_xhigh_po_1p41 l=35
X26 dvdd.t69 a_36122_30341# por_dig_0.net29 dvdd.t68 sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.26 ps=2.52 w=1 l=0.15
X27 a_34387_32909# osc_ck.t8 dvss.t887 dvss.t886 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X28 por_ana_0.ibias_gen_0.vp0.t0 avdd.t175 avdd.t177 avdd.t176 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X29 dvdd.t1530 dvss.t2236 dvdd.t1529 dvdd.t1528 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X30 dvss.t1165 por_ana_0.sky130_fd_sc_hd__inv_4_4.Y por.t14 dvss.t1164 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X31 a_31016_13935# a_31394_6535# avss.t1 sky130_fd_pr__res_xhigh_po_1p41 l=35
X32 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[3] a_33121_24371# avdd.t557 avdd.t556 sky130_fd_pr__pfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.24375 ps=1.825 w=1.5 l=0.5
X33 dvdd.t1533 dvss.t2237 dvdd.t1532 dvdd.t1531 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X34 a_34762_36173# por_dig_0.net23.t4 dvdd.t755 dvdd.t754 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.1725 ps=1.345 w=1 l=0.15
X35 por_dig_0.net10 a_31651_30341# dvdd.t980 dvdd.t979 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X36 avdd.t402 por_ana_0.comparator_1.vpp.t47 por_ana_0.comparator_1.n0.t0 avdd.t401 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X37 dvss.t79 por_ana_0.sky130_fd_sc_hd__inv_4_3.Y dcomp.t15 dvss.t78 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X38 dvss.t616 a_33926_22885# a_34026_22973# dvss.t615 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X39 por_ana_0.rstring_mux_0.vtrip3.t4 por_ana_0.rstring_mux_0.vtrip2.t2 avss.t149 sky130_fd_pr__res_xhigh_po_1p41 l=35
X40 dvss.t1123 a_33172_28165# por_dig_0.net12 dvss.t523 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.221 ps=1.98 w=0.65 l=0.15
X41 a_35202_29877# a_35298_29619# dvss.t391 dvss.t390 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.5
X42 dvss.t1958 dvdd.t1810 dvss.t1957 dvss.t1956 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X43 dvss.t1955 dvdd.t1811 dvss.t1954 dvss.t1872 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X44 por_ana_0.rstring_mux_0.vtrip_decoded_b_avdd[6] por_ana_0.rstring_mux_0.vtrip_decoded_avdd[6].t2 avdd.t391 avdd.t390 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X45 dvss.t1133 a_23734_23637# a_24159_23593# dvss.t1132 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X46 por_dig_0._034_.t9 por_dig_0.cnt_por\[2\] dvdd.t1279 dvdd.t1278 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X47 a_34482_34541# por_dig_0.cnt_por\[2\] a_34398_34541# dvss.t1581 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X48 avdd.t379 por_ana_0.ibias_gen_0.vp.t7 por_ana_0.ibias_gen_0.ibias0.t1 avdd.t378 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X49 a_26288_32594# a_25863_32638# dvss.t538 dvss.t537 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X50 a_39417_31795# force_short_oneshot.t2 dvdd.t730 dvdd.t729 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X51 a_31651_30341# por_dig_0.net2 dvdd.t147 dvdd.t146 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14575 ps=1.335 w=0.42 l=0.15
X52 a_39887_21959# a_39887_23089# avdd.t273 avdd.t272 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.1197 ps=1.41 w=0.42 l=0.5
X53 a_33334_28557# por_dig_0.net7.t2 dvdd.t732 dvdd.t731 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14575 ps=1.335 w=1 l=0.15
X54 dcomp.t14 por_ana_0.sky130_fd_sc_hd__inv_4_3.Y dvss.t77 dvss.t76 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X55 avdd.t257 a_31914_22973# a_32607_21859# avdd.t256 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.1365 ps=1.49 w=0.42 l=1
X56 por_dig_0._032_ por_dig_0._031_ dvdd.t145 dvdd.t144 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X57 dvdd.t1536 dvss.t2238 dvdd.t1535 dvdd.t1534 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X58 dvdd.t943 por_dig_0._048_ por_dig_0._006_ dvdd.t942 sky130_fd_pr__pfet_01v8_hvt ad=0.182 pd=1.92 as=0.174 ps=1.39 w=0.7 l=0.15
X59 por_ana_0.rstring_mux_0.vtrip5.t0 por_ana_0.rstring_mux_0.vtrip6.t0 avss.t0 sky130_fd_pr__res_xhigh_po_1p41 l=35
X60 por_ana_0.schmitt_trigger_0.m.t7 por_ana_0.schmitt_trigger_0.in.t1 dvdd.t559 dvdd.t558 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X61 por_ana_0.comparator_1.vpp.t15 por_ana_0.comparator_1.vpp.t14 avdd.t400 avdd.t395 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X62 dvdd.t367 por_dig_0.net24 a_35092_33427# dvdd.t366 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X63 dvdd.t306 por_dig_0._028_ a_34746_29645# dvdd.t70 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X64 dvdd.t384 por_dig_0.cnt_por\[3\] por_dig_0._034_.t1 dvdd.t383 sky130_fd_pr__pfet_01v8_hvt ad=0.215 pd=1.43 as=0.135 ps=1.27 w=1 l=0.15
X65 por_ana_0.comparator_0.vnn.t13 por_ana_0.comparator_0.vpp.t47 avdd.t206 avdd.t182 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X66 dvdd.t1 por_dig_0.cnt_rsb a_34510_31277# dvdd.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X67 dvss.t1953 dvdd.t1812 dvss.t1952 dvss.t1951 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X68 por_ana_0.comparator_0.vinn.t18 avss.t134 por_ana_0.comparator_0.vinn.t18 avss.t135 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=0.6
X69 a_36138_22973# a_36038_22885# dvss.t282 dvss.t281 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X70 por_dig_0._022_ por_dig_0.cnt_por\[6\] a_34212_33997# dvdd.t393 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X71 a_37961_33453# a_37046_33453# a_37614_33695# dvss.t19 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X72 por_dig_0.cnt_por\[0\].t3 a_36756_35603# dvss.t564 dvss.t563 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X73 a_39881_33703# por_dig_0.cnt_st\[1\] dvdd.t511 dvdd.t510 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.14575 ps=1.335 w=0.42 l=0.15
X74 dvdd.t322 por_dig_0.net32 a_34594_32615# dvdd.t321 sky130_fd_pr__pfet_01v8_hvt ad=0.365 pd=1.73 as=0.105 ps=1.21 w=1 l=0.15
X75 por_dig_0._018_ por_dig_0.cnt_por\[4\] dvss.t1552 dvss.t1551 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X76 dvdd.t749 por_dig_0._034_.t10 a_35942_31821# dvdd.t748 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X77 dvss.t832 a_38320_34301# a_38254_34375# dvss.t831 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X78 a_32019_33819# a_31893_33721# a_31615_33705# dvss.t477 sky130_fd_pr__special_nfet_01v8 ad=0.0999 pd=0.985 as=0.0711 ps=0.755 w=0.36 l=0.15
X79 dvss.t75 por_ana_0.sky130_fd_sc_hd__inv_4_3.Y dcomp.t13 dvss.t74 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X80 avdd.t205 por_ana_0.comparator_0.vpp.t48 por_ana_0.comparator_0.vnn.t12 avdd.t180 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X81 a_3299_22912# a_2921_15512# avss.t27 sky130_fd_pr__res_xhigh_po_1p41 l=35
X82 a_24159_23593# a_23734_23637# dvss.t1131 dvss.t1130 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X83 avss.t133 avss.t132 avss.t133 avss.t68 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=8
X84 pwup_filt.t31 por_ana_0.sky130_fd_sc_hd__inv_4_0.Y dvdd.t225 dvdd.t224 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X85 a_31526_31827# a_31360_31827# dvss.t33 dvss.t32 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X86 avss.t131 avss.t129 avss.t130 avss.t81 sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0 ps=0 w=5 l=8
X87 a_34746_31277# a_34510_31277# dvss.t464 dvss.t463 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.5
X88 dvss.t226 por_ana_0.sky130_fd_sc_hd__inv_4_1.A por_ana_0.sky130_fd_sc_hd__inv_4_1.Y dvss.t225 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X89 avss.t144 por_ana_0.sky130_fd_sc_hvl__inv_4_0.A por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.t7 avss.t143 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.105 ps=1.03 w=0.75 l=0.5
X90 a_32233_33819# a_32019_33819# dvdd.t1281 dvdd.t1280 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07035 ps=0.755 w=0.42 l=0.15
X91 por_dig_0.net7.t1 a_34615_28013# dvdd.t937 dvdd.t936 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X92 dvss.t5 a_32701_28531# por_dig_0.otrip_decoded[1] dvss.t4 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X93 dvdd.t413 por_dig_0.clknet_1_0__leaf_osc_ck.t32 a_36972_30189# dvdd.t412 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X94 por_ana_0.schmitt_trigger_0.m.t8 por_ana_0.schmitt_trigger_0.out.t4 dvdd.t702 dvdd.t701 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X95 dvdd.t684 por_dig_0.por_unbuf.t4 por_ana_0.sky130_fd_sc_hd__inv_4_1.A dvdd.t683 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X96 a_35640_32517# por_dig_0.net23.t5 dvdd.t757 dvdd.t756 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.142225 ps=1.335 w=0.42 l=0.15
X97 dvdd.t223 por_ana_0.sky130_fd_sc_hd__inv_4_0.Y pwup_filt.t30 dvdd.t222 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X98 dvdd.t1240 por_dig_0.net22.t5 a_33600_34335# dvdd.t1239 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X99 dvss.t1532 por_dig_0.cnt_st\[4\] a_37616_32141# dvss.t1531 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X100 dvss.t2143 isrc_sel.t2 a_38150_24619# dvss.t2142 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X101 a_32088_31514# a_31893_31545# a_32398_31277# dvss.t21 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.1401 ps=1.1 w=0.36 l=0.15
X102 por_dig_0.clknet_1_1__leaf_osc_ck.t15 a_35583_34541# dvss.t596 dvss.t595 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X103 a_35645_31277# por_dig_0._015_ dvss.t378 dvss.t377 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X104 dvss.t280 a_36038_22885# a_36138_22973# dvss.t279 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X105 por_dig_0.net4 a_39417_31795# dvdd.t456 dvdd.t455 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X106 avdd.t174 avdd.t172 avdd.t173 avdd.t3 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=8
X107 por_ana_0.comparator_0.vinn.t6 avdd.t170 por_ana_0.comparator_0.vinn.t6 avdd.t171 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=0.6
X108 dvdd.t33 por_dig_0._033_ a_35640_32517# dvdd.t32 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.06615 ps=0.735 w=0.42 l=0.15
X109 dvss.t1950 dvdd.t1813 dvss.t1949 dvss.t1948 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X110 a_8591_22912# a_8213_15512# avss.t27 sky130_fd_pr__res_xhigh_po_1p41 l=35
X111 dvdd.t97 a_38053_30189# a_38228_30163# dvdd.t96 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X112 a_32088_31514# a_31932_31419# a_32233_31643# dvdd.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.1155 ps=0.97 w=0.42 l=0.15
X113 a_33161_36539# por_dig_0._007_ dvdd.t7 dvdd.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X114 avdd.t249 por_ana_0.rstring_mux_0.ena_b por_ana_0.rstring_mux_0.vtop.t15 avdd.t248 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X115 dvss.t323 a_39162_33453# a_39268_33453# dvss.t322 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.5
X116 a_5567_22912# a_5189_15512# avss.t27 sky130_fd_pr__res_xhigh_po_1p41 l=35
X117 dvss.t368 a_25846_23637# a_26271_23593# dvss.t367 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X118 dvdd.t399 a_32616_32125# a_32603_31821# dvdd.t398 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X119 por_dig_0.clknet_1_0__leaf_osc_ck.t15 a_34098_30707# dvss.t210 dvss.t209 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X120 a_34098_30707# por_dig_0.clknet_0_osc_ck.t32 dvss.t2127 dvss.t2126 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X121 dvss.t1947 dvdd.t1814 dvss.t1946 dvss.t1860 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X122 a_35030_28557# por_dig_0.net5.t2 dvss.t2112 dvss.t2111 sky130_fd_pr__nfet_01v8 ad=0.10785 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X123 avss.t128 avss.t126 avss.t127 avss.t64 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=8
X124 a_34734_34363# por_dig_0.net22.t6 a_34662_34363# dvss.t1525 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X125 por_dig_0.cnt_por\[2\] a_33996_36477# dvss.t1571 dvss.t1570 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X126 a_33012_33997# por_dig_0._047_ a_32794_33971# dvdd.t728 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.26 ps=2.52 w=1 l=0.15
X127 a_32607_23593# a_32182_23637# dvss.t15 dvss.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X128 a_33804_31251# por_dig_0.cnt_por\[8\] dvdd.t267 dvdd.t266 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.175 ps=1.35 w=1 l=0.15
X129 dvss.t1163 por_ana_0.sky130_fd_sc_hd__inv_4_4.Y por.t13 dvss.t1162 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X130 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.t6 por_ana_0.sky130_fd_sc_hvl__inv_4_0.A avss.t142 avss.t141 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X131 a_38250_22973# a_38150_22885# dvss.t114 dvss.t113 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X132 por_ana_0.rstring_mux_0.vtrip2.t1 por_ana_0.rstring_mux_0.otrip_decoded_avdd[2] vin.t1 avss.t5 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X133 por_ana_0.comparator_0.vinn.t17 avss.t124 por_ana_0.comparator_0.vinn.t17 avss.t125 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=0.6
X134 dvdd.t245 por_ana_0.rc_osc_0.in por_ana_0.rc_osc_0.m dvdd.t244 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X135 a_32607_21859# a_32182_21903# dvss.t1122 dvss.t1121 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X136 por_ana_0.rstring_mux_0.vtop.t14 por_ana_0.rstring_mux_0.ena_b avdd.t247 avdd.t246 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=0.6
X137 a_33930_36551# a_32740_36179# a_33821_36551# dvss.t448 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X138 a_37488_30189# a_36972_30189# a_37393_30189# dvss.t29 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X139 por_ana_0.ibias_gen_0.vstart.t9 vbg_1v2.t2 por_ana_0.ibias_gen_0.vn0.t6 avss.t150 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X140 dvdd.t253 por_dig_0._042_ a_37528_31527# dvdd.t252 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X141 a_34102_29965# por_dig_0.net30 dvss.t375 dvss.t374 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X142 dvss.t837 a_31413_32339# por_timed_out.t1 dvss.t836 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X143 a_7835_22912# a_7457_15512# avss.t27 sky130_fd_pr__res_xhigh_po_1p41 l=35
X144 por_ana_0.rstring_mux_0.otrip_decoded_b_avdd[1] por_ana_0.rstring_mux_0.otrip_decoded_avdd[1] avss.t33 avss.t32 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X145 a_33161_36539# por_dig_0._007_ dvss.t17 dvss.t16 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X146 dvdd.t1096 otrip[2].t2 a_34615_28013# dvdd.t1095 sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X147 a_33444_31037# por_dig_0.net24 dvdd.t365 dvdd.t364 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X148 por_dig_0.clknet_0_osc_ck.t15 a_34387_32909# dvss.t165 dvss.t164 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X149 a_19676_13935# a_20054_6535# avss.t136 sky130_fd_pr__res_xhigh_po_1p41 l=35
X150 por_ana_0.comparator_1.vnn.t15 por_ana_0.comparator_1.vnn.t14 avdd.t632 avdd.t403 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X151 a_35666_35629# a_35500_35629# dvdd.t442 dvdd.t441 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X152 a_38136_33427# a_37961_33453# a_38315_33453# dvss.t621 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X153 por_ana_0.sky130_fd_sc_hd__inv_4_4.Y por_dig_0.por_unbuf.t5 dvdd.t686 dvdd.t685 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X154 dvdd.t1294 dvdd.t1292 dvdd.t1294 dvdd.t1293 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.18
X155 dvss.t1945 dvdd.t1815 dvss.t1944 dvss.t1740 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X156 dvss.t604 a_33162_35603# por_dig_0._008_ dvss.t603 sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X157 por_ana_0.comparator_1.vt.t53 vbg_1v2.t3 por_ana_0.comparator_1.vnn por_ana_0.comparator_1.vt.t41 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X158 avdd.t478 por_ana_0.comparator_0.n1.t4 por_ana_0.dcomp3v3uv avdd.t477 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X159 avdd.t323 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.t8 porb_h.t15 avdd.t322 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X160 dvss.t1943 dvdd.t1816 dvss.t1942 dvss.t1941 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X161 a_36382_31795# por_dig_0._037_ a_36669_31821# dvdd.t99 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.21 ps=1.42 w=1 l=0.15
X162 dvdd.t688 por_dig_0.por_unbuf.t6 por_ana_0.sky130_fd_sc_hd__inv_4_4.Y dvdd.t687 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X163 dvdd.t1249 por_dig_0.otrip_decoded[4] a_25478_22885# dvdd.t1248 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X164 a_29802_24707# a_29702_24619# dvss.t1546 dvss.t1545 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X165 dvdd.t497 a_35583_34541# por_dig_0.clknet_1_1__leaf_osc_ck.t29 dvdd.t496 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X166 a_34842_32365# por_dig_0.net32 dvss.t387 dvss.t386 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X167 dvdd.t299 por_ana_0.sky130_fd_sc_hd__inv_4_1.Y porb.t29 dvdd.t298 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X168 dvdd.t1539 dvss.t2239 dvdd.t1538 dvdd.t1537 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X169 a_16652_13935# a_17030_6535# avss.t319 sky130_fd_pr__res_xhigh_po_1p41 l=35
X170 dvdd.t1437 por_dig_0.otrip_decoded[5].t4 a_25478_24619# dvdd.t1436 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X171 a_37952_31037# a_37777_31111# a_38131_31099# dvss.t1472 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X172 a_35612_33595# por_dig_0.clknet_1_1__leaf_osc_ck.t32 dvss.t699 dvss.t698 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X173 a_25863_32638# a_25495_33620# dvss.t1467 dvss.t1466 sky130_fd_pr__nfet_01v8 ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X174 dvss.t1161 por_ana_0.sky130_fd_sc_hd__inv_4_4.Y por.t12 dvss.t1160 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X175 por_ana_0.rstring_mux_0.vtrip2.t7 por_ana_0.rstring_mux_0.otrip_decoded_b_avdd[2] vin.t37 avdd.t527 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X176 por_ana_0.comparator_0.vinn.t5 avdd.t168 por_ana_0.comparator_0.vinn.t5 avdd.t169 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=0.6
X177 por_ana_0.rc_osc_0.m por_ana_0.rc_osc_0.in dvss.t296 dvss.t295 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.1475 ps=1.295 w=1 l=0.5
X178 dvss.t787 a_27958_23637# a_28383_23593# dvss.t786 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X179 a_35776_28013# por_dig_0.net6 dvdd.t682 dvdd.t681 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X180 a_33161_35451# por_dig_0._008_ dvss.t389 dvss.t388 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X181 por_dig_0.otrip_decoded[3].t1 a_37800_28013# dvss.t1487 dvss.t523 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X182 por_ana_0.comparator_0.vpp.t16 vbg_1v2.t4 por_ana_0.comparator_0.vt.t53 por_ana_0.comparator_0.vt.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X183 por_dig_0.net8 a_32004_30189# dvdd.t1172 dvdd.t1171 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X184 vin.t21 avss.t122 vin.t21 avss.t123 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=0.6
X185 dvss.t516 a_33926_24619# a_34026_24707# dvss.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X186 a_37046_32915# a_36880_32915# dvdd.t434 dvdd.t433 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X187 a_35394_28013# a_35217_28013# dvss.t524 dvss.t523 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X188 a_39718_33605# por_dig_0.cnt_st\[0\] a_39881_33703# dvdd.t1117 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X189 dcomp.t12 por_ana_0.sky130_fd_sc_hd__inv_4_3.Y dvss.t73 dvss.t72 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X190 a_34719_23593# a_34294_23637# dvss.t1349 dvss.t1348 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X191 a_34824_30189# a_34378_30189# a_34728_30189# dvss.t1351 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X192 a_39328_34515# por_dig_0.cnt_st\[0\] dvdd.t1116 dvdd.t1115 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X193 a_34486_33703# por_dig_0.cnt_por\[4\] dvdd.t1260 dvdd.t1259 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X194 a_33983_36173# a_32906_36179# a_33821_36551# dvdd.t615 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X195 por_ana_0.rc_osc_0.in dvss.t294 sky130_fd_pr__cap_mim_m3_2 l=30 w=30
X196 dvss.t1940 dvdd.t1817 dvss.t1939 dvss.t1938 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X197 por_dig_0.net17 a_35130_28673# dvdd.t617 dvdd.t616 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X198 por_dig_0._009_ por_dig_0._048_ dvdd.t941 dvdd.t940 sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.39 as=0.182 ps=1.92 w=0.7 l=0.15
X199 avss.t314 a_2165_15512# avss.t27 sky130_fd_pr__res_xhigh_po_1p41 l=35
X200 a_34719_21859# a_34294_21903# dvss.t1497 dvss.t1496 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X201 por_dig_0.otrip_decoded[6].t1 a_35960_29101# dvss.t1501 dvss.t1500 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X202 a_34398_34541# por_dig_0.cnt_por\[0\].t8 a_34302_34541# dvss.t636 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X203 dvdd.t1222 por_dig_0._011_ a_32651_33819# dvdd.t1221 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X204 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[1] a_31009_24371# dvss.t1504 dvss.t517 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.121875 ps=1.075 w=0.75 l=0.5
X205 por_dig_0.cnt_por\[10\] a_36480_31251# dvdd.t1226 dvdd.t1225 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X206 dvss.t71 por_ana_0.sky130_fd_sc_hd__inv_4_3.Y dcomp.t11 dvss.t70 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X207 avdd.t204 por_ana_0.comparator_0.vpp.t49 por_ana_0.comparator_0.vnn.t11 avdd.t180 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X208 a_23734_23637# a_23366_24619# dvss.t1524 dvss.t1523 sky130_fd_pr__nfet_01v8 ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X209 a_36262_32365# por_dig_0._033_ dvss.t39 dvss.t38 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.13165 ps=1.14 w=0.42 l=0.15
X210 a_34570_32141# por_dig_0.cnt_por\[6\] dvss.t461 dvss.t460 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X211 a_21944_13935# a_21566_6535# avss.t306 sky130_fd_pr__res_xhigh_po_1p41 l=35
X212 a_34202_36717# por_dig_0._033_ por_dig_0._016_ dvss.t37 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X213 por_ana_0.comparator_0.vt.t35 avss.t410 por_ana_0.comparator_0.vnn.t22 por_ana_0.comparator_0.vt.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=8
X214 avss.t400 por_ana_0.ibias_gen_0.vn1.t10 por_ana_0.ibias_gen_0.vp1.t9 avss.t396 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=8
X215 vin.t34 por_ana_0.rstring_mux_0.otrip_decoded_avdd[0] por_ana_0.rstring_mux_0.vtrip0.t9 avss.t310 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X216 a_34762_36173# por_dig_0.cnt_por\[1\] dvdd.t1170 dvdd.t1169 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X217 a_34746_29645# por_dig_0.net29 dvdd.t183 dvdd.t70 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X218 a_24159_21859# a_23734_21903# dvss.t1415 dvss.t1414 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X219 a_36138_24707# a_36038_24619# dvss.t685 dvss.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X220 dvdd.t579 a_37798_33971# a_37688_33997# dvdd.t578 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X221 a_36564_32339# por_dig_0.net20.t2 dvss.t2102 dvss.t2101 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.06825 ps=0.745 w=0.42 l=0.15
X222 por_ana_0.ibias_gen_0.vp1.t8 por_ana_0.ibias_gen_0.vn1.t11 avss.t401 avss.t398 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=8
X223 dvss.t1678 dvss.t1676 por_ana_0.rc_osc_0.m dvss.t1677 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X224 por_dig_0.cnt_por\[8\] a_33444_31037# dvdd.t316 dvdd.t315 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X225 dvdd.t415 por_dig_0.clknet_1_0__leaf_osc_ck.t33 a_31728_32365# dvdd.t414 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X226 por_dig_0.net3 a_31360_28557# dvdd.t589 dvdd.t588 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X227 dvss.t869 por_dig_0.net23.t6 a_36500_33229# dvss.t868 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.095875 ps=0.945 w=0.65 l=0.15
X228 a_32244_32365# a_31728_32365# a_32149_32365# dvss.t695 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X229 dvss.t1361 a_34265_27987# por_dig_0.otrip_decoded[4] dvss.t523 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X230 a_4055_22912# a_4433_15512# avss.t27 sky130_fd_pr__res_xhigh_po_1p41 l=35
X231 avdd.t167 avdd.t165 avdd.t166 avdd.t3 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=8
X232 a_37961_33287# a_37046_32915# a_37614_32883# dvss.t19 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X233 dvss.t1937 dvdd.t1818 dvss.t1936 dvss.t1853 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X234 por_ana_0.comparator_0.vinn.t46 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[7].t2 por_ana_0.rstring_mux_0.vtrip7.t5 avss.t392 sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=0.6
X235 dvss.t562 a_36756_35603# por_dig_0.cnt_por\[0\].t2 dvss.t561 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X236 vin.t9 avdd.t163 vin.t9 avdd.t164 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=0.6
X237 dvdd.t1435 por_dig_0.otrip_decoded[6].t4 a_27590_22885# dvdd.t1434 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X238 dvdd.t452 a_35468_30163# a_35455_30555# dvdd.t451 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X239 a_18920_13935# a_18542_6535# avss.t304 sky130_fd_pr__res_xhigh_po_1p41 l=35
X240 dvss.t1347 a_34294_23637# a_34719_23593# dvss.t1346 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X241 dvdd.t1420 por_dig_0.otrip_decoded[7].t4 a_27590_24619# dvdd.t1419 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X242 dvdd.t1418 otrip[1].t2 a_33971_28557# dvdd.t1417 sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X243 por_ana_0.comparator_1.vnn.t13 por_ana_0.comparator_1.vnn.t12 avdd.t631 avdd.t403 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X244 dvdd.t1542 dvss.t2240 dvdd.t1541 dvdd.t1540 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X245 por_dig_0._045_ a_37789_31821# dvss.t1389 dvss.t1388 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X246 dvss.t208 a_34098_30707# por_dig_0.clknet_1_0__leaf_osc_ck.t14 dvss.t207 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X247 a_33198_32883# a_32980_33287# dvss.t627 dvss.t626 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X248 avss.t390 por_ana_0.comparator_0.vn.t7 por_ana_0.comparator_0.vt.t54 avss.t45 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X249 a_14384_13935# a_14006_6535# avss.t305 sky130_fd_pr__res_xhigh_po_1p41 l=35
X250 a_35699_33819# a_35612_33595# a_35295_33705# dvdd.t1209 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.0588 ps=0.7 w=0.42 l=0.15
X251 a_33450_33453# por_dig_0.cnt_por\[6\] a_33366_33453# dvss.t459 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X252 dvdd.t704 por_ana_0.schmitt_trigger_0.out.t5 por_ana_0.schmitt_trigger_0.m.t9 dvdd.t703 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X253 dvdd.t809 a_35958_31519# a_35848_31643# dvdd.t808 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X254 por_dig_0._022_ por_dig_0.net22.t7 a_34295_34317# dvss.t1526 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.095875 ps=0.945 w=0.65 l=0.15
X255 por_dig_0._042_ por_dig_0.cnt_st\[3\] a_38622_31053# dvss.t934 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X256 a_32704_31111# a_32188_30739# a_32609_31099# dvss.t938 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X257 a_36016_35629# a_35666_35629# a_35921_35629# dvdd.t519 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X258 por_ana_0.rc_osc_0.ena_b por_dig_0.osc_ena.t4 dvdd.t1422 dvdd.t1421 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X259 a_32818_28013# a_32641_28013# dvss.t943 dvss.t523 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X260 por_ana_0.comparator_1.vpp.t31 vin.t50 por_ana_0.comparator_1.vt.t35 por_ana_0.comparator_1.vt.t18 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X261 por_ana_0.comparator_0.vt.t55 por_ana_0.comparator_0.vn.t8 avss.t391 avss.t45 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X262 a_37952_31037# por_dig_0.net25 dvdd.t848 dvdd.t847 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X263 por_ana_0.comparator_1.vpp.t17 por_ana_0.comparator_1.vnn.t47 avdd.t633 avdd.t395 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X264 avdd.t162 avdd.t160 avdd.t162 avdd.t161 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=4
X265 a_35666_35629# a_35500_35629# dvss.t528 dvss.t527 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X266 a_33600_34335# por_dig_0.net4 dvdd.t89 dvdd.t88 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X267 a_6323_22912# a_6701_15512# avss.t27 sky130_fd_pr__res_xhigh_po_1p41 l=35
X268 por_ana_0.comparator_0.vinn.t16 avss.t120 por_ana_0.comparator_0.vinn.t16 avss.t121 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=0.6
X269 vin.t23 por_ana_0.rstring_mux_0.otrip_decoded_b_avdd[0] por_ana_0.rstring_mux_0.vtrip0.t6 avdd.t430 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X270 dvss.t684 a_36038_24619# a_36138_24707# dvss.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X271 dvdd.t852 a_33752_28013# por_dig_0.otrip_decoded[2].t3 dvdd.t851 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X272 dvss.t969 a_38974_34693# por_dig_0.net31 dvss.t968 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X273 dvss.t800 por_dig_0.net6 a_34290_28557# dvss.t799 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X274 a_36831_23593# a_36406_23637# dvss.t982 dvss.t981 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X275 a_38136_33427# por_dig_0.net25 dvdd.t846 dvdd.t845 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X276 a_38228_30163# por_dig_0.net25 dvdd.t844 dvdd.t843 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X277 a_29802_22973# a_29702_22885# dvss.t489 dvss.t488 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X278 por_dig_0.clknet_1_0__leaf_osc_ck.t13 a_34098_30707# dvss.t206 dvss.t205 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X279 a_32630_32915# a_32464_32915# dvss.t471 dvss.t470 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X280 dvdd.t1545 dvss.t2241 dvdd.t1544 dvdd.t1543 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X281 a_37064_13935# a_36686_6535# avss.t225 sky130_fd_pr__res_xhigh_po_1p41 l=35
X282 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[3] a_33121_24371# dvss.t1567 dvss.t517 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.121875 ps=1.075 w=0.75 l=0.5
X283 por_ana_0.comparator_0.vinn.t27 por_ana_0.rstring_mux_0.vtrip_decoded_b_avdd[7] por_ana_0.rstring_mux_0.vtrip7.t1 avdd.t434 sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=0.6
X284 por_ana_0.rstring_mux_0.vtrip7.t3 por_ana_0.rstring_mux_0.otrip_decoded_avdd[7] vin.t25 avss.t229 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X285 dvss.t635 pwup_filt.t32 a_32004_30189# dvss.t634 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X286 dvdd.t1548 dvss.t2242 dvdd.t1547 dvdd.t1546 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X287 a_25846_23637# a_25478_24619# dvss.t1484 dvss.t1483 sky130_fd_pr__nfet_01v8 ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X288 avdd.t159 avdd.t158 avdd.t159 avdd.t33 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=8
X289 dvdd.t87 por_dig_0.net4 a_35040_34587# dvdd.t86 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.1092 ps=1.36 w=0.42 l=0.15
X290 avdd.t604 por_ana_0.rstring_mux_0.ena.t1 por_ana_0.ibias_gen_0.vp1.t17 avdd.t603 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X291 por_ana_0.rc_osc_0.m por_ana_0.rc_osc_0.n.t6 dvss.t2020 dvss.t2019 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X292 dvss.t987 a_38146_31429# por_dig_0.net34 dvss.t986 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X293 a_36494_35091# a_36328_35091# dvss.t994 dvss.t993 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X294 a_26271_21859# a_25846_21903# dvss.t1006 dvss.t1005 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X295 dvss.t1935 dvdd.t1819 dvss.t1934 dvss.t1682 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X296 por.t11 por_ana_0.sky130_fd_sc_hd__inv_4_4.Y dvss.t1159 dvss.t1158 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X297 avdd.t362 por_ana_0.comparator_0.vnn.t47 por_ana_0.comparator_0.vm.t5 avdd.t195 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X298 por_dig_0._050_ a_35592_36286# dvdd.t876 dvdd.t875 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X299 a_38250_24707# a_38150_24619# dvss.t47 dvss.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X300 por_ana_0.comparator_1.vpp.t18 por_ana_0.comparator_1.vnn.t48 avdd.t634 avdd.t395 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X301 dvdd.t883 a_37584_35389# a_37571_35085# dvdd.t882 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X302 por_dig_0.net22.t3 a_36380_33971# dvdd.t887 dvdd.t886 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X303 avss.t345 por_ana_0.comparator_1.vm.t4 por_ana_0.comparator_1.vm.t5 avss.t290 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X304 porb_h.t31 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.t9 avss.t179 avss.t178 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X305 a_36100_32517# por_dig_0._033_ dvdd.t31 dvdd.t30 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.142225 ps=1.335 w=0.42 l=0.15
X306 por_dig_0._020_ por_dig_0.net22.t8 a_33378_34317# dvss.t1169 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X307 a_37658_33275# a_37614_32883# a_37492_33287# dvss.t356 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X308 dvss.t2150 a_36381_36691# por_dig_0.por_unbuf.t1 dvss.t2149 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X309 dvdd.t1477 por_dig_0.net13 a_33752_28013# dvdd.t1476 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X310 dvdd.t862 a_35040_34587# por_dig_0._046_ dvdd.t861 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X311 dvdd.t1550 dvss.t2243 a_29702_22885# dvdd.t1549 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X312 por_dig_0.net1 a_31360_33997# dvss.t2154 dvss.t2153 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X313 dvss.t395 a_35092_33427# por_dig_0.cnt_por\[4\] dvss.t394 sky130_fd_pr__nfet_01v8 ad=0.2087 pd=2.02 as=0.169 ps=1.82 w=0.65 l=0.15
X314 por_dig_0.clknet_0_osc_ck.t14 a_34387_32909# dvss.t163 dvss.t162 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X315 por_ana_0.comparator_0.vinn.t4 avdd.t156 por_ana_0.comparator_0.vinn.t4 avdd.t157 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=0.6
X316 por_ana_0.comparator_0.vn.t5 por_ana_0.comparator_0.ena_b.t2 avss.t332 avss.t331 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X317 dvss.t980 a_36406_23637# a_36831_23593# dvss.t979 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X318 dvdd.t1258 por_dig_0.cnt_por\[4\] a_36100_32517# dvdd.t1257 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.06615 ps=0.735 w=0.42 l=0.15
X319 por_ana_0.dcomp3v3uv por_ana_0.comparator_0.n1.t5 avdd.t480 avdd.t479 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X320 por_ana_0.comparator_0.vt.t17 por_ana_0.comparator_0.vinn.t48 por_ana_0.comparator_0.vnn por_ana_0.comparator_0.vt.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X321 dvss.t2168 a_31814_22885# a_31914_22973# dvss.t2167 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X322 dvss.t2170 a_33852_29645# por_dig_0._014_ dvss.t2169 sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.25025 ps=1.42 w=0.65 l=0.15
X323 a_33934_32615# por_dig_0._019_ dvdd.t1496 dvdd.t1495 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.1725 ps=1.345 w=1 l=0.15
X324 avdd.t580 por_ana_0.ibias_gen_0.isrc_sel.t2 por_ana_0.ibias_gen_0.isrc_sel_b.t2 avdd.t579 sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=1
X325 por_ana_0.ibias_gen_0.vstart.t8 vbg_1v2.t5 por_ana_0.ibias_gen_0.vn0.t7 avss.t150 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X326 dvdd.t1552 dvss.t2244 a_29702_24619# dvdd.t1551 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X327 a_35227_32141# por_dig_0.cnt_por\[9\] a_35000_31795# dvss.t2186 sky130_fd_pr__nfet_01v8 ad=0.118625 pd=1.015 as=0.19825 ps=1.91 w=0.65 l=0.15
X328 a_39510_31251# por_dig_0._030_ dvss.t2192 dvss.t2191 sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.25675 ps=1.44 w=0.65 l=0.15
X329 avdd.t285 a_29802_22973# a_31009_22637# avdd.t284 sky130_fd_pr__pfet_g5v0d10v5 ad=0.24375 pd=1.825 as=0.3975 ps=3.53 w=1.5 l=0.5
X330 por_ana_0.rstring_mux_0.otrip_decoded_avdd[2] a_24673_22637# dvss.t2196 dvss.t2195 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.121875 ps=1.075 w=0.75 l=0.5
X331 dvss.t2206 a_27958_21903# a_28383_21859# dvss.t2205 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X332 a_36382_31795# por_dig_0.cnt_st\[4\] dvdd.t1247 dvdd.t1225 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.15 ps=1.3 w=1 l=0.15
X333 dvss.t1933 dvdd.t1820 dvss.t1932 dvss.t1931 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X334 avdd.t582 por_ana_0.ibias_gen_0.isrc_sel.t3 a_12598_23626# avdd.t581 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X335 por_ana_0.rstring_mux_0.vtrip7.t9 por_ana_0.rstring_mux_0.otrip_decoded_b_avdd[7] vin.t49 avdd.t654 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X336 a_19094_2382# a_41694_2004# dvss.t2207 sky130_fd_pr__res_xhigh_po_1p41 l=111
X337 avdd.t155 avdd.t153 avdd.t154 avdd.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=8
X338 dvdd.t1508 a_36581_35629# a_36756_35603# dvdd.t1507 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X339 a_32094_31795# a_31876_32199# dvss.t2210 dvss.t2209 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X340 dvdd.t133 a_34387_32909# por_dig_0.clknet_0_osc_ck.t31 dvdd.t132 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X341 a_32535_28013# a_32358_28013# dvss.t2212 dvss.t523 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X342 a_17398_35244# a_17020_27844# avss.t408 sky130_fd_pr__res_xhigh_po_1p41 l=35
X343 a_39554_33997# por_dig_0.net4 dvdd.t85 dvdd.t84 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X344 dvss.t385 por_dig_0.net32 a_34486_32365# dvss.t384 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X345 dvdd.t1291 dvdd.t1289 por_ana_0.schmitt_trigger_0.m.t13 dvdd.t1290 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X346 dvss.t1930 dvdd.t1821 dvss.t1929 dvss.t1720 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X347 a_36334_32365# por_dig_0.cnt_por\[4\] a_36262_32365# dvss.t1550 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X348 a_38943_23593# a_38518_23637# dvss.t2223 dvss.t2222 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X349 a_25595_33708# a_25495_33620# dvss.t1465 dvss.t1464 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X350 por_dig_0.cnt_st\[4\] a_37952_31037# dvdd.t1203 dvdd.t1202 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X351 dvss.t493 por_dig_0.clknet_1_0__leaf_osc_ck.t34 a_31728_32365# dvss.t492 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X352 dvss.t2151 por_dig_0.net13 a_33752_28013# dvss.t677 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X353 a_31413_29075# por_dig_0.net9 dvdd.t1517 dvdd.t618 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X354 dvss.t1928 dvdd.t1822 dvss.t1927 dvss.t1926 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X355 a_38576_13935# a_38954_6535# avss.t409 sky130_fd_pr__res_xhigh_po_1p41 l=35
X356 a_31914_22973# a_31814_22885# dvss.t2166 dvss.t2165 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X357 porb_h.t30 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.t10 avss.t181 avss.t180 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X358 dvdd.t734 por_dig_0.net7.t3 a_35776_28013# dvdd.t733 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X359 a_32354_30739# a_32188_30739# dvss.t937 dvss.t936 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X360 a_21178_35244# a_20800_27844# avss.t251 sky130_fd_pr__res_xhigh_po_1p41 l=35
X361 por_ana_0.ibias_gen_0.vn1.t5 por_ana_0.ibias_gen_0.vn1.t4 avss.t399 avss.t398 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=8
X362 por_ana_0.comparator_1.vpp.t19 por_ana_0.comparator_1.vnn.t49 avdd.t635 avdd.t395 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X363 a_27958_23637# a_27590_24619# dvss.t1385 dvss.t1384 sky130_fd_pr__nfet_01v8 ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X364 por_ana_0.comparator_1.ena_b por_ana_0.rstring_mux_0.ena.t2 avss.t381 avss.t380 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X365 a_33256_35463# a_32740_35091# a_33161_35451# dvss.t1222 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X366 a_22047_23593# a_21622_23637# dvss.t1234 dvss.t1233 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X367 a_19666_35244# a_19288_27844# avss.t258 sky130_fd_pr__res_xhigh_po_1p41 l=35
X368 a_28383_21859# a_27958_21903# dvss.t2204 dvss.t2203 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X369 a_32984_32339# por_dig_0.net24 dvdd.t363 dvdd.t362 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X370 dvss.t2014 por_dig_0._036_.t3 a_33374_31277# dvss.t2013 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X371 por_dig_0.net24 a_35100_32339# dvss.t1246 dvss.t1245 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X372 dvss.t1925 dvdd.t1823 dvss.t1924 dvss.t1825 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X373 a_38136_33213# por_dig_0.net24 dvdd.t361 dvdd.t360 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X374 dcomp.t31 por_ana_0.sky130_fd_sc_hd__inv_4_3.Y dvdd.t67 dvdd.t66 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X375 dvss.t1250 a_37751_31251# a_37392_31251# dvss.t1249 sky130_fd_pr__nfet_01v8 ad=0.1359 pd=1.1 as=0.08775 ps=0.92 w=0.65 l=0.15
X376 avdd.t152 avdd.t151 avdd.t152 avdd.t33 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=8
X377 por_ana_0.comparator_0.vt.t16 por_ana_0.comparator_0.vinn.t49 por_ana_0.comparator_0.vnn por_ana_0.comparator_0.vt.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X378 dvss.t1923 dvdd.t1824 dvss.t1922 dvss.t1921 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X379 a_31413_29075# por_dig_0.net9 dvss.t2227 dvss.t2226 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X380 pwup_filt.t29 por_ana_0.sky130_fd_sc_hd__inv_4_0.Y dvdd.t221 dvdd.t220 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X381 dvss.t1920 dvdd.t1825 dvss.t1919 dvss.t1918 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X382 avdd.t255 a_31914_22973# a_33121_22637# avdd.t254 sky130_fd_pr__pfet_g5v0d10v5 ad=0.24375 pd=1.825 as=0.3975 ps=3.53 w=1.5 l=0.5
X383 dvdd.t814 por_dig_0.cnt_st\[3\] a_38956_32339# dvdd.t813 sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0588 ps=0.7 w=0.42 l=0.15
X384 por_ana_0.comparator_1.vpp.t20 por_ana_0.comparator_1.vnn.t50 avdd.t636 avdd.t395 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X385 dvss.t443 por_dig_0.net24 a_35330_33453# dvss.t442 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.06405 ps=0.725 w=0.42 l=0.15
X386 dvdd.t1059 a_40247_24823# a_40247_23627# dvdd.t1058 sky130_fd_pr__pfet_01v8_hvt ad=0.2968 pd=2.77 as=0.2968 ps=2.77 w=1.12 l=0.15
X387 dvdd.t65 por_ana_0.sky130_fd_sc_hd__inv_4_3.Y dcomp.t30 dvdd.t64 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X388 dvss.t965 por_dig_0.net25 a_36002_31277# dvss.t964 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X389 dvss.t1917 dvdd.t1826 dvss.t1916 dvss.t1915 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X390 a_37320_30733# a_36696_30739# a_37212_31111# dvdd.t1066 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X391 dvdd.t1555 dvss.t2245 dvdd.t1554 dvdd.t1553 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X392 por_ana_0.rstring_mux_0.vtrip_decoded_b_avdd[1] por_ana_0.rstring_mux_0.vtrip_decoded_avdd[1] avss.t318 avss.t317 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X393 dvdd.t736 por_dig_0.net7.t4 a_35130_28673# dvdd.t735 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.074375 ps=0.815 w=0.42 l=0.15
X394 por_ana_0.comparator_0.vpp.t17 vbg_1v2.t6 por_ana_0.comparator_0.vt.t52 por_ana_0.comparator_0.vt.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X395 dvss.t204 a_34098_30707# por_dig_0.clknet_1_0__leaf_osc_ck.t12 dvss.t203 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X396 a_33996_35389# por_dig_0.net24 dvdd.t359 dvdd.t358 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X397 dvdd.t982 por_dig_0.net22.t9 a_33804_31251# dvdd.t981 sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.22 ps=1.44 w=1 l=0.15
X398 a_33366_33453# por_dig_0.net22.t10 a_33282_33453# dvss.t1170 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X399 por_ana_0.rstring_mux_0.vtop.t13 por_ana_0.rstring_mux_0.ena_b avdd.t245 avdd.t244 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X400 por_ana_0.rc_osc_0.vr dvss.t1673 dvss.t1675 dvss.t1674 sky130_fd_pr__nfet_01v8 ad=0.1475 pd=1.295 as=0.145 ps=1.29 w=1 l=0.6
X401 por_ana_0.comparator_0.vpp.t18 vbg_1v2.t7 por_ana_0.comparator_0.vt.t51 por_ana_0.comparator_0.vt.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X402 dvdd.t1558 dvss.t2246 dvdd.t1557 dvdd.t1556 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X403 a_37688_33997# a_37064_34003# a_37580_34375# dvdd.t1076 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X404 por_ana_0.rstring_mux_0.otrip_decoded_b_avdd[5] por_ana_0.rstring_mux_0.otrip_decoded_avdd[5] avss.t262 avss.t261 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X405 avdd.t150 avdd.t148 avdd.t149 avdd.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=8
X406 a_37308_31111# a_36862_30739# a_37212_31111# dvss.t1276 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X407 dvdd.t583 a_36564_32339# por_dig_0.net23.t3 dvdd.t582 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X408 dvdd.t1560 dvss.t2247 dvdd.t1559 dvdd.t1556 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X409 por_ana_0.rstring_mux_0.vtrip_decoded_b_avdd[4] por_ana_0.rstring_mux_0.vtrip_decoded_avdd[4].t2 avdd.t573 avdd.t572 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X410 por_dig_0.otrip_decoded[2].t2 a_33752_28013# dvdd.t850 dvdd.t849 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X411 a_32651_31643# a_31932_31419# a_32088_31514# dvss.t25 sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0594 ps=0.69 w=0.36 l=0.15
X412 dvss.t1914 dvdd.t1827 dvss.t1913 dvss.t1734 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X413 por_ana_0.dcomp3v3 por_ana_0.comparator_1.n1.t4 avss.t25 avss.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X414 por_ana_0.comparator_0.vt.t34 avss.t411 por_ana_0.comparator_0.vnn.t21 por_ana_0.comparator_0.vt.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=8
X415 dvss.t403 a_39887_23089# a_39887_21959# dvss.t402 sky130_fd_pr__nfet_g5v0d10v5 ad=0.178875 pd=1.26 as=0.1197 ps=1.41 w=0.42 l=0.5
X416 por_dig_0.clknet_1_0__leaf_osc_ck.t11 a_34098_30707# dvss.t202 dvss.t201 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X417 dvdd.t1506 por_dig_0._030_ a_39738_32909# dvdd.t1505 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X418 a_29802_24707# a_29702_24619# dvss.t1544 dvss.t1543 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X419 por_ana_0.ibias_gen_0.ena_b.t3 por_ana_0.rstring_mux_0.ena.t3 avss.t383 avss.t382 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=1
X420 por_ana_0.comparator_0.vinn.t35 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[2] por_ana_0.rstring_mux_0.vtrip2.t4 avss.t266 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X421 avss.t269 por_ana_0.comparator_0.n1.t6 por_ana_0.dcomp3v3uv avss.t268 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X422 dvdd.t448 por_ana_0.rc_osc_0.m por_ana_0.rc_osc_0.n.t3 dvdd.t447 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X423 dvss.t495 por_dig_0.clknet_1_0__leaf_osc_ck.t35 a_32464_32915# dvss.t494 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X424 a_34378_30189# a_34212_30189# dvdd.t1084 dvdd.t1083 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X425 a_32019_31643# a_31932_31419# a_31615_31529# dvdd.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.0588 ps=0.7 w=0.42 l=0.15
X426 dvdd.t1563 dvss.t2248 dvdd.t1562 dvdd.t1561 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X427 por_ana_0.ibias_gen_0.vn0.t8 vbg_1v2.t8 por_ana_0.ibias_gen_0.vstart.t7 avss.t150 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X428 por_ana_0.comparator_0.vt.t33 avss.t412 por_ana_0.comparator_0.vnn.t20 por_ana_0.comparator_0.vt.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=8
X429 a_30260_13935# a_30638_6535# avss.t267 sky130_fd_pr__res_xhigh_po_1p41 l=35
X430 avss.t140 por_ana_0.sky130_fd_sc_hvl__inv_4_0.A por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.t5 avss.t139 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X431 dvdd.t269 a_32610_35603# por_dig_0._007_ dvdd.t268 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X432 a_35848_31643# a_35224_31277# a_35740_31277# dvdd.t1092 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X433 dvss.t1672 dvss.t1670 force_ena_rc_osc.t1 dvss.t1671 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X434 dvss.t1300 a_30070_23637# a_30495_23593# dvss.t1299 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X435 a_39262_34317# por_dig_0.cnt_st\[1\] por_dig_0._029_ dvss.t602 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X436 por_ana_0.comparator_1.vpp.t32 vin.t51 por_ana_0.comparator_1.vt.t34 por_ana_0.comparator_1.vt.t18 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X437 por_ana_0.comparator_1.vnn.t29 por_ana_0.comparator_1.vpp.t48 avdd.t404 avdd.t403 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X438 a_15886_35244# a_16264_27844# avss.t365 sky130_fd_pr__res_xhigh_po_1p41 l=35
X439 dvss.t871 por_dig_0.net23.t7 a_35746_36539# dvss.t870 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X440 a_31772_13935# a_31394_6535# avss.t366 sky130_fd_pr__res_xhigh_po_1p41 l=35
X441 por_dig_0.cnt_st\[2\] a_38136_33213# dvdd.t1052 dvdd.t1051 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X442 dvss.t1357 por_dig_0.net3 por_dig_0.net9 dvss.t1356 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X443 avdd.t269 a_34026_22973# a_35233_22637# avdd.t268 sky130_fd_pr__pfet_g5v0d10v5 ad=0.24375 pd=1.825 as=0.3975 ps=3.53 w=1.5 l=0.5
X444 avss.t119 avss.t118 por_ana_0.ibias_gen_0.ve.t1 sky130_fd_pr__pnp_05v5_W0p68L0p68
**devattr s=18496,544 d=4547244,10712
X445 por_ana_0.comparator_1.vpp.t33 vin.t52 por_ana_0.comparator_1.vt.t33 por_ana_0.comparator_1.vt.t18 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X446 dvss.t1912 dvdd.t1828 dvss.t1911 dvss.t1910 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X447 a_33378_34317# por_dig_0._019_ dvss.t2182 dvss.t2181 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X448 a_31615_33705# a_31893_33721# a_31849_33819# dvdd.t409 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0567 ps=0.69 w=0.42 l=0.15
X449 por.t10 por_ana_0.sky130_fd_sc_hd__inv_4_4.Y dvss.t1157 dvss.t1156 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X450 por_ana_0.rstring_mux_0.vtrip3.t9 por_ana_0.rstring_mux_0.vtrip4.t7 avss.t367 sky130_fd_pr__res_xhigh_po_1p41 l=35
X451 dvdd.t1268 a_33996_36477# a_33983_36173# dvdd.t1267 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X452 a_37584_30189# a_37138_30189# a_37488_30189# dvss.t2037 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X453 por_dig_0._046_ por_dig_0.net23.t8 dvdd.t759 dvdd.t758 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14575 ps=1.335 w=1 l=0.15
X454 a_35647_30189# por_dig_0.net25 dvss.t963 dvss.t962 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X455 a_32980_33287# a_32630_32915# a_32885_33275# dvdd.t860 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X456 a_19666_35244# a_20044_27844# avss.t368 sky130_fd_pr__res_xhigh_po_1p41 l=35
X457 dvss.t2039 a_36476_30163# a_36218_30163# dvss.t2038 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.5
X458 dvdd.t297 por_ana_0.sky130_fd_sc_hd__inv_4_1.Y porb.t28 dvdd.t296 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X459 por_dig_0.net21 a_38936_32159# dvss.t2043 dvss.t2042 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X460 dvss.t2056 a_31814_24619# a_31914_24707# dvss.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X461 a_22700_13935# a_23078_6535# avss.t369 sky130_fd_pr__res_xhigh_po_1p41 l=35
X462 dvss.t1909 dvdd.t1829 dvss.t1908 dvss.t1907 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X463 por_dig_0.net3 a_31360_28557# dvss.t697 dvss.t696 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X464 a_18154_35244# a_18532_27844# avss.t370 sky130_fd_pr__res_xhigh_po_1p41 l=35
X465 a_36690_35629# a_35500_35629# a_36581_35629# dvss.t526 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X466 por_ana_0.comparator_0.vinn.t45 por_ana_0.rstring_mux_0.vtrip_decoded_b_avdd[2] por_ana_0.rstring_mux_0.vtrip2.t9 avdd.t591 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X467 avdd.t630 por_ana_0.comparator_1.vnn.t10 por_ana_0.comparator_1.vnn.t11 avdd.t401 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X468 por_ana_0.comparator_1.vpp.t21 por_ana_0.comparator_1.vnn.t51 avdd.t637 avdd.t395 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X469 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.t4 por_ana_0.sky130_fd_sc_hvl__inv_4_0.A avss.t138 avss.t137 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.21375 ps=2.07 w=0.75 l=0.5
X470 por_ana_0.rstring_mux_0.otrip_decoded_b_avdd[6] por_ana_0.rstring_mux_0.otrip_decoded_avdd[6] avdd.t593 avdd.t592 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X471 a_15130_35244# a_15508_27844# avss.t375 sky130_fd_pr__res_xhigh_po_1p41 l=35
X472 a_38250_22973# a_38150_22885# dvss.t112 dvss.t111 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X473 porb.t27 por_ana_0.sky130_fd_sc_hd__inv_4_1.Y dvdd.t295 dvdd.t294 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X474 avdd.t599 a_23466_22973# a_24159_21859# avdd.t598 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.1365 ps=1.49 w=0.42 l=1
X475 avdd.t529 por_ana_0.comparator_1.n1.t5 por_ana_0.dcomp3v3 avdd.t528 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X476 por_dig_0.cnt_por\[3\] a_33996_35389# dvdd.t1072 dvdd.t1071 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X477 por_dig_0.clknet_1_1__leaf_osc_ck.t28 a_35583_34541# dvdd.t495 dvdd.t494 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X478 dvdd.t131 a_34387_32909# por_dig_0.clknet_0_osc_ck.t30 dvdd.t130 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X479 por_ana_0.schmitt_trigger_0.out.t3 por_ana_0.schmitt_trigger_0.m.t14 dvdd.t553 dvdd.t552 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X480 por_dig_0._034_.t0 por_dig_0.cnt_por\[3\] dvdd.t382 dvdd.t381 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X481 dvdd.t63 por_ana_0.sky130_fd_sc_hd__inv_4_3.Y dcomp.t29 dvdd.t62 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X482 vin.t47 por_ana_0.rstring_mux_0.otrip_decoded_avdd[4] por_ana_0.rstring_mux_0.vtrip4.t9 avss.t379 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X483 por_dig_0.clknet_1_1__leaf_osc_ck.t14 a_35583_34541# dvss.t594 dvss.t593 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X484 dcomp.t10 por_ana_0.sky130_fd_sc_hd__inv_4_3.Y dvss.t69 dvss.t68 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X485 dvss.t2049 por_dig_0.net21 a_38957_32883# dvss.t2048 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.091 ps=0.93 w=0.65 l=0.15
X486 dvdd.t1566 dvss.t2249 dvdd.t1565 dvdd.t1564 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X487 por_ana_0.schmitt_trigger_0.m.t1 por_ana_0.schmitt_trigger_0.in.t2 dvss.t651 dvss.t650 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X488 a_31914_24707# a_31814_24619# dvss.t2055 dvss.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X489 a_19094_1626# a_41694_2004# dvss.t2062 sky130_fd_pr__res_xhigh_po_1p41 l=111
X490 a_35942_31821# por_dig_0._035_ a_35858_31821# dvdd.t1390 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X491 por_ana_0.comparator_0.vnn avss.t413 por_ana_0.comparator_0.vt.t32 por_ana_0.comparator_0.vt.t18 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=8
X492 dvdd.t680 por_dig_0.net6 a_36649_28789# dvdd.t679 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1087 ps=1.36 w=0.42 l=0.15
X493 dvss.t13 a_32182_23637# a_32607_23593# dvss.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X494 por_dig_0.net27 a_34852_31277# dvss.t2071 dvss.t2070 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X495 dvdd.t1399 a_31413_29619# por_dig_0.osc_ena.t3 dvdd.t70 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X496 por_ana_0.rstring_mux_0.vtrip0.t8 por_ana_0.rstring_mux_0.otrip_decoded_avdd[0] vin.t35 avss.t309 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=0.6
X497 dvdd.t1568 dvss.t2250 dvdd.t1567 dvdd.t1522 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X498 dvss.t497 por_dig_0.clknet_1_0__leaf_osc_ck.t36 a_31360_31827# dvss.t496 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X499 avdd.t325 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.t11 porb_h.t14 avdd.t324 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X500 avdd.t147 avdd.t146 avdd.t147 avdd.t13 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=8
X501 dvss.t1906 dvdd.t1830 dvss.t1905 dvss.t1904 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X502 a_34357_33427# por_dig_0.cnt_por\[5\] a_34486_33703# dvdd.t1404 sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X503 por_ana_0.ibias_gen_0.vn0.t17 por_ana_0.ibias_gen_0.ena_b.t4 avss.t324 avss.t323 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X504 por_dig_0.otrip_decoded[1] a_32701_28531# dvss.t3 dvss.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X505 avdd.t211 a_36138_22973# a_37345_22637# avdd.t210 sky130_fd_pr__pfet_g5v0d10v5 ad=0.24375 pd=1.825 as=0.3975 ps=3.53 w=1.5 l=0.5
X506 dvss.t1903 dvdd.t1831 dvss.t1902 dvss.t1700 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X507 a_35930_28013# por_dig_0.net6 a_35858_28013# dvss.t677 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X508 dvdd.t1410 a_36512_28013# por_dig_0.otrip_decoded[5].t3 dvdd.t1409 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X509 por_ana_0.sky130_fd_sc_hd__inv_4_1.A por_dig_0.por_unbuf.t7 dvdd.t690 dvdd.t689 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X510 por_ana_0.sky130_fd_sc_hd__inv_4_0.Y por_ana_0.schmitt_trigger_0.out.t6 dvdd.t706 dvdd.t705 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X511 dvdd.t1571 dvss.t2251 dvdd.t1570 dvdd.t1569 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X512 a_39328_34515# por_dig_0.cnt_st\[0\] dvss.t1337 dvss.t1336 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X513 a_36480_31251# a_36305_31277# a_36659_31277# dvss.t2089 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X514 pwup_filt.t28 por_ana_0.sky130_fd_sc_hd__inv_4_0.Y dvdd.t219 dvdd.t218 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X515 a_31615_33705# a_31932_33595# a_31890_33453# dvss.t2093 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0669 ps=0.75 w=0.36 l=0.15
X516 a_36567_32141# por_dig_0._034_.t11 dvss.t863 dvss.t862 sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.203125 ps=1.275 w=0.65 l=0.15
X517 por_ana_0.rstring_mux_0.vtrip7.t4 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[7].t3 por_ana_0.comparator_0.vinn.t47 avss.t393 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X518 dvss.t224 por_ana_0.sky130_fd_sc_hd__inv_4_1.A por_ana_0.sky130_fd_sc_hd__inv_4_1.Y dvss.t223 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X519 vin.t41 por_ana_0.rstring_mux_0.otrip_decoded_b_avdd[4] por_ana_0.rstring_mux_0.vtrip4.t6 avdd.t561 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X520 a_24968_13935# a_24590_6535# avss.t320 sky130_fd_pr__res_xhigh_po_1p41 l=35
X521 a_40247_24823# a_40247_23627# dvdd.t1062 dvdd.t1061 sky130_fd_pr__pfet_01v8_hvt ad=0.2968 pd=2.77 as=0.1568 ps=1.4 w=1.12 l=0.15
X522 dvdd.t61 por_ana_0.sky130_fd_sc_hd__inv_4_3.Y dcomp.t28 dvdd.t60 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X523 a_37392_31251# por_dig_0.net34 a_37611_31277# dvss.t990 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.091 ps=0.93 w=0.65 l=0.15
X524 por_dig_0._002_ por_dig_0._039_ dvdd.t1298 dvdd.t1297 sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.39 as=0.182 ps=1.92 w=0.7 l=0.15
X525 dvdd.t1057 a_38956_32339# por_dig_0._031_ dvdd.t1056 sky130_fd_pr__pfet_01v8_hvt ad=0.31245 pd=1.68 as=0.26 ps=2.52 w=1 l=0.15
X526 a_33012_33997# por_dig_0._025_ dvdd.t1302 dvdd.t1301 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X527 pwup_filt.t15 por_ana_0.sky130_fd_sc_hd__inv_4_0.Y dvss.t258 dvss.t257 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X528 dvdd.t1574 dvss.t2252 dvdd.t1573 dvdd.t1572 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
R0 por_dig_0.net26 dvdd sky130_fd_pr__res_generic_po w=0.48 l=0.045
X529 dvdd.t446 por_ana_0.rc_osc_0.m por_ana_0.rc_osc_0.n.t2 dvdd.t445 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X530 dvdd.t243 por_ana_0.rc_osc_0.in por_ana_0.rc_osc_0.m dvdd.t242 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X531 dvdd.t692 por_dig_0.por_unbuf.t8 por_ana_0.sky130_fd_sc_hd__inv_4_1.A dvdd.t691 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X532 dvdd.t93 a_35030_28557# a_35130_28673# dvdd.t92 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1085 ps=1.36 w=0.42 l=0.15
X533 a_37430_30707# a_37212_31111# dvdd.t1068 dvdd.t1067 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X534 dvdd.t217 por_ana_0.sky130_fd_sc_hd__inv_4_0.Y pwup_filt.t27 dvdd.t216 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X535 por_dig_0.cnt_por\[9\] a_35468_30163# dvss.t544 dvss.t543 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X536 a_36124_35995# a_35500_35629# a_36016_35629# dvdd.t440 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X537 por_dig_0._043_ a_39497_30849# dvdd.t1306 dvdd.t1305 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X538 dvdd.t1451 por_dig_0.clknet_0_osc_ck.t33 a_34098_30707# dvdd.t1450 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X539 por_ana_0.comparator_1.vt.t32 vin.t53 por_ana_0.comparator_1.vpp.t34 por_ana_0.comparator_1.vt.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X540 a_32462_32607# a_32244_32365# dvss.t1359 dvss.t1358 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X541 por_ana_0.rstring_mux_0.vtrip_decoded_b_avdd[3] por_ana_0.rstring_mux_0.vtrip_decoded_avdd[3] avdd.t179 avdd.t178 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X542 a_32340_32365# a_31894_32365# a_32244_32365# dvss.t1972 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X543 avdd.t564 a_25578_22973# a_26271_21859# avdd.t563 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.1365 ps=1.49 w=0.42 l=1
X544 dvss.t1976 a_38444_28013# por_dig_0.otrip_decoded[0].t1 dvss.t523 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X545 avdd.t145 avdd.t144 avdd.t145 avdd.t13 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=8
X546 avss.t29 por_ana_0.rstring_mux_0.ena_b por_ana_0.rstring_mux_0.vtop.t16 avss.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X547 a_34282_35629# por_dig_0.cnt_por\[0\].t9 a_34198_35629# dvss.t637 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X548 dvdd.t1577 dvss.t2253 dvdd.t1576 dvdd.t1575 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X549 a_36331_33819# a_35573_33721# a_35768_33690# dvdd.t1318 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.07245 ps=0.765 w=0.42 l=0.15
X550 por_ana_0.comparator_1.vt.t31 vin.t54 por_ana_0.comparator_1.vpp.t35 por_ana_0.comparator_1.vt.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X551 por_ana_0.rstring_mux_0.vtrip0.t5 por_ana_0.rstring_mux_0.otrip_decoded_b_avdd[0] vin.t22 avdd.t429 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=0.6
X552 dvss.t1901 dvdd.t1832 dvss.t1900 dvss.t1812 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X553 dvdd.t1149 a_33198_32883# a_33088_32909# dvdd.t1148 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X554 otrip[1].t1 dvss.t1667 dvss.t1669 dvss.t1668 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X555 dvdd.t1397 por_dig_0.net27 a_36328_29645# dvdd.t70 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.265 ps=2.53 w=1 l=0.15
X556 a_15130_35244# a_14752_27844# avss.t321 sky130_fd_pr__res_xhigh_po_1p41 l=35
X557 avss.t117 avss.t115 avss.t116 avss.t81 sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0 ps=0 w=5 l=8
X558 a_20432_13935# a_20054_6535# avss.t322 sky130_fd_pr__res_xhigh_po_1p41 l=35
X559 avdd.t629 por_ana_0.comparator_1.vnn.t8 por_ana_0.comparator_1.vnn.t9 avdd.t401 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X560 por_timed_out.t0 a_31413_32339# dvss.t835 dvss.t834 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X561 dvss.t1899 dvdd.t1833 dvss.t1898 dvss.t1897 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X562 dvss.t1155 por_ana_0.sky130_fd_sc_hd__inv_4_4.Y por.t9 dvss.t1154 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X563 a_32800_31111# a_32354_30739# a_32704_31111# dvss.t2233 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X564 por_dig_0.cnt_st\[0\] a_38320_34301# dvss.t830 dvss.t829 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X565 por_ana_0.rstring_mux_0.vtrip7.t0 por_ana_0.rstring_mux_0.vtrip_decoded_b_avdd[7] por_ana_0.comparator_0.vinn.t26 avdd.t433 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X566 vin.t20 avss.t113 vin.t20 avss.t114 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=0.6
X567 avdd.t143 avdd.t142 avdd.t143 avdd.t33 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=8
X568 dvss.t2092 a_31932_33595# a_31893_33721# dvss.t2091 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X569 dvdd.t1580 dvss.t2254 dvdd.t1579 dvdd.t1578 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X570 porb.t26 por_ana_0.sky130_fd_sc_hd__inv_4_1.Y dvdd.t293 dvdd.t292 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X571 ibg_200n.t0 por_ana_0.rstring_mux_0.ena.t4 a_13894_21948# avss.t384 sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=0.6
X572 por_ana_0.comparator_1.vt.t30 vin.t55 por_ana_0.comparator_1.vpp.t36 por_ana_0.comparator_1.vt.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X573 a_36581_35629# a_35666_35629# a_36234_35871# dvss.t620 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X574 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[4].t0 a_35233_22637# avdd.t586 avdd.t268 sky130_fd_pr__pfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.24375 ps=1.825 w=1.5 l=0.5
X575 dvss.t1896 dvdd.t1834 dvss.t1895 dvss.t1894 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X576 por.t8 por_ana_0.sky130_fd_sc_hd__inv_4_4.Y dvss.t1153 dvss.t1152 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X577 a_34580_34110# por_dig_0.net22.t11 dvdd.t984 dvdd.t983 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X578 dvss.t101 por_dig_0.net4 a_35040_34587# dvss.t100 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X579 dvss.t1987 a_27690_22973# a_28897_22637# dvss.t1986 sky130_fd_pr__nfet_g5v0d10v5 ad=0.121875 pd=1.075 as=0.19875 ps=2.03 w=0.75 l=0.5
X580 a_36122_30341# a_36218_30163# dvss.t2041 dvss.t2040 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.5
X581 avss.t148 por_ana_0.comparator_1.n0.t6 por_ana_0.comparator_1.n1.t3 avss.t147 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X582 dvdd.t291 por_ana_0.sky130_fd_sc_hd__inv_4_1.Y porb.t25 dvdd.t290 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X583 por_ana_0.comparator_1.vt.t29 vin.t56 por_ana_0.comparator_1.vpp.t37 por_ana_0.comparator_1.vt.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X584 a_33896_35603# por_dig_0.cnt_por\[3\] dvss.t455 dvss.t454 sky130_fd_pr__nfet_01v8 ad=0.183625 pd=1.215 as=0.160875 ps=1.145 w=0.65 l=0.15
X585 a_38315_33453# por_dig_0.net25 dvss.t961 dvss.t408 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X586 a_32885_33275# por_dig_0._010_ dvss.t1993 dvss.t1992 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X587 dvss.t1995 por_dig_0._026_ a_34486_32365# dvss.t460 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X588 a_34024_33703# por_dig_0._047_ a_33806_33427# dvdd.t727 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.26 ps=2.52 w=1 l=0.15
X589 dvdd.t1582 dvss.t2255 dvdd.t1581 dvdd.t1556 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X590 por_ana_0.ibias_gen_0.vn0.t9 vbg_1v2.t9 por_ana_0.ibias_gen_0.vstart.t6 avss.t150 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X591 dvdd.t1326 a_33896_35603# por_dig_0._053_ dvdd.t1325 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X592 a_34387_32909# osc_ck.t9 dvdd.t774 dvdd.t773 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X593 por_ana_0.comparator_0.vpp.t13 por_ana_0.comparator_0.vpp.t12 avdd.t203 avdd.t191 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X594 dvss.t1534 por_dig_0.otrip_decoded[4] a_25478_22885# dvss.t1533 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X595 a_36002_31277# a_35958_31519# a_35836_31277# dvss.t930 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X596 por_dig_0.clknet_0_osc_ck.t29 a_34387_32909# dvdd.t129 dvdd.t128 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X597 dvdd.t1439 por_dig_0.net5.t3 a_35776_28013# dvdd.t1438 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X598 dvdd.t1337 a_36376_28789# por_dig_0.net16 dvdd.t1336 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.26 ps=2.52 w=1 l=0.15
X599 dvss.t2129 por_dig_0.clknet_0_osc_ck.t34 a_35583_34541# dvss.t2128 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X600 a_36831_23593# a_36406_23637# dvss.t978 dvss.t977 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X601 a_35330_32141# por_dig_0.cnt_por\[8\] a_35227_32141# dvss.t319 sky130_fd_pr__nfet_01v8 ad=0.118625 pd=1.015 as=0.118625 ps=1.015 w=0.65 l=0.15
X602 a_30070_23637# a_29702_24619# dvss.t1542 dvss.t1541 sky130_fd_pr__nfet_01v8 ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X603 avdd.t217 a_26288_32594# a_25595_33708# avdd.t216 sky130_fd_pr__pfet_g5v0d10v5 ad=0.2142 pd=1.99 as=0.2142 ps=1.99 w=0.42 l=1
X604 vin.t8 avdd.t140 vin.t8 avdd.t141 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=0.6
X605 por_ana_0.rstring_mux_0.vtop.t12 por_ana_0.rstring_mux_0.ena_b avdd.t243 avdd.t242 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X606 dvss.t2005 a_31412_31251# por_dig_0.cnt_rsb_stg1 dvss.t2004 sky130_fd_pr__nfet_01v8 ad=0.2087 pd=2.02 as=0.169 ps=1.82 w=0.65 l=0.15
X607 avdd.t139 avdd.t137 avdd.t138 avdd.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=8
X608 a_31849_33819# a_31412_33427# dvdd.t1347 dvdd.t1346 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X609 dvss.t286 a_38136_33427# a_38070_33453# dvss.t285 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X610 a_12598_23626# por_ana_0.ibias_gen_0.ena_b.t5 por_ana_0.ibias_gen_0.vstart.t10 avdd.t570 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=0.6
X611 dvss.t1151 por_ana_0.sky130_fd_sc_hd__inv_4_4.Y por.t7 dvss.t1150 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X612 avdd.t568 a_27690_22973# a_28383_21859# avdd.t567 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.1365 ps=1.49 w=0.42 l=1
X613 a_29802_22973# a_29702_22885# dvss.t487 dvss.t486 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X614 a_36526_28917# por_dig_0.net7.t5 dvss.t849 dvss.t848 sky130_fd_pr__nfet_01v8 ad=0.05355 pd=0.675 as=0.122275 ps=1.08 w=0.42 l=0.15
X615 dvss.t960 por_dig_0.net25 a_37658_33453# dvss.t406 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X616 dvss.t161 a_34387_32909# por_dig_0.clknet_0_osc_ck.t13 dvss.t160 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X617 dvdd.t1585 dvss.t2256 dvdd.t1584 dvdd.t1583 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X618 por_ana_0.rc_osc_0.in a_41694_492# dvss.t1178 sky130_fd_pr__res_xhigh_po_1p41 l=111
X619 por_ana_0.comparator_1.vpp.t16 por_ana_0.rstring_mux_0.ena.t5 avdd.t606 avdd.t605 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X620 avdd.t432 a_36831_23593# a_36138_24707# avdd.t431 sky130_fd_pr__pfet_g5v0d10v5 ad=0.2142 pd=1.99 as=0.2142 ps=1.99 w=0.42 l=1
X621 dvss.t1893 dvdd.t1835 dvss.t1892 dvss.t1891 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X622 porb.t24 por_ana_0.sky130_fd_sc_hd__inv_4_1.Y dvdd.t289 dvdd.t288 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X623 dvss.t1180 a_32088_33690# a_32019_33819# dvss.t1179 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0999 ps=0.985 w=0.64 l=0.15
X624 por_ana_0.sky130_fd_sc_hd__inv_4_3.Y por_ana_0.vl dvss.t1188 dvss.t1187 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X625 avdd.t457 a_30495_21859# a_29802_22973# avdd.t456 sky130_fd_pr__pfet_g5v0d10v5 ad=0.2142 pd=1.99 as=0.2142 ps=1.99 w=0.42 l=1
X626 a_26271_21859# a_25846_21903# dvss.t1004 dvss.t1003 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X627 dcomp.t9 por_ana_0.sky130_fd_sc_hd__inv_4_3.Y dvss.t67 dvss.t66 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X628 por_dig_0.clknet_1_1__leaf_osc_ck.t27 a_35583_34541# dvdd.t493 dvdd.t492 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X629 a_38250_24707# a_38150_24619# dvss.t46 dvss.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X630 dvss.t1192 a_39732_31829# startup_timed_out.t1 dvss.t1191 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X631 a_34830_35629# por_dig_0.cnt_por\[0\].t10 a_35024_35629# dvss.t638 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X632 dvss.t2221 a_38518_23637# a_38943_23593# dvss.t2220 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X633 dvss.t373 por_dig_0.net30 a_33852_29645# dvss.t372 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X634 por_ana_0.comparator_1.n0.t1 por_ana_0.comparator_1.vpp.t49 avdd.t405 avdd.t403 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X635 dvdd.t1277 por_dig_0.cnt_por\[2\] por_dig_0._034_.t8 dvdd.t1276 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X636 dvss.t873 por_dig_0.net23.t9 a_34482_34541# dvss.t872 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X637 a_39022_32159# por_dig_0.cnt_st\[4\] a_38936_32159# dvss.t1530 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X638 dcomp.t27 por_ana_0.sky130_fd_sc_hd__inv_4_3.Y dvdd.t59 dvdd.t58 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X639 a_35433_32141# por_dig_0.net23.t10 a_35330_32141# dvss.t874 sky130_fd_pr__nfet_01v8 ad=0.19825 pd=1.26 as=0.118625 ps=1.015 w=0.65 l=0.15
X640 por_ana_0.dcomp3v3 por_ana_0.comparator_1.n1.t6 avdd.t531 avdd.t530 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X641 a_39177_33229# por_dig_0._040_ dvss.t1194 dvss.t1193 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.26 ps=1.45 w=0.65 l=0.15
X642 dvss.t653 por_ana_0.schmitt_trigger_0.in.t3 por_ana_0.schmitt_trigger_0.m.t0 dvss.t652 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X643 dvss.t65 por_ana_0.sky130_fd_sc_hd__inv_4_3.Y dcomp.t8 dvss.t64 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X644 a_13628_13935# a_13250_6535# avss.t247 sky130_fd_pr__res_xhigh_po_1p41 l=35
X645 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[6].t0 a_37345_22637# avdd.t602 avdd.t210 sky130_fd_pr__pfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.24375 ps=1.825 w=1.5 l=0.5
X646 dvss.t1252 a_37392_31251# por_dig_0._004_ dvss.t1251 sky130_fd_pr__nfet_01v8 ad=0.258375 pd=1.445 as=0.169 ps=1.82 w=0.65 l=0.15
X647 por_dig_0.cnt_rsb a_32616_32125# dvdd.t397 dvdd.t396 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X648 dvss.t2047 por_dig_0.net21 por_dig_0._039_ dvss.t2046 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X649 dvdd.t1119 a_39718_33605# por_dig_0._040_ dvdd.t1118 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.34 ps=2.68 w=1 l=0.15
X650 dvdd.t1182 por_dig_0.net8 a_31864_30823# dvdd.t1181 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X651 a_34746_31277# a_34510_31277# dvdd.t395 dvdd.t394 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.5
X652 a_35858_31821# por_dig_0._037_ por_dig_0.net19 dvdd.t98 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X653 por_ana_0.comparator_1.n0.t2 por_ana_0.comparator_1.ena_b avss.t257 avss.t256 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X654 a_14384_13935# a_14762_6535# avss.t248 sky130_fd_pr__res_xhigh_po_1p41 l=35
X655 dvss.t1666 dvss.t1664 otrip[0].t1 dvss.t1665 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X656 dvdd.t491 a_35583_34541# por_dig_0.clknet_1_1__leaf_osc_ck.t26 dvdd.t490 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X657 por_ana_0.rstring_mux_0.vtrip_decoded_b_avdd[5] por_ana_0.rstring_mux_0.vtrip_decoded_avdd[5].t2 avss.t301 avss.t300 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X658 dvss.t1405 por_dig_0.cnt_por\[1\] por_dig_0._049_ dvss.t1404 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X659 dvdd.t1104 force_dis_rc_osc.t2 a_31360_33997# dvdd.t1103 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X660 a_32609_31099# por_dig_0._013_ dvss.t1206 dvss.t1205 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X661 dvdd.t1587 dvss.t2257 dvdd.t1586 dvdd.t1556 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X662 dvss.t499 por_dig_0.clknet_1_0__leaf_osc_ck.t37 a_34212_30189# dvss.t498 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X663 dvdd.t251 por_dig_0._042_ a_39728_31527# dvdd.t250 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X664 avdd.t327 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.t12 porb_h.t13 avdd.t326 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X665 dvdd.t1494 por_dig_0._019_ a_34212_33997# dvdd.t1493 sky130_fd_pr__pfet_01v8_hvt ad=0.1475 pd=1.295 as=0.265 ps=2.53 w=1 l=0.15
X666 a_32326_31277# por_dig_0.net8 dvss.t1427 dvss.t1426 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1346 ps=1.15 w=0.42 l=0.15
X667 force_pdn.t1 dvss.t1661 dvss.t1663 dvss.t1662 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X668 a_32704_31111# a_32354_30739# a_32609_31099# dvdd.t1521 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X669 por_ana_0.comparator_1.vnn.t45 vbg_1v2.t10 por_ana_0.comparator_1.vt.t52 por_ana_0.comparator_1.vt.t36 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X670 dvss.t560 a_36756_35603# por_dig_0.cnt_por\[0\].t1 dvss.t559 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X671 dvdd.t1589 dvss.t2258 dvdd.t1588 dvdd.t1583 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X672 ibg_200n.t1 por_ana_0.ibias_gen_0.ena_b.t6 a_13844_23626# avdd.t571 sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=0.6
X673 por_ana_0.rstring_mux_0.otrip_decoded_b_avdd[1] por_ana_0.rstring_mux_0.otrip_decoded_avdd[1] avdd.t259 avdd.t258 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X674 a_31890_31277# a_31412_31251# dvss.t2003 dvss.t2002 sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.12495 ps=1.015 w=0.42 l=0.15
X675 por_ana_0.comparator_1.vt.t17 avss.t414 por_ana_0.comparator_1.vnn.t37 por_ana_0.comparator_1.vt.t3 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=8
X676 a_33352_35463# a_32906_35091# a_33256_35463# dvss.t1208 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X677 dvdd.t357 por_dig_0.net24 a_32233_33819# dvdd.t356 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1092 ps=1.36 w=0.42 l=0.15
X678 por_dig_0.cnt_st\[1\] a_38136_33427# dvss.t284 dvss.t283 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X679 a_31781_32187# por_dig_0.net28 dvss.t1210 dvss.t1209 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X680 dvss.t2108 por_dig_0.otrip_decoded[6].t5 a_27590_22885# dvss.t2107 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X681 a_36308_13935# a_35930_6535# avss.t249 sky130_fd_pr__res_xhigh_po_1p41 l=35
X682 a_38943_23593# a_38518_23637# dvss.t2219 dvss.t2218 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X683 a_32182_23637# a_31814_24619# dvss.t2054 dvss.t2053 sky130_fd_pr__nfet_01v8 ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X684 por_dig_0.otrip_decoded[5].t2 a_36512_28013# dvdd.t1408 dvdd.t1407 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X685 dvdd.t708 por_ana_0.schmitt_trigger_0.out.t7 por_ana_0.sky130_fd_sc_hd__inv_4_0.Y dvdd.t707 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X686 a_33474_35059# a_33256_35463# dvdd.t1036 dvdd.t1035 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X687 por_ana_0.comparator_0.vnn.t23 por_ana_0.comparator_0.vinn.t50 por_ana_0.comparator_0.vt.t15 por_ana_0.comparator_0.vt.t3 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X688 a_31914_22973# a_31814_22885# dvss.t2164 dvss.t2163 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X689 a_33374_31277# por_dig_0.net4 dvss.t99 dvss.t98 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X690 a_31727_30849# por_dig_0.net1 dvdd.t1482 dvdd.t1481 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.14825 ps=1.34 w=0.42 l=0.15
X691 por_ana_0.comparator_1.vt.t16 avss.t415 por_ana_0.comparator_1.vnn.t36 por_ana_0.comparator_1.vt.t3 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=8
X692 force_short_oneshot.t1 dvss.t1658 dvss.t1660 dvss.t1659 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X693 por_dig_0.net5.t0 a_32039_28013# dvss.t1212 dvss.t523 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X694 a_37064_13935# a_37442_6535# avss.t250 sky130_fd_pr__res_xhigh_po_1p41 l=35
X695 avdd.t656 a_38943_23593# a_38250_24707# avdd.t655 sky130_fd_pr__pfet_g5v0d10v5 ad=0.2142 pd=1.99 as=0.2142 ps=1.99 w=0.42 l=1
X696 dvdd.t1592 dvss.t2259 dvdd.t1591 dvdd.t1590 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X697 dvdd.t1275 por_dig_0.cnt_por\[2\] a_34672_35451# dvdd.t1274 sky130_fd_pr__pfet_01v8_hvt ad=0.31245 pd=1.68 as=0.0588 ps=0.7 w=0.42 l=0.15
X698 a_37138_30189# a_36972_30189# dvdd.t19 dvdd.t18 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X699 a_34022_31527# por_dig_0.net4 dvdd.t83 dvdd.t82 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.26 ps=2.52 w=1 l=0.15
X700 dvss.t1425 por_dig_0.net8 a_31650_31277# dvss.t1424 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.06405 ps=0.725 w=0.42 l=0.15
X701 por_ana_0.comparator_0.vt.t50 vbg_1v2.t11 por_ana_0.comparator_0.vpp.t19 por_ana_0.comparator_0.vt.t36 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X702 dvdd.t179 a_34098_30707# por_dig_0.clknet_1_0__leaf_osc_ck.t31 dvdd.t178 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X703 dvdd.t1595 dvss.t2260 dvdd.t1594 dvdd.t1593 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X704 por_ana_0.comparator_0.vinn.t21 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[6].t3 por_ana_0.rstring_mux_0.vtrip6.t2 avss.t210 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X705 dvdd.t177 a_34098_30707# por_dig_0.clknet_1_0__leaf_osc_ck.t30 dvdd.t176 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X706 avdd.t241 por_ana_0.rstring_mux_0.ena_b por_ana_0.rstring_mux_0.vtop.t11 avdd.t240 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X707 avdd.t263 a_32607_21859# a_31914_22973# avdd.t262 sky130_fd_pr__pfet_g5v0d10v5 ad=0.2142 pd=1.99 as=0.2142 ps=1.99 w=0.42 l=1
X708 a_28383_21859# a_27958_21903# dvss.t2202 dvss.t2201 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X709 dvdd.t1597 dvss.t2261 a_36038_22885# dvdd.t1596 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X710 dvss.t1890 dvdd.t1836 dvss.t1889 dvss.t1888 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X711 dvdd.t1028 a_31776_29864# por_dig_0.net2 dvdd.t1027 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X712 a_35640_32517# por_dig_0.cnt_por\[4\] dvdd.t1256 dvdd.t1255 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X713 avdd.t638 por_ana_0.comparator_1.vnn.t52 por_ana_0.comparator_1.vpp.t22 avdd.t392 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X714 dvdd.t1599 dvss.t2262 a_36038_24619# dvdd.t1598 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X715 a_31776_29864# force_ena_rc_osc.t2 dvdd.t1348 dvdd.t1027 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X716 por_dig_0._042_ por_dig_0.net4 dvdd.t81 dvdd.t80 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X717 por_ana_0.comparator_1.vt.t15 avss.t416 por_ana_0.comparator_1.vnn.t35 por_ana_0.comparator_1.vt.t3 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=8
X718 por_ana_0.comparator_0.vnn avss.t417 por_ana_0.comparator_0.vt.t31 por_ana_0.comparator_0.vt.t18 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=8
X719 a_34198_35629# por_dig_0.cnt_por\[1\] a_33896_35603# dvss.t1403 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.183625 ps=1.215 w=0.65 l=0.15
X720 a_37789_31821# por_dig_0._042_ a_37698_31821# dvdd.t249 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.1525 ps=1.305 w=1 l=0.15
X721 por_ana_0.comparator_1.vnn avss.t418 por_ana_0.comparator_1.vt.t14 por_ana_0.comparator_1.vt.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=8
X722 a_33097_34317# por_dig_0._024_ a_32794_33971# dvss.t1039 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.089375 ps=0.925 w=0.65 l=0.15
X723 dvdd.t1602 dvss.t2263 dvdd.t1601 dvdd.t1600 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X724 dvss.t2075 por_dig_0.net27 a_36328_29645# dvss.t2074 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.1113 ps=1.37 w=0.42 l=0.15
X725 dvdd.t1605 dvss.t2264 dvdd.t1604 dvdd.t1603 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X726 a_37842_34363# a_37798_33971# a_37676_34375# dvss.t687 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X727 dvdd.t718 a_38320_34301# a_38307_33997# dvdd.t717 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X728 por_ana_0.rstring_mux_0.ena.t0 a_39457_22637# avdd.t448 avdd.t447 sky130_fd_pr__pfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.24375 ps=1.825 w=1.5 l=0.5
X729 a_34580_33453# por_dig_0._033_ a_34486_33453# dvss.t36 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X730 por_ana_0.comparator_1.vt.t13 avss.t419 por_ana_0.comparator_1.vnn.t34 por_ana_0.comparator_1.vt.t3 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=8
X731 por_ana_0.comparator_0.vnn avss.t420 por_ana_0.comparator_0.vt.t30 por_ana_0.comparator_0.vt.t18 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=8
X732 a_39634_32615# por_dig_0.net33 por_dig_0._041_ dvdd.t903 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X733 por_ana_0.rstring_mux_0.vtrip2.t3 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[2] por_ana_0.comparator_0.vinn.t34 avss.t265 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X734 dvdd.t1345 a_31412_33427# por_dig_0.cnt_por\[6\] dvdd.t1103 sky130_fd_pr__pfet_01v8_hvt ad=0.3012 pd=2.66 as=0.26 ps=2.52 w=1 l=0.15
X735 por_ana_0.comparator_1.vnn avss.t421 por_ana_0.comparator_1.vt.t12 por_ana_0.comparator_1.vt.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=8
X736 a_33805_32339# por_dig_0.cnt_por\[6\] a_34028_32365# dvss.t458 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X737 por.t6 por_ana_0.sky130_fd_sc_hd__inv_4_4.Y dvss.t1149 dvss.t1148 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X738 por_ana_0.schmitt_trigger_0.m.t6 por_ana_0.schmitt_trigger_0.in.t4 dvdd.t561 dvdd.t560 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X739 dvdd.t761 por_dig_0.net23.t11 a_35776_36967# dvdd.t760 sky130_fd_pr__pfet_01v8_hvt ad=0.1475 pd=1.295 as=0.265 ps=2.53 w=1 l=0.15
X740 a_35954_34317# por_dig_0.net22.t12 dvss.t1172 dvss.t1171 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X741 dvdd.t1608 dvss.t2265 dvdd.t1607 dvdd.t1606 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X742 dvss.t83 a_35202_29877# por_dig_0.net30 dvss.t82 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X743 avdd.t422 a_29802_24707# a_30495_23593# avdd.t421 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.1365 ps=1.49 w=0.42 l=1
X744 por_dig_0._014_ por_dig_0._027_ a_34102_29965# dvss.t1050 sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.08775 ps=0.92 w=0.65 l=0.15
X745 a_32651_31643# a_31893_31545# a_32088_31514# dvdd.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.07245 ps=0.765 w=0.42 l=0.15
X746 dvss.t1147 por_ana_0.sky130_fd_sc_hd__inv_4_4.Y por.t5 dvss.t1146 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X747 por_ana_0.comparator_0.vinn.t41 por_ana_0.rstring_mux_0.vtrip_decoded_b_avdd[6] por_ana_0.rstring_mux_0.vtrip6.t4 avdd.t559 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X748 dvdd.t909 a_33269_31111# a_33444_31037# dvdd.t908 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X749 dvdd.t1224 a_36480_31251# a_36467_31643# dvdd.t1223 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X750 a_33076_33287# a_32630_32915# a_32980_33287# dvss.t984 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X751 dvss.t1657 dvss.t1655 a_29702_22885# dvss.t1656 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X752 por_ana_0.dcomp3v3uv por_ana_0.comparator_0.n1.t7 avss.t271 avss.t270 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X753 a_33088_32909# a_32464_32915# a_32980_33287# dvdd.t403 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X754 a_36756_35603# por_dig_0.net24 dvdd.t355 dvdd.t354 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X755 a_34028_32365# por_dig_0.net22.t13 a_33934_32365# dvss.t1173 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X756 por_ana_0.comparator_0.vnn.t10 por_ana_0.comparator_0.vpp.t50 avdd.t202 avdd.t182 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X757 a_34294_23637# a_33926_24619# dvss.t515 dvss.t514 sky130_fd_pr__nfet_01v8 ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X758 por_ana_0.comparator_1.vnn avss.t422 por_ana_0.comparator_1.vt.t11 por_ana_0.comparator_1.vt.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=8
X759 a_34026_22973# a_33926_22885# dvss.t614 dvss.t613 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X760 dvdd.t1273 por_dig_0.cnt_por\[2\] a_34114_35879# dvdd.t1272 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X761 dvdd.t509 por_dig_0.cnt_st\[1\] a_39634_32615# dvdd.t508 sky130_fd_pr__pfet_01v8_hvt ad=0.1475 pd=1.295 as=0.14 ps=1.28 w=1 l=0.15
X762 a_34486_32365# a_34444_32517# por_dig_0._013_ dvss.t1052 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.195 ps=1.9 w=0.65 l=0.15
X763 a_32462_32607# a_32244_32365# dvdd.t1129 dvdd.t1128 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X764 a_34387_32909# osc_ck.t10 dvdd.t776 dvdd.t775 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X765 por_ana_0.comparator_1.vnn avss.t423 por_ana_0.comparator_1.vt.t10 por_ana_0.comparator_1.vt.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=8
X766 dvss.t1054 por_dig_0._052_ a_32913_35629# dvss.t1053 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X767 a_34796_13935# a_34418_6535# avss.t236 sky130_fd_pr__res_xhigh_po_1p41 l=35
X768 dvss.t441 por_dig_0.net24 a_33518_36539# dvss.t440 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X769 a_37230_34003# a_37064_34003# dvdd.t1075 dvdd.t1074 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X770 avdd.t406 por_ana_0.comparator_1.vpp.t50 por_ana_0.comparator_1.vnn.t28 avdd.t401 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X771 dvdd.t1611 dvss.t2266 dvdd.t1610 dvdd.t1609 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X772 por_ana_0.rstring_mux_0.vtrip2.t8 por_ana_0.rstring_mux_0.vtrip_decoded_b_avdd[2] por_ana_0.comparator_0.vinn.t44 avdd.t590 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X773 avdd.t516 a_34719_21859# a_34026_22973# avdd.t515 sky130_fd_pr__pfet_g5v0d10v5 ad=0.2142 pd=1.99 as=0.2142 ps=1.99 w=0.42 l=1
X774 dvss.t159 a_34387_32909# por_dig_0.clknet_0_osc_ck.t12 dvss.t158 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X775 a_29802_24707# a_29702_24619# dvss.t1540 dvss.t1539 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X776 dvss.t1887 dvdd.t1837 dvss.t1886 dvss.t1682 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X777 avdd.t136 avdd.t135 avdd.t136 avdd.t33 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=8
X778 por_ana_0.rc_osc_0.in dvss.t293 sky130_fd_pr__cap_mim_m3_2 l=30 w=30
X779 a_38904_31277# por_dig_0._032_ dvss.t301 dvss.t300 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.08775 ps=0.92 w=0.65 l=0.15
X780 por_ana_0.rstring_mux_0.vtrip4.t8 por_ana_0.rstring_mux_0.otrip_decoded_avdd[4] vin.t46 avss.t378 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X781 dvss.t1885 dvdd.t1838 dvss.t1884 dvss.t1863 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X782 avdd.t201 por_ana_0.comparator_0.vpp.t10 por_ana_0.comparator_0.vpp.t11 avdd.t195 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X783 a_33364_35085# por_dig_0.net24 dvdd.t353 dvdd.t352 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X784 por_ana_0.rstring_mux_0.vtop.t10 por_ana_0.rstring_mux_0.ena_b avdd.t239 avdd.t238 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X785 a_19094_3138# a_41694_2760# dvss.t1057 sky130_fd_pr__res_xhigh_po_1p41 l=111
X786 dvss.t278 a_36038_22885# a_36138_22973# dvss.t277 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X787 dvss.t1883 dvdd.t1839 dvss.t1882 dvss.t1881 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X788 avdd.t200 por_ana_0.comparator_0.vpp.t51 por_ana_0.comparator_0.n0.t1 avdd.t180 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X789 dvss.t1298 a_30070_23637# a_30495_23593# dvss.t1297 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X790 dvdd.t916 a_35556_29619# a_35298_29619# dvdd.t325 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.5
X791 dvdd.t1106 por_dig_0.otrip_decoded[0].t4 a_21254_22885# dvdd.t1105 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X792 a_35583_34541# por_dig_0.clknet_0_osc_ck.t35 dvdd.t1453 dvdd.t1452 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X793 por_ana_0.rstring_mux_0.otrip_decoded_b_avdd[3] por_ana_0.rstring_mux_0.otrip_decoded_avdd[3] avss.t240 avss.t239 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X794 a_32398_31277# a_32019_31643# a_32326_31277# dvss.t1284 sky130_fd_pr__nfet_01v8 ad=0.1401 pd=1.1 as=0.0441 ps=0.63 w=0.42 l=0.15
X795 a_36124_35995# por_dig_0.net24 dvdd.t351 dvdd.t350 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X796 por_dig_0.clknet_1_1__leaf_osc_ck.t25 a_35583_34541# dvdd.t489 dvdd.t488 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X797 dvss.t1186 por_ana_0.vl por_ana_0.sky130_fd_sc_hd__inv_4_3.Y dvss.t1185 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X798 dvdd.t185 por_dig_0.otrip_decoded[1] a_21254_24619# dvdd.t184 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X799 a_37396_33453# a_37046_33453# a_37301_33453# dvdd.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X800 por_dig_0._011_ por_dig_0._048_ a_35040_34317# dvss.t1112 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X801 por_ana_0.comparator_0.n0.t0 por_ana_0.comparator_0.vpp.t52 avdd.t199 avdd.t182 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X802 dvss.t1880 dvdd.t1840 dvss.t1879 dvss.t1878 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X803 startup_timed_out.t0 a_39732_31829# dvss.t1190 dvss.t1189 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X804 a_37488_30189# a_37138_30189# a_37393_30189# dvdd.t1374 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X805 por_ana_0.dcomp3v3 por_ana_0.comparator_1.n1.t7 avss.t23 avss.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X806 por_dig_0.clknet_0_osc_ck.t11 a_34387_32909# dvss.t157 dvss.t156 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X807 a_30260_13935# a_29882_6535# avss.t241 sky130_fd_pr__res_xhigh_po_1p41 l=35
X808 dvdd.t1168 por_dig_0.cnt_por\[1\] por_dig_0._034_.t7 dvdd.t1167 sky130_fd_pr__pfet_01v8_hvt ad=0.42 pd=2.84 as=0.135 ps=1.27 w=1 l=0.15
X809 por_ana_0.rstring_mux_0.otrip_decoded_avdd[3] a_24673_24371# avdd.t454 avdd.t453 sky130_fd_pr__pfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.24375 ps=1.825 w=1.5 l=0.5
X810 avdd.t407 por_ana_0.comparator_1.vpp.t51 por_ana_0.comparator_1.vnn.t27 avdd.t401 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X811 dvss.t2061 a_38957_32883# por_dig_0._001_ dvss.t2060 sky130_fd_pr__nfet_01v8 ad=0.26 pd=1.45 as=0.17225 ps=1.83 w=0.65 l=0.15
X812 avdd.t134 avdd.t132 avdd.t133 avdd.t3 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=8
X813 por_ana_0.rc_osc_0.m por_ana_0.rc_osc_0.in dvdd.t241 dvdd.t240 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X814 dvss.t439 por_dig_0.net24 a_33518_35451# dvss.t438 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X815 a_25724_13935# por_ana_0.rstring_mux_0.vtrip0.t7 avss.t242 sky130_fd_pr__res_xhigh_po_1p41 l=35
X816 dvdd.t1614 dvss.t2267 dvdd.t1613 dvdd.t1612 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X817 a_34010_31821# a_33774_31821# dvss.t1090 dvss.t1089 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.5
X818 a_34654_32141# por_dig_0.cnt_por\[7\] a_34570_32141# dvss.t1096 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X819 dcomp.t26 por_ana_0.sky130_fd_sc_hd__inv_4_3.Y dvdd.t57 dvdd.t56 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X820 dvss.t2104 por_dig_0.net20.t3 a_34202_36717# dvss.t2103 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X821 a_35768_33690# a_35573_33721# a_36078_33453# dvss.t1978 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.1401 ps=1.1 w=0.36 l=0.15
X822 avdd.t198 por_ana_0.comparator_0.vpp.t8 por_ana_0.comparator_0.vpp.t9 avdd.t195 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X823 a_21622_21903# a_21254_22885# dvdd.t918 dvdd.t917 sky130_fd_pr__pfet_01v8_hvt ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X824 avdd.t131 avdd.t129 avdd.t130 avdd.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=8
X825 a_38499_34363# por_dig_0.net25 dvss.t959 dvss.t958 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X826 a_30495_23593# a_30070_23637# dvss.t1296 dvss.t1295 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X827 a_38974_34693# a_39070_34515# dvdd.t935 dvdd.t934 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14075 ps=1.325 w=0.42 l=0.5
X828 a_36406_23637# a_36038_24619# dvss.t683 dvss.t682 sky130_fd_pr__nfet_01v8 ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X829 por_ana_0.comparator_0.n1.t0 por_ana_0.comparator_0.n0.t5 avdd.t500 avdd.t499 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.6
X830 dvss.t1654 dvss.t1652 force_pdn.t0 dvss.t1653 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X831 a_21622_23637# a_21254_24619# dvdd.t920 dvdd.t919 sky130_fd_pr__pfet_01v8_hvt ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X832 dvss.t1877 dvdd.t1841 dvss.t1876 dvss.t1875 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X833 dvdd.t694 por_dig_0.por_unbuf.t9 a_25495_33620# dvdd.t693 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X834 dvss.t1874 dvdd.t1842 dvss.t1873 dvss.t1872 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X835 por_ana_0.rstring_mux_0.vtrip4.t5 por_ana_0.rstring_mux_0.otrip_decoded_b_avdd[4] vin.t40 avdd.t560 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X836 a_30495_23593# a_30070_23637# dvss.t1294 dvss.t1293 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X837 por_dig_0.clknet_1_0__leaf_osc_ck.t29 a_34098_30707# dvdd.t175 dvdd.t174 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X838 por_ana_0.ibias_gen_0.vp1.t7 por_ana_0.ibias_gen_0.vn1.t12 avss.t402 avss.t398 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=8
X839 dvss.t1871 dvdd.t1843 dvss.t1870 dvss.t1869 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X840 dvdd.t1296 por_dig_0._039_ por_dig_0._000_ dvdd.t1295 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X841 a_31894_32365# a_31728_32365# dvdd.t587 dvdd.t586 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X842 avss.t112 avss.t111 avss.t112 avss.t100 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=8
X843 dvdd.t1617 dvss.t2268 dvdd.t1616 dvdd.t1615 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X844 por_dig_0.cnt_por\[1\] a_37584_35389# dvdd.t881 dvdd.t880 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3012 ps=2.66 w=1 l=0.15
X845 a_31932_33595# por_dig_0.clknet_1_1__leaf_osc_ck.t33 dvss.t701 dvss.t700 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X846 avdd.t128 avdd.t127 avdd.t128 avdd.t13 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=8
X847 a_34467_28557# a_34290_28557# dvdd.t858 dvdd.t857 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X848 dvdd.t181 a_32088_31514# a_32019_31643# dvdd.t180 sky130_fd_pr__pfet_01v8_hvt ad=0.2184 pd=2.2 as=0.12915 ps=1.185 w=0.84 l=0.15
X849 avdd.t126 avdd.t124 avdd.t125 avdd.t3 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=8
X850 a_38053_30189# a_36972_30189# a_37706_30431# dvdd.t17 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X851 a_31914_24707# a_31814_24619# dvss.t2052 dvss.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X852 a_31876_32199# a_31360_31827# a_31781_32187# dvss.t31 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X853 avdd.t329 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.t13 porb_h.t12 avdd.t328 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X854 dvdd.t533 por_dig_0.cnt_por\[0\].t11 a_34672_35451# dvdd.t532 sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X855 dvdd.t173 a_34098_30707# por_dig_0.clknet_1_0__leaf_osc_ck.t28 dvdd.t172 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X856 dvdd.t1620 dvss.t2269 dvdd.t1619 dvdd.t1618 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X857 dvss.t292 por_ana_0.rc_osc_0.in por_ana_0.rc_osc_0.m dvss.t291 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X858 dvss.t110 a_38150_22885# a_38250_22973# dvss.t109 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X859 a_32094_31795# a_31876_32199# dvdd.t1510 dvdd.t1509 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X860 dvss.t1651 dvss.t1649 osc_ck.t1 dvss.t1650 sky130_fd_pr__nfet_01v8 ad=0.1475 pd=1.295 as=0.15 ps=1.3 w=1 l=0.18
X861 dvss.t11 a_32182_23637# a_32607_23593# dvss.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X862 dvdd.t1365 por_dig_0.otrip_decoded[2].t4 a_23366_22885# dvdd.t1364 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X863 avdd.t253 a_38250_22973# a_39457_22637# avdd.t252 sky130_fd_pr__pfet_g5v0d10v5 ad=0.24375 pd=1.825 as=0.3975 ps=3.53 w=1.5 l=0.5
X864 por_ana_0.rstring_mux_0.vtrip_decoded_b_avdd[0] por_ana_0.rstring_mux_0.vtrip_decoded_avdd[0] avdd.t424 avdd.t423 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X865 dvdd.t1622 dvss.t2270 dvdd.t1621 dvdd.t1522 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X866 dvdd.t1625 dvss.t2271 dvdd.t1624 dvdd.t1623 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X867 avdd.t408 por_ana_0.comparator_1.vpp.t52 por_ana_0.comparator_1.vnn.t26 avdd.t401 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X868 avss.t339 por_ana_0.ibias_gen_0.isrc_sel.t4 por_ana_0.ibias_gen_0.isrc_sel_b.t3 avss.t338 sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=1
X869 dvdd.t1433 por_dig_0.otrip_decoded[3].t4 a_23366_24619# dvdd.t1432 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X870 por_ana_0.comparator_1.vt.t51 vbg_1v2.t12 por_ana_0.comparator_1.vnn por_ana_0.comparator_1.vt.t41 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X871 dvdd.t1627 dvss.t2272 dvdd.t1626 dvdd.t1612 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X872 por_dig_0._047_ a_33600_34335# dvdd.t377 dvdd.t376 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X873 dvdd.t521 a_37961_33453# a_38136_33427# dvdd.t520 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X874 por_dig_0._037_ por_dig_0.cnt_por\[9\] dvdd.t1501 dvdd.t1500 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.165 ps=1.33 w=1 l=0.15
X875 dvss.t1106 a_21622_21903# a_22047_21859# dvss.t1105 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X876 avdd.t308 a_36138_24707# a_36831_23593# avdd.t307 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.1365 ps=1.49 w=0.42 l=1
X877 otrip[0].t0 dvss.t1646 dvss.t1648 dvss.t1647 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X878 a_13894_21948# por_ana_0.ibias_gen_0.isrc_sel.t5 por_ana_0.ibias_gen_0.vn1.t9 avss.t340 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X879 dvdd.t318 a_35293_30189# a_35468_30163# dvdd.t317 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X880 a_34946_30431# a_34728_30189# dvss.t1353 dvss.t1352 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X881 dvss.t1868 dvdd.t1844 dvss.t1867 dvss.t1866 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X882 porb.t15 por_ana_0.sky130_fd_sc_hd__inv_4_1.Y dvss.t355 dvss.t354 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X883 a_38307_33997# a_37230_34003# a_38145_34375# dvdd.t915 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X884 dvss.t437 por_dig_0.net24 a_33242_33275# dvss.t436 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X885 por_ana_0.schmitt_trigger_0.out.t0 por_ana_0.schmitt_trigger_0.m.t15 dvss.t649 dvss.t648 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X886 por_dig_0.net24 a_35100_32339# dvdd.t1048 dvdd.t1047 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X887 a_34719_23593# a_34294_23637# dvss.t1345 dvss.t1344 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X888 por_dig_0.clknet_0_osc_ck.t28 a_34387_32909# dvdd.t127 dvdd.t126 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X889 dvss.t2145 a_36100_32517# por_dig_0._019_ dvss.t2144 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X890 a_23456_13935# a_23078_6535# avss.t223 sky130_fd_pr__res_xhigh_po_1p41 l=35
X891 a_32244_32365# a_31894_32365# a_32149_32365# dvdd.t1312 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X892 a_38518_23637# a_38150_24619# dvss.t45 dvss.t44 sky130_fd_pr__nfet_01v8 ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X893 porb_h.t11 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.t14 avdd.t331 avdd.t330 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X894 dvss.t592 a_35583_34541# por_dig_0.clknet_1_1__leaf_osc_ck.t13 dvss.t591 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X895 a_38500_31251# por_dig_0.cnt_st\[4\] dvss.t1529 dvss.t1528 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X896 dvss.t590 a_35583_34541# por_dig_0.clknet_1_1__leaf_osc_ck.t12 dvss.t589 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X897 dvdd.t885 a_36380_33971# por_dig_0.net22.t2 dvdd.t884 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X898 por_ana_0.comparator_0.vnn.t24 por_ana_0.comparator_0.vinn.t51 por_ana_0.comparator_0.vt.t14 por_ana_0.comparator_0.vt.t3 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X899 avdd.t409 por_ana_0.comparator_1.vpp.t53 por_ana_0.comparator_1.vnn.t25 avdd.t401 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X900 dvss.t200 a_34098_30707# por_dig_0.clknet_1_0__leaf_osc_ck.t10 dvss.t199 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X901 a_24212_13935# a_24590_6535# avss.t224 sky130_fd_pr__res_xhigh_po_1p41 l=35
X902 dvss.t1865 dvdd.t1845 dvss.t1864 dvss.t1863 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X903 a_37396_33287# a_37046_32915# a_37301_33275# dvdd.t436 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X904 dvss.t1645 dvss.t1643 isrc_sel.t1 dvss.t1644 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X905 avdd.t197 por_ana_0.comparator_0.vpp.t53 por_ana_0.comparator_0.vnn.t9 avdd.t180 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X906 dvdd.t798 a_31592_30965# por_dig_0._038_ dvdd.t797 sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.275 ps=2.55 w=1 l=0.15
X907 por_ana_0.comparator_1.vm.t3 por_ana_0.comparator_1.vm.t2 avss.t344 avss.t288 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X908 dvss.t176 por_dig_0._031_ a_39022_32159# dvss.t175 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X909 a_36467_31643# a_35390_31277# a_36305_31277# dvdd.t802 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X910 dvss.t1862 dvdd.t1846 dvss.t1861 dvss.t1860 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X911 por_ana_0.comparator_0.vt.t49 vbg_1v2.t13 por_ana_0.comparator_0.vpp.t20 por_ana_0.comparator_0.vt.t36 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X912 por_ana_0.comparator_0.vnn.t25 por_ana_0.comparator_0.vinn.t52 por_ana_0.comparator_0.vt.t13 por_ana_0.comparator_0.vt.t3 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X913 a_36100_32517# por_dig_0.cnt_por\[5\] dvdd.t1403 dvdd.t1402 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X914 por_ana_0.ibias_gen_0.vr.t1 avss.t110 por_ana_0.ibias_gen_0.ve.t2 avss.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X915 a_36607_28917# por_dig_0.net5.t4 a_36526_28917# dvss.t2113 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.05355 ps=0.675 w=0.42 l=0.15
X916 dvdd.t1630 dvss.t2273 dvdd.t1629 dvdd.t1628 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X917 a_22047_21859# a_21622_21903# dvss.t1104 dvss.t1103 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X918 a_34026_24707# a_33926_24619# dvss.t513 dvss.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X919 a_32616_32125# por_dig_0.net8 dvdd.t1180 dvdd.t1179 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X920 avss.t297 por_ana_0.comparator_0.n0.t6 por_ana_0.comparator_0.n1.t1 avss.t296 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X921 por_ana_0.comparator_0.vt.t48 vbg_1v2.t14 por_ana_0.comparator_0.vpp.t21 por_ana_0.comparator_0.vt.t36 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X922 a_32701_28531# por_dig_0.net12 dvss.t474 dvss.t473 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X923 dvdd.t1633 dvss.t2274 dvdd.t1632 dvdd.t1631 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X924 a_33940_31277# por_dig_0._036_.t4 dvss.t2016 dvss.t2015 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.105625 ps=0.975 w=0.65 l=0.15
X925 dvss.t1580 por_dig_0.cnt_por\[2\] a_34580_35629# dvss.t1579 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X926 dvss.t1343 a_34294_23637# a_34719_23593# dvss.t1342 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X927 por_dig_0._014_ a_33852_29645# a_34102_29645# dvdd.t70 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.26 ps=2.52 w=1 l=0.15
X928 avdd.t123 avdd.t121 avdd.t122 avdd.t3 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=8
X929 a_32088_33690# a_31932_33595# a_32233_33819# dvdd.t1416 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.1155 ps=0.97 w=0.42 l=0.15
X930 dvdd.t55 por_ana_0.sky130_fd_sc_hd__inv_4_3.Y dcomp.t25 dvdd.t54 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X931 por_ana_0.rstring_mux_0.vtrip_decoded_b_avdd[1] por_ana_0.rstring_mux_0.vtrip_decoded_avdd[1] avdd.t519 avdd.t518 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X932 dvdd.t591 por_dig_0.clknet_1_1__leaf_osc_ck.t34 a_37064_34003# dvdd.t590 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X933 dvss.t889 osc_ck.t11 a_34387_32909# dvss.t888 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X934 a_33256_35463# a_32906_35091# a_33161_35451# dvdd.t1018 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X935 dvss.t155 a_34387_32909# por_dig_0.clknet_0_osc_ck.t10 dvss.t154 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X936 a_38956_32339# por_dig_0.cnt_st\[1\] a_39354_32365# dvss.t601 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0609 ps=0.71 w=0.42 l=0.15
X937 dvss.t501 por_dig_0.clknet_1_0__leaf_osc_ck.t38 a_36972_30189# dvss.t500 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X938 a_34580_35629# por_dig_0.cnt_por\[3\] a_34830_35629# dvss.t453 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X939 dvss.t2018 por_dig_0._036_.t5 a_35433_32141# dvss.t2017 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.19825 ps=1.26 w=0.65 l=0.15
X940 a_31894_32365# a_31728_32365# dvss.t694 dvss.t693 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X941 por_dig_0.osc_ena.t2 a_31413_29619# dvdd.t1398 dvdd.t70 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X942 dvss.t1413 a_23734_21903# a_24159_21859# dvss.t1412 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X943 dvss.t1059 a_35556_29619# a_35298_29619# dvss.t1058 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.5
X944 dvdd.t1636 dvss.t2275 dvdd.t1635 dvdd.t1634 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X945 dcomp.t24 por_ana_0.sky130_fd_sc_hd__inv_4_3.Y dvdd.t53 dvdd.t52 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X946 avdd.t442 a_38250_24707# a_38943_23593# avdd.t441 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.1365 ps=1.49 w=0.42 l=1
X947 dvss.t681 a_36038_24619# a_36138_24707# dvss.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X948 dvdd.t531 pwup_filt.t33 a_32004_30189# dvdd.t530 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X949 a_35583_34541# por_dig_0.clknet_0_osc_ck.t36 dvdd.t1455 dvdd.t1454 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X950 dvss.t1204 por_dig_0._049_ a_36328_36493# dvss.t1203 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X951 avdd.t482 por_ana_0.comparator_0.n1.t8 por_ana_0.dcomp3v3uv avdd.t481 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.6
X952 a_34633_36147# por_dig_0.cnt_por\[2\] a_34762_36173# dvdd.t1271 sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X953 a_35040_34317# por_dig_0._023_ dvss.t928 dvss.t927 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X954 a_31984_31821# por_dig_0.net8 dvdd.t1178 dvdd.t1177 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X955 a_4811_22912# a_5189_15512# avss.t27 sky130_fd_pr__res_xhigh_po_1p41 l=35
X956 dvss.t1423 por_dig_0.net8 a_32138_32187# dvss.t1422 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X957 dvdd.t807 a_32809_32365# a_32984_32339# dvdd.t806 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X958 por_dig_0._034_.t6 por_dig_0.cnt_por\[1\] dvdd.t1166 dvdd.t1165 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.335 ps=1.67 w=1 l=0.15
X959 a_37798_33971# a_37580_34375# dvss.t1274 dvss.t1273 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X960 dvdd.t563 por_ana_0.schmitt_trigger_0.in.t5 por_ana_0.schmitt_trigger_0.m.t5 dvdd.t562 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X961 avdd.t547 por_ana_0.comparator_1.n0.t7 por_ana_0.comparator_1.n1.t0 avdd.t546 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X962 a_38254_34375# a_37064_34003# a_38145_34375# dvss.t1272 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X963 a_13844_23626# por_ana_0.ibias_gen_0.isrc_sel_b.t4 por_ana_0.ibias_gen_0.vn1.t7 avdd.t575 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X964 por_dig_0.net7.t0 a_34615_28013# dvss.t1109 dvss.t523 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X965 dvdd.t1137 a_37961_33287# a_38136_33213# dvdd.t1136 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X966 dvss.t318 por_dig_0.cnt_por\[8\] a_33774_31821# dvss.t317 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X967 dvdd.t1335 por_dig_0._053_ a_33380_35879# dvdd.t1334 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X968 dvdd.t51 por_ana_0.sky130_fd_sc_hd__inv_4_3.Y dcomp.t23 dvdd.t50 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X969 dvss.t401 a_39887_23089# a_40246_23089# dvss.t400 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.19875 ps=2.03 w=0.75 l=0.5
X970 dvss.t1859 dvdd.t1847 dvss.t1858 dvss.t1847 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X971 porb_h.t10 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.t15 avdd.t333 avdd.t332 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X972 a_38352_32365# por_dig_0.cnt_st\[0\] dvdd.t1114 dvdd.t1113 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X973 pwup_filt.t14 por_ana_0.sky130_fd_sc_hd__inv_4_0.Y dvss.t256 dvss.t255 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X974 dvss.t1857 dvdd.t1848 dvss.t1856 dvss.t1794 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X975 dvdd.t215 por_ana_0.sky130_fd_sc_hd__inv_4_0.Y pwup_filt.t26 dvdd.t214 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X976 a_17408_13935# a_17786_6535# avss.t174 sky130_fd_pr__res_xhigh_po_1p41 l=35
X977 dvss.t1455 a_37952_31037# a_37886_31111# dvss.t1454 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X978 a_36234_35871# a_36016_35629# dvdd.t822 dvdd.t821 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X979 dvdd.t1102 force_pdn.t2 a_31360_28557# dvdd.t1101 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X980 a_20432_13935# a_20810_6535# avss.t175 sky130_fd_pr__res_xhigh_po_1p41 l=35
X981 a_35674_28557# por_dig_0.net7.t6 dvss.t851 dvss.t850 sky130_fd_pr__nfet_01v8 ad=0.10785 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X982 dvdd.t1373 por_dig_0.cnt_st\[2\] a_38352_32365# dvdd.t1372 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X983 dvss.t169 a_34746_31277# a_34852_31277# dvss.t168 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.5
X984 avdd.t410 por_ana_0.comparator_1.vpp.t54 por_ana_0.comparator_1.vnn.t24 avdd.t401 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X985 dvss.t2084 a_34357_33427# por_dig_0._021_ dvss.t886 sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.17225 ps=1.83 w=0.65 l=0.15
X986 a_7079_22912# a_7457_15512# avss.t27 sky130_fd_pr__res_xhigh_po_1p41 l=35
X987 dvss.t254 por_ana_0.sky130_fd_sc_hd__inv_4_0.Y pwup_filt.t13 dvss.t253 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X988 por_dig_0.net14 a_35774_28673# dvdd.t633 dvdd.t632 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X989 dvss.t853 por_dig_0.net7.t7 a_35289_28917# dvss.t852 sky130_fd_pr__nfet_01v8 ad=0.122275 pd=1.08 as=0.05355 ps=0.675 w=0.42 l=0.15
X990 dvss.t976 a_36406_23637# a_36831_23593# dvss.t975 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X991 por_dig_0._048_ por_dig_0.net4 a_35954_34317# dvss.t97 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X992 por.t30 por_ana_0.sky130_fd_sc_hd__inv_4_4.Y dvdd.t976 dvdd.t975 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X993 dvdd.t1639 dvss.t2276 dvdd.t1638 dvdd.t1637 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X994 dvdd.t637 a_33821_35463# a_33996_35389# dvdd.t636 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X995 otrip[2].t1 dvss.t1640 dvss.t1642 dvss.t1641 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X996 a_35690_33997# por_dig_0._018_ por_dig_0._009_ dvdd.t457 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.174 ps=1.39 w=1 l=0.15
X997 por_ana_0.rstring_mux_0.otrip_decoded_avdd[0] a_22561_22637# dvss.t740 dvss.t739 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.121875 ps=1.075 w=0.75 l=0.5
X998 a_36756_35603# a_36581_35629# a_36935_35629# dvss.t2208 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X999 dvss.t1002 a_25846_21903# a_26271_21859# dvss.t1001 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X1000 dvdd.t171 a_34098_30707# por_dig_0.clknet_1_0__leaf_osc_ck.t27 dvdd.t170 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1001 a_34024_33703# por_dig_0._021_ dvdd.t631 dvdd.t630 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X1002 por_ana_0.comparator_0.vt.t12 por_ana_0.comparator_0.vinn.t53 por_ana_0.comparator_0.vnn por_ana_0.comparator_0.vt.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1003 dvss.t43 a_38150_24619# a_38250_24707# dvss.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X1004 dvss.t1503 por_dig_0._011_ a_32651_33819# dvss.t1502 sky130_fd_pr__nfet_01v8 ad=0.2205 pd=1.89 as=0.066 ps=0.745 w=0.42 l=0.15
X1005 por_dig_0.net6 a_33971_28557# dvss.t1387 dvss.t1386 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X1006 avdd.t335 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.t16 porb_h.t9 avdd.t334 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X1007 dvss.t1855 dvdd.t1849 dvss.t1854 dvss.t1853 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1008 por_ana_0.rstring_mux_0.vtop.t17 a_13250_6535# avss.t176 sky130_fd_pr__res_xhigh_po_1p41 l=35
X1009 porb.t23 por_ana_0.sky130_fd_sc_hd__inv_4_1.Y dvdd.t287 dvdd.t286 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1010 a_33720_33213# a_33545_33287# a_33899_33275# dvss.t741 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X1011 avdd.t363 por_ana_0.comparator_0.vnn.t48 por_ana_0.comparator_0.vpp.t32 avdd.t195 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1012 dvss.t2131 por_dig_0.clknet_0_osc_ck.t37 a_34098_30707# dvss.t2130 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X1013 a_37614_32883# a_37396_33287# dvss.t918 dvss.t917 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X1014 a_39152_32365# por_dig_0.cnt_st\[2\] dvss.t2033 dvss.t2032 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.196275 ps=1.33 w=0.42 l=0.15
X1015 porb.t14 por_ana_0.sky130_fd_sc_hd__inv_4_1.Y dvss.t353 dvss.t352 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1016 por.t4 por_ana_0.sky130_fd_sc_hd__inv_4_4.Y dvss.t1145 dvss.t1144 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1017 avdd.t196 por_ana_0.comparator_0.vpp.t6 por_ana_0.comparator_0.vpp.t7 avdd.t195 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1018 dvss.t1852 dvdd.t1850 dvss.t1851 dvss.t1850 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X1019 por_ana_0.dcomp3v3 por_ana_0.comparator_1.n1.t8 avdd.t535 avdd.t534 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X1020 a_36376_28789# a_36649_28789# a_36607_28917# dvss.t2069 sky130_fd_pr__nfet_01v8 ad=0.107825 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X1021 a_34750_28557# a_34573_28557# dvdd.t645 dvdd.t644 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X1022 a_37062_35059# a_36844_35463# dvdd.t647 dvdd.t646 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X1023 a_37301_33275# por_dig_0._002_ dvss.t1962 dvss.t1087 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X1024 a_35468_30163# por_dig_0.net25 dvdd.t842 dvdd.t841 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X1025 dvss.t1639 dvss.t1637 vin.t39 dvss.t1638 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X1026 por_dig_0._023_ a_34580_34110# dvdd.t1030 dvdd.t1029 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X1027 a_28383_21859# a_27958_21903# dvss.t2200 dvss.t2199 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X1028 dvdd.t1376 a_36476_30163# a_36218_30163# dvdd.t1375 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.5
X1029 dvss.t351 por_ana_0.sky130_fd_sc_hd__inv_4_1.Y porb.t13 dvss.t350 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1030 a_37396_33453# a_36880_33453# a_37301_33453# dvss.t522 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X1031 dvss.t1335 por_dig_0.cnt_st\[0\] a_39262_34317# dvss.t1334 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1032 por_dig_0.clknet_0_osc_ck.t27 a_34387_32909# dvdd.t125 dvdd.t124 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1033 dvdd.t1642 dvss.t2277 dvdd.t1641 dvdd.t1640 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1034 dvss.t588 a_35583_34541# por_dig_0.clknet_1_1__leaf_osc_ck.t11 dvss.t587 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1035 por_ana_0.rstring_mux_0.otrip_decoded_avdd[3] a_24673_24371# dvss.t1086 dvss.t1085 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.121875 ps=1.075 w=0.75 l=0.5
X1036 dvdd.t657 a_37156_28013# por_dig_0.otrip_decoded[7].t3 dvdd.t656 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X1037 a_36844_35463# a_36328_35091# a_36749_35451# dvss.t992 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X1038 a_40246_23089# a_39887_23089# dvss.t399 dvss.t396 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.105 ps=1.03 w=0.75 l=0.5
X1039 dvss.t1095 por_dig_0.cnt_por\[7\] a_33805_32339# dvss.t1094 sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.10725 ps=0.98 w=0.65 l=0.15
X1040 a_40247_24823# a_39888_24823# dvss.t761 dvss.t754 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.105 ps=1.03 w=0.75 l=0.5
X1041 dvdd.t1645 dvss.t2278 dvdd.t1644 dvdd.t1643 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X1042 por_ana_0.comparator_1.vt.t50 vbg_1v2.t15 por_ana_0.comparator_1.vnn por_ana_0.comparator_1.vt.t41 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1043 avss.t183 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.t17 porb_h.t29 avss.t182 sky130_fd_pr__nfet_g5v0d10v5 ad=0.2025 pd=2.04 as=0.105 ps=1.03 w=0.75 l=0.5
X1044 dvss.t1324 force_dis_rc_osc.t3 a_31360_33997# dvss.t1323 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X1045 dvss.t2217 a_38518_23637# a_38943_23593# dvss.t2216 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X1046 dvss.t1969 por_dig_0._043_ a_39813_31277# dvss.t1968 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X1047 por_ana_0.sky130_fd_sc_hd__inv_4_1.Y por_ana_0.sky130_fd_sc_hd__inv_4_1.A dvdd.t193 dvdd.t192 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1048 por_dig_0.net9 por_dig_0.net3 dvdd.t1127 dvdd.t1126 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1049 porb.t22 por_ana_0.sky130_fd_sc_hd__inv_4_1.Y dvdd.t285 dvdd.t284 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1050 por_ana_0.comparator_1.vt.t49 vbg_1v2.t16 por_ana_0.comparator_1.vnn por_ana_0.comparator_1.vt.t41 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1051 por_ana_0.rstring_mux_0.otrip_decoded_avdd[4] a_26785_22637# dvss.t763 dvss.t762 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.121875 ps=1.075 w=0.75 l=0.5
X1052 por_dig_0.clknet_1_1__leaf_osc_ck.t24 a_35583_34541# dvdd.t487 dvdd.t486 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1053 a_33852_29645# por_dig_0._027_ dvss.t1049 dvss.t1048 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1054 por_ana_0.schmitt_trigger_0.in.t6 dvss.t654 sky130_fd_pr__cap_mim_m3_2 l=30 w=30
X1055 a_38145_34375# a_37230_34003# a_37798_33971# dvss.t1056 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X1056 a_34114_35879# por_dig_0.net20.t4 dvdd.t1425 dvdd.t1265 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.165 ps=1.33 w=1 l=0.15
X1057 a_34836_30555# por_dig_0.net25 dvdd.t840 dvdd.t158 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X1058 vin.t19 avss.t108 vin.t19 avss.t109 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=0.6
X1059 avdd.t318 a_27690_24707# a_28897_24371# avdd.t317 sky130_fd_pr__pfet_g5v0d10v5 ad=0.24375 pd=1.825 as=0.3975 ps=3.53 w=1.5 l=0.5
X1060 avdd.t281 por_ana_0.sky130_fd_sc_hvl__inv_4_0.A por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.t3 avdd.t280 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.21 ps=1.78 w=1.5 l=0.5
X1061 a_4055_22912# a_3677_15512# avss.t27 sky130_fd_pr__res_xhigh_po_1p41 l=35
X1062 por_ana_0.comparator_0.vinn.t42 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[4].t3 por_ana_0.rstring_mux_0.vtrip4.t2 avss.t327 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X1063 dvdd.t283 por_ana_0.sky130_fd_sc_hd__inv_4_1.Y porb.t21 dvdd.t282 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1064 avdd.t237 por_ana_0.rstring_mux_0.ena_b por_ana_0.rstring_mux_0.vtop.t9 avdd.t236 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X1065 por_ana_0.comparator_0.vpp.t22 vbg_1v2.t17 por_ana_0.comparator_0.vt.t47 por_ana_0.comparator_0.vt.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1066 dvss.t1636 dvss.t1634 otrip[1].t0 dvss.t1635 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X1067 dvss.t891 osc_ck.t12 a_34387_32909# dvss.t890 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1068 dvdd.t1264 a_35640_32517# por_dig_0._017_ dvdd.t1263 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.26 ps=2.52 w=1 l=0.15
X1069 por_ana_0.ibias_gen_0.vn0.t10 vbg_1v2.t18 por_ana_0.ibias_gen_0.vstart.t5 avss.t153 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X1070 dvdd.t661 por_dig_0.net18 a_37156_28013# dvdd.t660 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X1071 por_ana_0.comparator_1.vnn.t7 por_ana_0.comparator_1.vnn.t6 avdd.t628 avdd.t403 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1072 por_dig_0._039_ por_dig_0.net4 dvss.t96 dvss.t95 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1073 dcomp.t22 por_ana_0.sky130_fd_sc_hd__inv_4_3.Y dvdd.t49 dvdd.t48 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1074 a_33444_31037# a_33269_31111# a_33623_31099# dvss.t1051 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X1075 dvss.t252 por_ana_0.sky130_fd_sc_hd__inv_4_0.Y pwup_filt.t12 dvss.t251 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1076 dvss.t63 por_ana_0.sky130_fd_sc_hd__inv_4_3.Y dcomp.t7 dvss.t62 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1077 dvss.t1849 dvdd.t1851 dvss.t1848 dvss.t1847 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1078 a_37584_35389# por_dig_0.net24 dvdd.t349 dvdd.t348 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X1079 por_ana_0.ibias_gen_0.vp.t0 avdd.t119 por_ana_0.ibias_gen_0.vp.t0 avdd.t120 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=0.6
X1080 a_37393_30189# por_dig_0._003_ dvss.t772 dvss.t771 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X1081 dvdd.t665 por_dig_0._051_ a_32828_35879# dvdd.t664 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X1082 avss.t107 avss.t105 avss.t106 avss.t81 sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0 ps=0 w=5 l=8
X1083 dvdd.t47 por_ana_0.sky130_fd_sc_hd__inv_4_3.Y dcomp.t21 dvdd.t46 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1084 por_ana_0.comparator_0.vn.t0 avss.t103 por_ana_0.comparator_0.ibias.t0 avss.t104 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X1085 dvdd.t1648 dvss.t2279 dvdd.t1647 dvdd.t1646 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1086 dvss.t1092 a_34010_31821# a_34116_31821# dvss.t1091 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.5
X1087 por_ana_0.rc_osc_0.n.t1 por_ana_0.rc_osc_0.m dvdd.t444 dvdd.t443 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X1088 a_6323_22912# a_5945_15512# avss.t27 sky130_fd_pr__res_xhigh_po_1p41 l=35
X1089 a_34828_29253# por_dig_0.net7.t8 dvdd.t738 dvdd.t737 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14575 ps=1.335 w=0.42 l=0.15
X1090 dvss.t1569 a_33996_36477# a_33930_36551# dvss.t1568 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X1091 por_ana_0.sky130_fd_sc_hd__inv_4_0.Y por_ana_0.schmitt_trigger_0.out.t8 dvdd.t710 dvdd.t709 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1092 dvdd.t1651 dvss.t2280 dvdd.t1650 dvdd.t1649 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1093 avdd.t364 por_ana_0.comparator_0.vnn.t49 por_ana_0.comparator_0.vpp.t33 avdd.t195 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1094 a_37820_13935# a_37442_6535# avss.t177 sky130_fd_pr__res_xhigh_po_1p41 l=35
X1095 a_23466_22973# a_23366_22885# dvss.t912 dvss.t911 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X1096 a_32922_30707# a_32704_31111# dvdd.t820 dvdd.t819 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X1097 a_34828_29253# por_dig_0.net7.t9 dvss.t855 dvss.t854 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.10025 ps=0.985 w=0.42 l=0.15
X1098 avss.t102 avss.t99 avss.t101 avss.t100 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=8
X1099 por_ana_0.schmitt_trigger_0.in.t7 dvss.t655 sky130_fd_pr__cap_mim_m3_2 l=30 w=30
X1100 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.t2 por_ana_0.sky130_fd_sc_hvl__inv_4_0.A avdd.t279 avdd.t278 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X1101 a_33284_13935# a_32906_6535# avss.t311 sky130_fd_pr__res_xhigh_po_1p41 l=35
X1102 vin.t7 avdd.t117 vin.t7 avdd.t118 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=0.6
X1103 por_ana_0.comparator_0.vinn.t33 por_ana_0.rstring_mux_0.vtrip_decoded_b_avdd[4] por_ana_0.rstring_mux_0.vtrip4.t4 avdd.t471 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X1104 dvss.t770 por_dig_0.net18 a_37156_28013# dvss.t677 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X1105 dvdd.t712 por_ana_0.schmitt_trigger_0.out.t9 por_ana_0.sky130_fd_sc_hd__inv_4_0.Y dvdd.t711 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1106 dvdd.t659 por_dig_0._017_ a_35690_33997# dvdd.t658 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1107 a_34672_35451# por_dig_0.cnt_por\[1\] dvdd.t1164 dvdd.t1163 sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.1092 ps=1.36 w=0.42 l=0.15
X1108 dvss.t760 a_39888_24823# a_40247_24823# dvss.t759 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.19875 ps=2.03 w=0.75 l=0.5
X1109 por_ana_0.rstring_mux_0.vtrip7.t6 a_29126_6535# avss.t312 sky130_fd_pr__res_xhigh_po_1p41 l=35
X1110 a_36500_33229# por_dig_0._033_ por_dig_0._018_ dvss.t35 sky130_fd_pr__nfet_01v8 ad=0.095875 pd=0.945 as=0.091 ps=0.93 w=0.65 l=0.15
X1111 dvss.t435 por_dig_0.net24 a_36278_35629# dvss.t434 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X1112 a_37485_34363# por_dig_0._000_ dvdd.t782 dvdd.t781 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X1113 vin.t43 por_ana_0.rstring_mux_0.otrip_decoded_avdd[6] por_ana_0.rstring_mux_0.vtrip6.t7 avss.t374 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X1114 por_ana_0.rstring_mux_0.otrip_decoded_avdd[6] a_28897_22637# dvss.t1989 dvss.t1988 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.121875 ps=1.075 w=0.75 l=0.5
X1115 a_34982_29351# por_dig_0.net5.t5 a_34898_29351# dvdd.t668 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1116 dvss.t250 por_ana_0.sky130_fd_sc_hd__inv_4_0.Y pwup_filt.t11 dvss.t249 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1117 a_36331_33819# a_35612_33595# a_35768_33690# dvss.t1471 sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0594 ps=0.69 w=0.36 l=0.15
X1118 a_36414_32909# por_dig_0.cnt_por\[4\] por_dig_0._018_ dvdd.t1254 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X1119 dvss.t967 a_33752_28013# por_dig_0.otrip_decoded[2].t1 dvss.t523 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X1120 a_35130_28673# por_dig_0.net6 dvdd.t678 dvdd.t677 sky130_fd_pr__pfet_01v8_hvt ad=0.074375 pd=0.815 as=0.0567 ps=0.69 w=0.42 l=0.15
X1121 a_35770_29351# por_dig_0.net6 a_35686_29351# dvdd.t668 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1122 dvss.t1430 a_21354_22973# a_22561_22637# dvss.t1429 sky130_fd_pr__nfet_g5v0d10v5 ad=0.121875 pd=1.075 as=0.19875 ps=2.03 w=0.75 l=0.5
X1123 a_31650_31277# a_31615_31529# a_31412_31251# dvss.t1283 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.1092 ps=1.36 w=0.42 l=0.15
X1124 avdd.t289 a_34026_24707# a_34719_23593# avdd.t288 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.1365 ps=1.49 w=0.42 l=1
X1125 dvss.t1846 dvdd.t1852 dvss.t1845 dvss.t1844 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X1126 a_38974_34693# a_39070_34515# dvss.t1108 dvss.t1107 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.5
X1127 dvss.t1633 dvss.t1631 a_36038_22885# dvss.t1632 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X1128 dvss.t1268 a_33996_35389# a_33930_35463# dvss.t1267 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X1129 por_ana_0.comparator_0.vpp.t23 vbg_1v2.t19 por_ana_0.comparator_0.vt.t46 por_ana_0.comparator_0.vt.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1130 dvss.t1432 a_31802_32909# a_31908_32909# dvss.t1431 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.5
X1131 dvdd.t459 a_32794_33971# por_dig_0._012_ dvdd.t458 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1132 a_35645_31277# por_dig_0._015_ dvdd.t312 dvdd.t311 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X1133 dvdd.t593 por_dig_0.clknet_1_1__leaf_osc_ck.t35 a_36880_33453# dvdd.t592 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1134 a_37698_31821# por_dig_0.cnt_st\[4\] dvdd.t1246 dvdd.t1245 sky130_fd_pr__pfet_01v8_hvt ad=0.1525 pd=1.305 as=0.26 ps=2.52 w=1 l=0.15
X1135 dvdd.t1654 dvss.t2281 dvdd.t1653 dvdd.t1652 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1136 a_35858_28013# por_dig_0.net7.t10 a_35776_28013# dvss.t677 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X1137 a_36122_30341# a_36218_30163# dvdd.t1378 dvdd.t1377 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14075 ps=1.325 w=0.42 l=0.5
X1138 dvdd.t1331 por_dig_0._026_ a_34444_32517# dvdd.t1330 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.135 ps=1.27 w=1 l=0.15
X1139 a_31972_32199# a_31526_31827# a_31876_32199# dvss.t1135 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X1140 dvdd.t1220 a_35960_29101# por_dig_0.otrip_decoded[6].t3 dvdd.t668 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X1141 por_ana_0.ibias_gen_0.vn1.t1 avss.t97 por_ana_0.ibias_gen_0.vp1.t1 avss.t98 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X1142 por_ana_0.sky130_fd_sc_hd__inv_4_4.Y por_dig_0.por_unbuf.t10 dvss.t802 dvss.t801 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1143 a_37777_31111# a_36696_30739# a_37430_30707# dvdd.t1065 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X1144 por.t3 por_ana_0.sky130_fd_sc_hd__inv_4_4.Y dvss.t1143 dvss.t1142 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1145 a_36138_22973# a_36038_22885# dvss.t276 dvss.t275 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X1146 avdd.t511 a_21354_22973# a_22047_21859# avdd.t510 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.1365 ps=1.49 w=0.42 l=1
X1147 dvss.t1438 a_34496_29645# por_dig_0._015_ dvss.t1437 sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.25025 ps=1.42 w=0.65 l=0.15
X1148 dvss.t198 a_34098_30707# por_dig_0.clknet_1_0__leaf_osc_ck.t9 dvss.t197 sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X1149 por_dig_0._003_ a_39077_31527# dvdd.t1192 dvdd.t1191 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.3275 ps=1.655 w=1 l=0.15
X1150 dvss.t1843 dvdd.t1853 dvss.t1842 dvss.t1841 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X1151 vin.t45 por_ana_0.rstring_mux_0.otrip_decoded_b_avdd[6] por_ana_0.rstring_mux_0.vtrip6.t9 avdd.t595 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X1152 dvdd.t281 por_ana_0.sky130_fd_sc_hd__inv_4_1.Y porb.t20 dvdd.t280 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1153 por_ana_0.comparator_1.vnn.t5 por_ana_0.comparator_1.vnn.t4 avdd.t627 avdd.t403 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1154 por_dig_0._046_ a_35040_34587# a_35219_34541# dvss.t985 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1155 dvdd.t1657 dvss.t2282 dvdd.t1656 dvdd.t1655 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1156 avdd.t116 avdd.t114 avdd.t116 avdd.t115 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=4
X1157 dvss.t1141 por_ana_0.sky130_fd_sc_hd__inv_4_4.Y por.t2 dvss.t1140 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1158 por_ana_0.ibias_gen_0.vn1.t8 por_ana_0.ibias_gen_0.isrc_sel_b.t5 avss.t336 avss.t335 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=2
X1159 dvss.t1630 dvss.t1628 vbg_1v2.t0 dvss.t1629 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X1160 dvdd.t635 por_dig_0.net14 a_37800_28013# dvdd.t634 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X1161 dvdd.t1660 dvss.t2283 dvdd.t1659 dvdd.t1658 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X1162 avss.t326 por_ana_0.ibias_gen_0.ena_b.t7 por_ana_0.ibias_gen_0.vn1.t6 avss.t325 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X1163 dvdd.t485 a_35583_34541# por_dig_0.clknet_1_1__leaf_osc_ck.t23 dvdd.t484 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1164 dvss.t1840 dvdd.t1854 dvss.t1839 dvss.t1838 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X1165 avdd.t337 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.t18 porb_h.t8 avdd.t336 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X1166 dvss.t108 a_38150_22885# a_38250_22973# dvss.t107 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X1167 por_dig_0.cnt_st\[3\] a_38228_30163# dvdd.t257 dvdd.t256 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X1168 avdd.t438 a_26271_21859# a_25578_22973# avdd.t437 sky130_fd_pr__pfet_g5v0d10v5 ad=0.2142 pd=1.99 as=0.2142 ps=1.99 w=0.42 l=1
X1169 a_18910_35244# a_19288_27844# avss.t313 sky130_fd_pr__res_xhigh_po_1p41 l=35
X1170 a_39888_24823# por_ana_0.dcomp3v3 avdd.t472 avdd.t311 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.1197 ps=1.41 w=0.42 l=0.5
X1171 a_37396_33287# a_36880_32915# a_37301_33275# dvss.t522 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X1172 por_ana_0.comparator_0.vinn.t9 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[3] por_ana_0.rstring_mux_0.vtrip3.t1 avss.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X1173 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[0] a_31009_22637# avdd.t649 avdd.t284 sky130_fd_pr__pfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.24375 ps=1.825 w=1.5 l=0.5
X1174 dvdd.t517 por_dig_0._009_ a_36331_33819# dvdd.t516 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X1175 dvss.t153 a_34387_32909# por_dig_0.clknet_0_osc_ck.t9 dvss.t152 sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X1176 avss.t96 avss.t95 avss.t96 avss.t45 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=8
X1177 dvdd.t619 por_dig_0.net17 a_35960_29101# dvdd.t618 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X1178 por_ana_0.rc_osc_0.m por_ana_0.rc_osc_0.n.t7 dvdd.t1353 dvdd.t1352 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1179 dvss.t2059 a_23466_22973# a_24673_22637# dvss.t2058 sky130_fd_pr__nfet_g5v0d10v5 ad=0.121875 pd=1.075 as=0.19875 ps=2.03 w=0.75 l=0.5
X1180 dvss.t1627 dvss.t1625 force_short_oneshot.t0 dvss.t1626 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X1181 dvss.t703 por_dig_0.clknet_1_1__leaf_osc_ck.t36 a_36880_32915# dvss.t702 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1182 osc_ck.t3 por_ana_0.rc_osc_0.n.t8 dvdd.t1355 dvdd.t1354 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X1183 a_33256_36551# a_32740_36179# a_33161_36539# dvss.t447 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X1184 dvss.t1102 a_21622_21903# a_22047_21859# dvss.t1101 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X1185 por_ana_0.dcomp3v3 por_ana_0.comparator_1.n1.t9 avss.t21 avss.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X1186 dvss.t926 a_34633_36147# por_dig_0._052_ dvss.t925 sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.17225 ps=1.83 w=0.65 l=0.15
X1187 dvss.t899 a_34467_28557# a_34573_28557# dvss.t898 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X1188 avdd.t113 avdd.t112 avdd.t113 avdd.t33 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=8
X1189 por_ana_0.sky130_fd_sc_hd__inv_4_3.Y por_ana_0.vl dvss.t1184 dvss.t1183 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1190 por_ana_0.comparator_0.vt.t11 por_ana_0.comparator_0.vinn.t54 por_ana_0.comparator_0.vnn por_ana_0.comparator_0.vt.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1191 dvss.t1837 dvdd.t1855 dvss.t1836 dvss.t1682 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1192 por_ana_0.comparator_0.vinn.t15 avss.t93 por_ana_0.comparator_0.vinn.t15 avss.t94 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=0.6
X1193 dvdd.t1663 dvss.t2284 dvdd.t1662 dvdd.t1661 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1194 por_dig_0.clknet_1_1__leaf_osc_ck.t22 a_35583_34541# dvdd.t483 dvdd.t482 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1195 avss.t92 avss.t90 avss.t91 avss.t81 sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0 ps=0 w=5 l=8
X1196 a_39887_23089# por_ana_0.dcomp3v3uv avdd.t290 avdd.t272 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.1197 ps=1.41 w=0.42 l=0.5
X1197 dvdd.t1304 a_37430_30707# a_37320_30733# dvdd.t1303 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X1198 dvss.t1835 dvdd.t1856 dvss.t1834 dvss.t1833 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X1199 por_dig_0._025_ por_dig_0._019_ dvdd.t1492 dvdd.t1491 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1200 avdd.t365 por_ana_0.comparator_0.vnn.t50 por_ana_0.comparator_0.vpp.t34 avdd.t195 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1201 dvss.t737 por_dig_0.net14 a_37800_28013# dvss.t677 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X1202 dvss.t1322 force_pdn.t3 a_31360_28557# dvss.t1321 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X1203 dvss.t1327 por_dig_0.otrip_decoded[0].t5 a_21254_22885# dvss.t1326 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X1204 a_35674_36539# por_dig_0.cnt_por\[1\] a_35592_36286# dvss.t1402 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X1205 por_ana_0.comparator_0.vt.t10 por_ana_0.comparator_0.vinn.t55 por_ana_0.comparator_0.vnn por_ana_0.comparator_0.vt.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1206 dvss.t1182 por_ana_0.vl por_ana_0.sky130_fd_sc_hd__inv_4_3.Y dvss.t1181 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1207 a_34946_30431# a_34728_30189# dvdd.t1123 dvdd.t1122 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X1208 dvss.t1997 a_33806_33427# por_dig_0._010_ dvss.t1996 sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X1209 porb_h.t7 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.t19 avdd.t339 avdd.t338 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X1210 a_35024_35629# por_dig_0.cnt_por\[0\].t12 a_34830_35629# dvss.t639 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1211 a_35092_33427# a_35295_33705# dvdd.t1151 dvdd.t1150 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1134 ps=1.38 w=0.42 l=0.15
X1212 dvss.t725 por_dig_0.net17 a_35960_29101# dvss.t724 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X1213 avss.t291 por_ana_0.comparator_1.vn.t5 por_ana_0.comparator_1.vn.t6 avss.t290 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1214 a_32019_33819# a_31932_33595# a_31615_33705# dvdd.t1415 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.0588 ps=0.7 w=0.42 l=0.15
X1215 por_ana_0.comparator_0.vinn.t11 por_ana_0.rstring_mux_0.vtrip_decoded_b_avdd[3] por_ana_0.rstring_mux_0.vtrip3.t3 avdd.t261 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X1216 pwup_filt.t10 por_ana_0.sky130_fd_sc_hd__inv_4_0.Y dvss.t248 dvss.t247 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1217 por_ana_0.ibias_gen_0.vn0.t11 vbg_1v2.t20 por_ana_0.ibias_gen_0.vstart.t4 avss.t152 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X1218 a_31651_30341# por_dig_0.net2 dvss.t178 dvss.t177 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.10025 ps=0.985 w=0.42 l=0.15
X1219 avdd.t235 por_ana_0.rstring_mux_0.ena_b por_ana_0.rstring_mux_0.vtop.t8 avdd.t234 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X1220 dvss.t1832 dvdd.t1857 dvss.t1831 dvss.t1784 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X1221 a_19094_1626# a_41694_1248# dvss.t1443 sky130_fd_pr__res_xhigh_po_1p41 l=111
X1222 dvss.t1830 dvdd.t1858 dvss.t1829 dvss.t1828 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1223 avdd.t111 avdd.t109 avdd.t110 avdd.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=8
X1224 a_37658_33453# a_37614_33695# a_37492_33453# dvss.t356 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X1225 a_33996_36477# por_dig_0.net24 dvdd.t347 dvdd.t346 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X1226 a_21622_21903# a_21254_22885# dvss.t1071 dvss.t1070 sky130_fd_pr__nfet_01v8 ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X1227 dvss.t2045 por_dig_0.net21 a_39732_31829# dvss.t2044 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X1228 por_ana_0.ibias_gen_0.vn1.t0 avdd.t107 por_ana_0.ibias_gen_0.vp1.t0 avdd.t108 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X1229 por_ana_0.comparator_0.vinn.t3 avdd.t105 por_ana_0.comparator_0.vinn.t3 avdd.t106 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=0.6
X1230 a_35704_35124# por_dig_0._046_ a_35632_35124# dvdd.t1478 sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X1231 avdd.t484 por_ana_0.comparator_0.n1.t9 por_ana_0.dcomp3v3uv avdd.t483 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X1232 a_23466_24707# a_23366_24619# dvss.t1522 dvss.t1521 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X1233 a_34378_30189# a_34212_30189# dvss.t1282 dvss.t1281 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1234 dvdd.t1176 por_dig_0.net8 a_31412_31251# dvdd.t1175 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X1235 avdd.t652 a_28383_21859# a_27690_22973# avdd.t651 sky130_fd_pr__pfet_g5v0d10v5 ad=0.2142 pd=1.99 as=0.2142 ps=1.99 w=0.42 l=1
X1236 dvdd.t1665 dvss.t2285 dvdd.t1664 dvdd.t1556 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X1237 a_32809_32365# a_31728_32365# a_32462_32607# dvdd.t585 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X1238 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[2] a_33121_22637# avdd.t463 avdd.t254 sky130_fd_pr__pfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.24375 ps=1.825 w=1.5 l=0.5
X1239 a_33474_35059# a_33256_35463# dvss.t1224 dvss.t1223 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X1240 por_dig_0._051_ por_dig_0.cnt_por\[1\] dvdd.t1162 dvdd.t1161 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.3 ps=2.6 w=1 l=0.15
X1241 por_dig_0._035_ por_dig_0.cnt_por\[6\] dvdd.t392 dvdd.t391 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1242 por_dig_0.net13 a_33155_28640# dvss.t1449 dvss.t1448 sky130_fd_pr__nfet_01v8 ad=0.221 pd=1.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X1243 dvss.t1974 a_25578_22973# a_26785_22637# dvss.t1973 sky130_fd_pr__nfet_g5v0d10v5 ad=0.121875 pd=1.075 as=0.19875 ps=2.03 w=0.75 l=0.5
X1244 a_33380_35879# por_dig_0._047_ a_33162_35603# dvdd.t726 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.26 ps=2.52 w=1 l=0.15
X1245 dvss.t989 por_dig_0.net34 a_38904_31277# dvss.t988 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1246 a_31802_32909# a_31566_32909# dvss.t1451 dvss.t1450 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.5
X1247 dvss.t1047 a_33805_32339# por_dig_0._024_ dvss.t1046 sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.17225 ps=1.83 w=0.65 l=0.15
X1248 por_ana_0.comparator_1.vt.t28 vin.t57 por_ana_0.comparator_1.vpp.t38 por_ana_0.comparator_1.vt.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1249 a_37474_31099# a_37430_30707# a_37308_31111# dvss.t1965 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X1250 dvss.t1411 a_23734_21903# a_24159_21859# dvss.t1410 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X1251 por_dig_0.cnt_por\[7\] a_32984_32339# dvdd.t1040 dvdd.t1039 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X1252 a_36414_32909# por_dig_0.net23.t12 dvdd.t763 dvdd.t762 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.1475 ps=1.295 w=1 l=0.15
X1253 dvdd.t1668 dvss.t2286 dvdd.t1667 dvdd.t1666 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1254 por_ana_0.rstring_mux_0.otrip_decoded_b_avdd[0] por_ana_0.rstring_mux_0.otrip_decoded_avdd[0] avss.t308 avss.t307 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X1255 a_34898_29351# a_34828_29253# por_dig_0.net15 dvdd.t668 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.32 ps=2.64 w=1 l=0.15
X1256 por_dig_0.otrip_decoded[2].t0 a_33752_28013# dvss.t966 dvss.t523 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X1257 dvss.t2213 a_32535_28013# a_32641_28013# dvss.t677 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X1258 a_36831_23593# a_36406_23637# dvss.t974 dvss.t973 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X1259 a_35686_29351# por_dig_0.net7.t11 dvdd.t739 dvdd.t668 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1260 dvss.t2024 por_dig_0.otrip_decoded[2].t5 a_23366_22885# dvss.t2023 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X1261 dvdd.t1519 a_31413_29075# por_dig_0.force_pdnb dvdd.t668 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X1262 por_dig_0.clknet_1_0__leaf_osc_ck.t8 a_34098_30707# dvss.t196 dvss.t195 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1263 por_ana_0.sky130_fd_sc_hvl__inv_4_0.A por_ana_0.sky130_fd_sc_hvl__inv_1_0.A avss.t231 avss.t230 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X1264 a_23456_13935# a_23834_6535# avss.t232 sky130_fd_pr__res_xhigh_po_1p41 l=35
X1265 a_32812_30733# a_32188_30739# a_32704_31111# dvdd.t818 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X1266 dvss.t457 por_dig_0.cnt_por\[6\] por_dig_0._022_ dvss.t456 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X1267 dvss.t758 a_39888_24823# a_39888_23693# dvss.t757 sky130_fd_pr__nfet_g5v0d10v5 ad=0.178875 pd=1.26 as=0.1197 ps=1.41 w=0.42 l=0.5
X1268 dvdd.t5 a_32701_28531# por_dig_0.otrip_decoded[1] dvdd.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X1269 avdd.t104 avdd.t103 avdd.t104 avdd.t33 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=8
X1270 dvdd.t812 por_dig_0.cnt_st\[3\] por_dig_0._042_ dvdd.t256 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1271 por_ana_0.rstring_mux_0.vtrip_decoded_b_avdd[7] por_ana_0.rstring_mux_0.vtrip_decoded_avdd[7].t4 avss.t395 avss.t394 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X1272 dvss.t321 a_32610_35603# por_dig_0._007_ dvss.t320 sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X1273 a_33821_35463# a_32740_35091# a_33474_35059# dvdd.t1034 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X1274 por_dig_0._036_.t2 por_dig_0._035_ dvss.t2068 dvss.t2067 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1275 por_ana_0.comparator_0.vpp.t35 por_ana_0.comparator_0.vnn.t51 avdd.t366 avdd.t191 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1276 por_ana_0.rc_osc_0.in dvss.t290 sky130_fd_pr__cap_mim_m3_2 l=30 w=30
X1277 por_ana_0.comparator_1.vpp.t23 por_ana_0.comparator_1.vnn.t53 avdd.t639 avdd.t395 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1278 a_18154_35244# a_17776_27844# avss.t233 sky130_fd_pr__res_xhigh_po_1p41 l=35
X1279 dvss.t765 a_27690_24707# a_28897_24371# dvss.t764 sky130_fd_pr__nfet_g5v0d10v5 ad=0.121875 pd=1.075 as=0.19875 ps=2.03 w=0.75 l=0.5
X1280 porb_h.t6 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.t20 avdd.t341 avdd.t340 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X1281 a_36581_35629# a_35500_35629# a_36234_35871# dvdd.t439 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X1282 por_dig_0.clknet_1_0__leaf_osc_ck.t26 a_34098_30707# dvdd.t169 dvdd.t168 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1283 por_dig_0._025_ por_dig_0.cnt_por\[7\] a_33450_33453# dvss.t1093 sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.10725 ps=0.98 w=0.65 l=0.15
X1284 a_24159_21859# a_23734_21903# dvss.t1409 dvss.t1408 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X1285 a_33996_36477# a_33821_36551# a_34175_36539# dvss.t444 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X1286 dvdd.t1670 dvss.t2287 a_31814_22885# dvdd.t1669 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X1287 a_36138_24707# a_36038_24619# dvss.t680 dvss.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X1288 dvss.t804 por_dig_0.por_unbuf.t11 por_ana_0.sky130_fd_sc_hd__inv_4_4.Y dvss.t803 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1289 por_dig_0._000_ por_dig_0.net31 dvdd.t856 dvdd.t855 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1290 a_31413_32339# por_dig_0.net19 dvdd.t1012 dvdd.t1011 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X1291 dvdd.t1310 a_32462_32607# a_32352_32731# dvdd.t1309 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X1292 por_ana_0.schmitt_trigger_0.in.t8 dvss.t656 sky130_fd_pr__cap_mim_m3_2 l=30 w=30
X1293 dvss.t103 a_33804_31251# por_dig_0._027_ dvss.t102 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1294 dvss.t349 por_ana_0.sky130_fd_sc_hd__inv_4_1.Y porb.t12 dvss.t348 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1295 vin.t13 por_ana_0.rstring_mux_0.otrip_decoded_avdd[1] por_ana_0.rstring_mux_0.vtrip1.t3 avss.t31 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X1296 dvdd.t1672 dvss.t2288 a_31814_24619# dvdd.t1671 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X1297 a_35030_28557# por_dig_0.net5.t6 dvdd.t1441 dvdd.t1440 sky130_fd_pr__pfet_01v8_hvt ad=0.1087 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X1298 a_15896_13935# a_16274_6535# avss.t234 sky130_fd_pr__res_xhigh_po_1p41 l=35
X1299 a_35219_34541# por_dig_0.net23.t13 dvss.t876 dvss.t875 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10025 ps=0.985 w=0.65 l=0.15
X1300 por_dig_0.cnt_por\[2\] a_33996_36477# dvdd.t1266 dvdd.t1265 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X1301 a_35217_28917# a_35030_28557# a_35130_28673# dvss.t104 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.107825 ps=1.36 w=0.42 l=0.15
X1302 por_dig_0.clknet_1_0__leaf_osc_ck.t7 a_34098_30707# dvss.t194 dvss.t193 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X1303 dvdd.t1675 dvss.t2289 dvdd.t1674 dvdd.t1673 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1304 force_dis_rc_osc.t1 dvss.t1622 dvss.t1624 dvss.t1623 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X1305 por_ana_0.comparator_0.vpp.t36 por_ana_0.comparator_0.vnn.t52 avdd.t367 avdd.t191 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1306 dvss.t1421 por_dig_0.net8 a_31864_30823# dvss.t1420 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X1307 avdd.t102 avdd.t100 avdd.t101 avdd.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=8
X1308 a_35746_36539# por_dig_0.cnt_por\[0\].t13 a_35674_36539# dvss.t640 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X1309 dvss.t1827 dvdd.t1859 dvss.t1826 dvss.t1825 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1310 dvdd.t123 a_34387_32909# por_dig_0.clknet_0_osc_ck.t26 dvdd.t122 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1311 avdd.t368 por_ana_0.comparator_0.vnn.t53 por_ana_0.comparator_0.vpp.t37 avdd.t195 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1312 dvss.t1000 a_25846_21903# a_26271_21859# dvss.t999 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X1313 dvss.t398 a_39887_23089# a_40246_23089# dvss.t396 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X1314 a_34102_29645# por_dig_0.net30 dvdd.t308 dvdd.t70 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1315 dvdd.t1490 por_dig_0._019_ a_34580_34110# dvdd.t1489 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X1316 dvss.t756 a_39888_24823# a_40247_24823# dvss.t754 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X1317 dvss.t42 a_38150_24619# a_38250_24707# dvss.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X1318 avss.t89 avss.t88 avss.t89 avss.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=8
X1319 por_dig_0.clknet_1_1__leaf_osc_ck.t10 a_35583_34541# dvss.t586 dvss.t585 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1320 a_37492_33453# a_37046_33453# a_37396_33453# dvss.t18 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X1321 dvss.t151 a_34387_32909# por_dig_0.clknet_0_osc_ck.t8 dvss.t150 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1322 avdd.t343 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.t21 porb_h.t5 avdd.t342 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X1323 a_34830_35629# por_dig_0.cnt_por\[3\] a_34580_35629# dvss.t452 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1324 dvdd.t1677 dvss.t2290 dvdd.t1676 dvdd.t1537 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1325 a_32794_33971# por_dig_0._047_ dvss.t843 dvss.t842 sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.25675 ps=1.44 w=0.65 l=0.15
X1326 a_33996_35389# a_33821_35463# a_34175_35451# dvss.t738 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X1327 a_36940_35463# a_36494_35091# a_36844_35463# dvss.t996 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X1328 a_31413_32339# por_dig_0.net19 dvss.t1202 dvss.t1201 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X1329 a_38943_23593# a_38518_23637# dvss.t2215 dvss.t2214 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X1330 dvss.t2114 por_dig_0.net5.t7 a_32358_28013# dvss.t677 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X1331 dvdd.t1022 a_33474_35059# a_33364_35085# dvdd.t1021 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X1332 a_32607_21859# a_32182_21903# dvss.t1120 dvss.t1119 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X1333 a_31914_22973# a_31814_22885# dvss.t2162 dvss.t2161 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X1334 por_ana_0.rstring_mux_0.vtrip4.t1 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[4].t4 por_ana_0.comparator_0.vinn.t43 avss.t328 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X1335 vin.t11 por_ana_0.rstring_mux_0.otrip_decoded_b_avdd[1] por_ana_0.rstring_mux_0.vtrip1.t1 avdd.t215 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X1336 por_ana_0.comparator_1.vnn.t44 vbg_1v2.t21 por_ana_0.comparator_1.vt.t48 por_ana_0.comparator_1.vt.t36 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1337 dvdd.t1324 a_36234_35871# a_36124_35995# dvdd.t1323 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X1338 por_dig_0.net28 a_31908_32909# dvss.t1434 dvss.t1433 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X1339 por_ana_0.ibias_gen_0.vstart.t3 vbg_1v2.t22 por_ana_0.ibias_gen_0.vn0.t12 avss.t150 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X1340 por_ana_0.comparator_1.vnn.t23 por_ana_0.comparator_1.vpp.t55 avdd.t411 avdd.t403 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1341 dvss.t856 por_dig_0.net7.t12 a_34934_28013# dvss.t677 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X1342 dcomp.t20 por_ana_0.sky130_fd_sc_hd__inv_4_3.Y dvdd.t45 dvdd.t44 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1343 avss.t19 por_ana_0.comparator_1.n1.t10 por_ana_0.dcomp3v3 avss.t18 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X1344 a_33821_35463# a_32906_35091# a_33474_35059# dvss.t1207 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X1345 a_35111_28013# a_34934_28013# dvdd.t893 dvdd.t892 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X1346 dvss.t1031 a_39888_23693# a_40247_23627# dvss.t1029 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.105 ps=1.03 w=0.75 l=0.5
X1347 a_35570_33453# a_35092_33427# dvss.t393 dvss.t392 sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.12495 ps=1.015 w=0.42 l=0.15
X1348 por_ana_0.sky130_fd_sc_hd__inv_4_1.A por_dig_0.por_unbuf.t12 dvss.t806 dvss.t805 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1349 por_ana_0.dcomp3v3uv por_ana_0.comparator_0.n1.t10 avss.t273 avss.t272 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X1350 a_32019_31643# a_31893_31545# a_31615_31529# dvss.t20 sky130_fd_pr__special_nfet_01v8 ad=0.0999 pd=0.985 as=0.0711 ps=0.755 w=0.36 l=0.15
X1351 por_ana_0.comparator_0.vpp.t5 por_ana_0.comparator_0.vpp.t4 avdd.t194 avdd.t191 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1352 dvdd.t1679 dvss.t2291 a_33926_22885# dvdd.t1678 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X1353 a_40246_23089# a_39887_23089# dvss.t397 dvss.t396 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.178875 ps=1.26 w=0.75 l=0.5
X1354 dvdd.t676 por_dig_0.net6 a_34982_29351# dvdd.t668 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.135 ps=1.27 w=1 l=0.15
X1355 a_40247_24823# a_39888_24823# dvss.t755 dvss.t754 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.178875 ps=1.26 w=0.75 l=0.5
X1356 a_37320_30733# por_dig_0.net25 dvdd.t839 dvdd.t838 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X1357 por_dig_0.net33 a_39268_33453# dvdd.t135 dvdd.t134 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X1358 dvdd.t643 a_33720_33213# a_33707_32909# dvdd.t642 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X1359 dvdd.t1681 dvss.t2292 a_33926_24619# dvdd.t1680 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X1360 dvss.t2088 a_36512_28013# por_dig_0.otrip_decoded[5].t1 dvss.t523 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X1361 porb_h.t4 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.t22 avdd.t345 avdd.t344 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X1362 dvdd.t507 por_dig_0.cnt_st\[1\] a_38352_32365# dvdd.t506 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1363 dvss.t957 por_dig_0.net25 a_37474_31099# dvss.t956 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X1364 avss.t185 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.t23 porb_h.t28 avss.t184 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X1365 a_33518_36539# a_33474_36147# a_33352_36551# dvss.t1034 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X1366 a_38957_32883# por_dig_0.net4 dvss.t94 dvss.t93 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.10075 ps=0.96 w=0.65 l=0.15
X1367 dvss.t1824 dvdd.t1860 dvss.t1823 dvss.t1682 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1368 a_36380_33971# por_dig_0.net23.t14 dvss.t878 dvss.t877 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.06825 ps=0.745 w=0.42 l=0.15
X1369 a_34738_32141# por_dig_0.cnt_por\[4\] a_34654_32141# dvss.t1549 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X1370 a_35740_31277# a_35224_31277# a_35645_31277# dvss.t1288 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X1371 por_ana_0.comparator_1.vnn.t22 por_ana_0.comparator_1.vpp.t56 avdd.t412 avdd.t403 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1372 avss.t346 por_ana_0.comparator_1.vm.t7 por_ana_0.comparator_1.n0.t3 avss.t292 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1373 por_ana_0.comparator_1.vt.t9 avss.t424 por_ana_0.comparator_1.vnn.t33 por_ana_0.comparator_1.vt.t3 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=8
X1374 a_34265_27987# por_dig_0.net15 dvdd.t889 dvdd.t888 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X1375 pwup_filt.t9 por_ana_0.sky130_fd_sc_hd__inv_4_0.Y dvss.t246 dvss.t245 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1376 dvdd.t1684 dvss.t2293 dvdd.t1683 dvdd.t1682 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X1377 por_ana_0.rstring_mux_0.vtrip4.t3 por_ana_0.rstring_mux_0.vtrip_decoded_b_avdd[4] por_ana_0.comparator_0.vinn.t32 avdd.t470 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X1378 a_37046_33453# a_36880_33453# dvdd.t653 dvdd.t652 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1379 dvss.t2198 a_27958_21903# a_28383_21859# dvss.t2197 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X1380 avdd.t277 por_ana_0.sky130_fd_sc_hvl__inv_4_0.A por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.t1 avdd.t276 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X1381 por_dig_0.net23.t1 a_36564_32339# dvss.t691 dvss.t690 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1382 por_dig_0._003_ a_39077_31527# dvss.t1440 dvss.t1439 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1383 a_37504_33819# a_36880_33453# a_37396_33453# dvdd.t651 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X1384 por_ana_0.comparator_0.vpp.t3 por_ana_0.comparator_0.vpp.t2 avdd.t193 avdd.t191 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1385 por_ana_0.rstring_mux_0.vtrip6.t6 por_ana_0.rstring_mux_0.otrip_decoded_avdd[6] vin.t42 avss.t373 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X1386 a_40247_23627# a_39888_23693# dvss.t1030 dvss.t1029 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.178875 ps=1.26 w=0.75 l=0.5
X1387 a_37596_30555# a_36972_30189# a_37488_30189# dvdd.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X1388 a_31412_31251# a_31615_31529# dvdd.t1086 dvdd.t1085 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1134 ps=1.38 w=0.42 l=0.15
X1389 dvdd.t879 a_37584_35389# por_dig_0.cnt_por\[1\] dvdd.t878 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1390 a_40246_23089# a_40246_21893# dvdd.t900 dvdd.t899 sky130_fd_pr__pfet_01v8_hvt ad=0.2968 pd=2.77 as=0.1568 ps=1.4 w=1.12 l=0.15
X1391 dvss.t216 por_dig_0.net29 a_34496_29645# dvss.t215 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1392 dvss.t1200 por_dig_0.net19 a_31592_30965# dvss.t1199 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1393 dvss.t1822 dvdd.t1861 dvss.t1821 dvss.t1820 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X1394 dvdd.t1686 dvss.t2294 dvdd.t1685 dvdd.t1540 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1395 dvss.t2116 por_dig_0.net5.t8 por_dig_0.net13 dvss.t2115 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1396 dvss.t2188 a_35000_31795# por_dig_0._028_ dvss.t2187 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1397 a_34719_21859# a_34294_21903# dvss.t1495 dvss.t1494 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X1398 a_16642_35244# a_17020_27844# avss.t235 sky130_fd_pr__res_xhigh_po_1p41 l=35
X1399 por.t29 por_ana_0.sky130_fd_sc_hd__inv_4_4.Y dvdd.t974 dvdd.t973 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1400 por_ana_0.comparator_1.ena_b por_ana_0.rstring_mux_0.ena.t6 avdd.t608 avdd.t607 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X1401 dvss.t2007 por_dig_0.cnt_rsb_stg1 a_31566_32909# dvss.t2006 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1402 a_35582_34317# por_dig_0._048_ por_dig_0._009_ dvss.t1111 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1403 a_34026_22973# a_33926_22885# dvss.t612 dvss.t611 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X1404 por_ana_0.dcomp3v3 por_ana_0.comparator_1.n1.t11 avdd.t533 avdd.t532 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X1405 a_31876_32199# a_31526_31827# a_31781_32187# dvdd.t946 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X1406 avdd.t399 por_ana_0.comparator_1.vpp.t12 por_ana_0.comparator_1.vpp.t13 avdd.t392 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1407 a_33518_35451# a_33474_35059# a_33352_35463# dvss.t1211 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X1408 por_ana_0.sky130_fd_sc_hvl__inv_1_0.A a_26802_33372# avdd.t446 avdd.t445 sky130_fd_pr__pfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.24375 ps=1.825 w=1.5 l=0.5
X1409 dvdd.t972 por_ana_0.sky130_fd_sc_hd__inv_4_4.Y por.t28 dvdd.t971 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1410 vin.t18 avss.t86 vin.t18 avss.t87 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=0.6
X1411 por_ana_0.comparator_1.vnn avss.t425 por_ana_0.comparator_1.vt.t8 por_ana_0.comparator_1.vt.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=8
X1412 a_34265_27987# por_dig_0.net15 dvss.t1022 dvss.t677 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X1413 por_ana_0.comparator_1.vn.t1 por_ana_0.comparator_1.ena_b avss.t255 avss.t254 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X1414 a_35295_33705# a_35573_33721# a_35529_33819# dvdd.t1317 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0567 ps=0.69 w=0.42 l=0.15
X1415 dvss.t1333 por_dig_0.cnt_st\[0\] a_39720_32365# dvss.t1332 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.095875 ps=0.945 w=0.65 l=0.15
X1416 a_37798_33971# a_37580_34375# dvdd.t1078 dvdd.t1077 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X1417 a_35289_28917# por_dig_0.net6 a_35217_28917# dvss.t798 sky130_fd_pr__nfet_01v8 ad=0.05355 pd=0.675 as=0.0441 ps=0.63 w=0.42 l=0.15
X1418 por_ana_0.rc_osc_0.m por_ana_0.rc_osc_0.in dvdd.t239 dvdd.t238 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.1475 ps=1.295 w=1 l=0.5
X1419 dvdd.t1424 por_dig_0.osc_ena.t5 por_ana_0.rc_osc_0.in dvdd.t1423 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X1420 porb.t11 por_ana_0.sky130_fd_sc_hd__inv_4_1.Y dvss.t347 dvss.t346 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1421 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.t0 por_ana_0.sky130_fd_sc_hvl__inv_4_0.A avdd.t275 avdd.t274 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.4275 ps=3.57 w=1.5 l=0.5
X1422 dvss.t1819 dvdd.t1862 dvss.t1818 dvss.t1743 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X1423 a_38500_31251# por_dig_0.cnt_st\[4\] dvdd.t1244 dvdd.t1243 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1424 dvss.t2066 por_dig_0._035_ a_36567_32141# dvss.t2065 sky130_fd_pr__nfet_01v8 ad=0.1365 pd=1.07 as=0.117 ps=1.01 w=0.65 l=0.15
X1425 a_37046_32915# a_36880_32915# dvss.t521 dvss.t520 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1426 por_ana_0.comparator_1.vnn.t21 por_ana_0.comparator_1.vpp.t57 avdd.t413 avdd.t403 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1427 dvss.t558 a_36756_35603# a_36690_35629# dvss.t557 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X1428 por_dig_0.otrip_decoded[7].t2 a_37156_28013# dvdd.t655 dvdd.t654 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X1429 por_ana_0.rstring_mux_0.vtrip6.t8 por_ana_0.rstring_mux_0.otrip_decoded_b_avdd[6] vin.t44 avdd.t594 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X1430 dvdd.t1689 dvss.t2295 dvdd.t1688 dvdd.t1687 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1431 dvss.t1493 a_34294_21903# a_34719_21859# dvss.t1492 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X1432 dvss.t922 por_dig_0._038_ a_31717_30189# dvss.t921 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.08775 ps=0.92 w=0.65 l=0.15
X1433 por_dig_0.clknet_1_0__leaf_osc_ck.t25 a_34098_30707# dvdd.t167 dvdd.t166 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X1434 dvss.t345 por_ana_0.sky130_fd_sc_hd__inv_4_1.Y porb.t10 dvss.t344 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1435 a_37706_30431# a_37488_30189# dvss.t270 dvss.t269 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X1436 por_ana_0.ibias_gen_0.vr.t3 por_ana_0.ibias_gen_0.vn0.t19 por_ana_0.ibias_gen_0.vp0.t7 avss.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X1437 dvss.t1991 a_33896_35603# por_dig_0._053_ dvss.t1990 sky130_fd_pr__nfet_01v8 ad=0.160875 pd=1.145 as=0.169 ps=1.82 w=0.65 l=0.15
X1438 dvss.t745 a_33720_33213# a_33654_33287# dvss.t744 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X1439 a_32441_32199# a_31360_31827# a_32094_31795# dvdd.t23 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X1440 a_35402_30189# a_34212_30189# a_35293_30189# dvss.t1280 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1441 dvdd.t417 por_dig_0.clknet_1_0__leaf_osc_ck.t39 a_32188_30739# dvdd.t416 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1442 por_dig_0._030_ a_38352_32365# dvss.t731 dvss.t730 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X1443 dvss.t2110 por_dig_0.otrip_decoded[5].t5 a_25478_24619# dvss.t2109 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X1444 por_ana_0.rstring_mux_0.otrip_decoded_avdd[1] a_22561_24371# avdd.t493 avdd.t298 sky130_fd_pr__pfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.24375 ps=1.825 w=1.5 l=0.5
X1445 avss.t47 avss.t44 avss.t46 avss.t45 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=8
X1446 dvss.t174 por_dig_0._031_ por_dig_0._032_ dvss.t173 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1447 a_37706_30431# a_37488_30189# dvdd.t227 dvdd.t226 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X1448 dvss.t1017 a_37584_35389# a_37518_35463# dvss.t1016 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X1449 vin.t6 avdd.t98 vin.t6 avdd.t99 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=0.6
X1450 por_ana_0.sky130_fd_sc_hd__inv_4_1.Y por_ana_0.sky130_fd_sc_hd__inv_4_1.A dvdd.t191 dvdd.t190 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1451 a_32352_32731# por_dig_0.net24 dvdd.t345 dvdd.t344 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X1452 dvdd.t505 por_dig_0.cnt_st\[1\] a_38956_32339# dvdd.t504 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0735 ps=0.77 w=0.42 l=0.15
X1453 a_30495_23593# a_30070_23637# dvss.t1292 dvss.t1291 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X1454 por_ana_0.comparator_1.vnn.t20 por_ana_0.comparator_1.vpp.t58 avdd.t414 avdd.t403 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1455 a_36831_21859# a_36406_21903# dvss.t1316 dvss.t1315 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X1456 dvdd.t1692 dvss.t2296 dvdd.t1691 dvdd.t1690 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X1457 a_36078_33453# a_35699_33819# a_36006_33453# dvss.t1394 sky130_fd_pr__nfet_01v8 ad=0.1401 pd=1.1 as=0.0441 ps=0.63 w=0.42 l=0.15
X1458 dvdd.t121 a_34387_32909# por_dig_0.clknet_0_osc_ck.t25 dvdd.t120 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1459 por_ana_0.rstring_mux_0.vtrip_decoded_b_avdd[2] por_ana_0.rstring_mux_0.vtrip_decoded_avdd[2] avss.t264 avss.t263 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X1460 a_38146_31429# a_38242_31251# dvss.t1318 dvss.t1317 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.5
X1461 avdd.t97 avdd.t96 avdd.t97 avdd.t33 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=8
X1462 por_dig_0.clknet_1_1__leaf_osc_ck.t9 a_35583_34541# dvss.t584 dvss.t583 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1463 dvdd.t1098 a_32441_32199# a_32616_32125# dvdd.t1097 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X1464 dvdd.t248 por_dig_0._032_ a_37789_31821# dvdd.t247 sky130_fd_pr__pfet_01v8_hvt ad=0.3275 pd=1.655 as=0.195 ps=1.39 w=1 l=0.15
X1465 por_ana_0.comparator_0.vinn.t23 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[0] por_ana_0.rstring_mux_0.vtrip0.t2 avss.t222 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X1466 avdd.t476 a_30495_23593# a_29802_24707# avdd.t475 sky130_fd_pr__pfet_g5v0d10v5 ad=0.2142 pd=1.99 as=0.2142 ps=1.99 w=0.42 l=1
X1467 a_32352_32731# a_31728_32365# a_32244_32365# dvdd.t584 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X1468 osc_ck.t7 por_dig_0.osc_ena.t6 por_ana_0.rc_osc_0.vr dvss.t2098 sky130_fd_pr__nfet_01v8 ad=0.15 pd=1.3 as=0.1475 ps=1.295 w=1 l=0.18
X1469 dvss.t1621 dvss.t1619 otrip[2].t0 dvss.t1620 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X1470 dvss.t1817 dvdd.t1863 dvss.t1816 dvss.t1815 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X1471 a_36862_30739# a_36696_30739# dvdd.t1064 dvdd.t1063 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1472 a_34580_35629# por_dig_0.cnt_por\[2\] dvss.t1578 dvss.t1577 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1473 a_37492_33287# a_37046_32915# a_37396_33287# dvss.t18 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X1474 por_ana_0.sky130_fd_sc_hd__inv_4_3.Y por_ana_0.vl dvdd.t1000 dvdd.t999 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1475 a_36381_36691# por_dig_0.net20.t5 dvss.t2105 dvss.t1110 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X1476 dcomp.t19 por_ana_0.sky130_fd_sc_hd__inv_4_3.Y dvdd.t43 dvdd.t42 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1477 a_32528_13935# a_32150_6535# avss.t284 sky130_fd_pr__res_xhigh_po_1p41 l=35
X1478 a_25578_22973# a_25478_22885# dvss.t1564 dvss.t1563 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X1479 por_dig_0.net21 a_38936_32159# dvdd.t1380 dvdd.t1379 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X1480 a_37504_32909# a_36880_32915# a_37396_33287# dvdd.t432 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X1481 dvss.t244 por_ana_0.sky130_fd_sc_hd__inv_4_0.Y pwup_filt.t8 dvss.t243 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1482 a_31914_24707# a_31814_24619# dvss.t2051 dvss.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X1483 a_37138_30189# a_36972_30189# dvss.t28 dvss.t27 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1484 a_33352_36551# a_32906_36179# a_33256_36551# dvss.t721 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X1485 a_33623_31099# por_dig_0.net24 dvss.t433 dvss.t432 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X1486 a_35433_32141# por_dig_0.net4 dvss.t92 dvss.t91 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X1487 avdd.t398 por_ana_0.comparator_1.vpp.t10 por_ana_0.comparator_1.vpp.t11 avdd.t392 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1488 por_dig_0.clknet_0_osc_ck.t24 a_34387_32909# dvdd.t119 dvdd.t118 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1489 a_2543_22912# a_2921_15512# avss.t27 sky130_fd_pr__res_xhigh_po_1p41 l=35
X1490 a_33284_13935# a_33662_6535# avss.t285 sky130_fd_pr__res_xhigh_po_1p41 l=35
X1491 a_33474_36147# a_33256_36551# dvdd.t1194 dvdd.t1193 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X1492 dvdd.t41 por_ana_0.sky130_fd_sc_hd__inv_4_3.Y dcomp.t18 dvdd.t40 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1493 dvss.t582 a_35583_34541# por_dig_0.clknet_1_1__leaf_osc_ck.t8 dvss.t581 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1494 dvdd.t1512 a_32094_31795# a_31984_31821# dvdd.t1511 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X1495 dvss.t1814 dvdd.t1864 dvss.t1813 dvss.t1812 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1496 pwup_filt.t7 por_ana_0.sky130_fd_sc_hd__inv_4_0.Y dvss.t242 dvss.t241 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1497 dvss.t1618 dvss.t1616 por_ana_0.rc_osc_0.n.t4 dvss.t1617 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X1498 avdd.t95 avdd.t94 avdd.t95 avdd.t33 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=8
X1499 por_ana_0.ibias_gen_0.vstart.t2 vbg_1v2.t23 por_ana_0.ibias_gen_0.vn0.t13 avss.t151 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X1500 por_ana_0.rstring_mux_0.vtop.t7 por_ana_0.rstring_mux_0.ena_b avdd.t233 avdd.t232 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X1501 dvss.t1314 a_36406_21903# a_36831_21859# dvss.t1313 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X1502 por_dig_0.net24 a_35100_32339# dvss.t1244 dvss.t1243 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1218 ps=1.42 w=0.42 l=0.15
X1503 a_29504_13935# a_29126_6535# avss.t286 sky130_fd_pr__res_xhigh_po_1p41 l=35
X1504 dvss.t808 por_dig_0.por_unbuf.t13 por_ana_0.sky130_fd_sc_hd__inv_4_1.A dvss.t807 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1505 dvdd.t1694 dvss.t2297 dvdd.t1693 dvdd.t1522 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1506 avdd.t93 avdd.t91 avdd.t92 avdd.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=8
X1507 dvdd.t970 por_ana_0.sky130_fd_sc_hd__inv_4_4.Y por.t27 dvdd.t969 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1508 a_39349_32909# por_dig_0.net21 a_39094_32909# dvdd.t1384 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.14 ps=1.28 w=1 l=0.15
X1509 dvss.t382 a_33444_31037# a_33378_31111# dvss.t381 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X1510 por_ana_0.comparator_1.vnn.t46 por_ana_0.rstring_mux_0.ena.t7 avdd.t610 avdd.t609 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X1511 a_32651_33819# a_31893_33721# a_32088_33690# dvdd.t408 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.07245 ps=0.765 w=0.42 l=0.15
X1512 por_ana_0.rstring_mux_0.otrip_decoded_avdd[5] a_26785_24371# avdd.t496 avdd.t302 sky130_fd_pr__pfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.24375 ps=1.825 w=1.5 l=0.5
X1513 a_34109_33453# por_dig_0._020_ a_33806_33427# dvss.t2146 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.089375 ps=0.925 w=0.65 l=0.15
X1514 por_ana_0.comparator_0.vinn.t25 por_ana_0.rstring_mux_0.vtrip_decoded_b_avdd[0] por_ana_0.rstring_mux_0.vtrip0.t4 avdd.t426 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X1515 avdd.t231 por_ana_0.rstring_mux_0.ena_b por_ana_0.rstring_mux_0.vtop.t6 avdd.t230 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X1516 a_33364_35085# a_32740_35091# a_33256_35463# dvdd.t1033 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X1517 a_33707_32909# a_32630_32915# a_33545_33287# dvdd.t859 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X1518 por_ana_0.ibias_gen_0.vp1.t14 por_ana_0.ibias_gen_0.isrc_sel_b.t6 por_ana_0.ibias_gen_0.vp.t2 avdd.t576 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X1519 por_dig_0.otrip_decoded[5].t0 a_36512_28013# dvss.t2087 dvss.t523 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X1520 dvdd.t137 a_34746_31277# a_34852_31277# dvdd.t136 sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.5
X1521 dvss.t2097 por_dig_0.otrip_decoded[7].t5 a_27590_24619# dvss.t2096 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X1522 a_34728_30189# a_34378_30189# a_34633_30189# dvdd.t1121 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X1523 por_ana_0.comparator_1.vnn.t43 vbg_1v2.t24 por_ana_0.comparator_1.vt.t47 por_ana_0.comparator_1.vt.t36 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1524 dvdd.t724 a_31413_32339# por_timed_out.t3 dvdd.t723 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X1525 por_dig_0.cnt_por\[3\] a_33996_35389# dvss.t1266 dvss.t1265 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X1526 dvss.t2100 por_dig_0.osc_ena.t7 por_ana_0.rc_osc_0.ena_b dvss.t2099 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.6
X1527 por_ana_0.ibias_gen_0.ibias0.t0 por_ana_0.ibias_gen_0.vp.t8 avdd.t381 avdd.t380 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X1528 dvss.t865 por_dig_0._034_.t12 por_dig_0._036_.t0 dvss.t864 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1529 por_ana_0.comparator_0.vnn.t26 por_ana_0.comparator_0.vinn.t56 por_ana_0.comparator_0.vt.t9 por_ana_0.comparator_0.vt.t3 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1530 a_32607_23593# a_32182_23637# dvss.t9 dvss.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X1531 por_ana_0.comparator_1.vnn.t42 vbg_1v2.t25 por_ana_0.comparator_1.vt.t46 por_ana_0.comparator_1.vt.t36 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1532 a_38943_21859# a_38518_21903# dvss.t268 dvss.t267 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X1533 dvss.t240 por_ana_0.sky130_fd_sc_hd__inv_4_0.Y pwup_filt.t6 dvss.t239 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1534 por_ana_0.comparator_0.vinn.t39 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[1] por_ana_0.rstring_mux_0.vtrip1.t9 avss.t316 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X1535 porb_h.t3 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.t24 avdd.t347 avdd.t346 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X1536 avdd.t90 avdd.t88 avdd.t89 avdd.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=8
X1537 por_ana_0.comparator_0.vt.t45 vbg_1v2.t26 por_ana_0.comparator_0.vpp.t24 por_ana_0.comparator_0.vt.t36 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1538 avdd.t271 a_32607_23593# a_31914_24707# avdd.t270 sky130_fd_pr__pfet_g5v0d10v5 ad=0.2142 pd=1.99 as=0.2142 ps=1.99 w=0.42 l=1
X1539 a_36567_31821# por_dig_0._034_.t13 dvdd.t751 dvdd.t750 sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.3125 ps=1.625 w=1 l=0.15
X1540 a_22047_23593# a_21622_23637# dvss.t1232 dvss.t1231 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X1541 a_34444_32517# por_dig_0.net32 dvdd.t320 dvdd.t319 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.365 ps=1.73 w=1 l=0.15
X1542 a_34496_29645# por_dig_0._028_ dvss.t371 dvss.t370 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1543 a_35293_30189# a_34378_30189# a_34946_30431# dvss.t1350 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X1544 dvdd.t1208 a_35612_33595# a_35573_33721# dvdd.t1207 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1545 a_31592_30965# por_dig_0.net1 dvss.t2156 dvss.t2155 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.10025 ps=0.985 w=0.42 l=0.15
X1546 dvdd.t1697 dvss.t2298 dvdd.t1696 dvdd.t1695 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1547 a_38956_32339# por_dig_0.cnt_st\[2\] dvdd.t1371 dvdd.t1370 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.31245 ps=1.68 w=0.42 l=0.15
X1548 a_35100_32339# por_dig_0.net27 dvss.t2073 dvss.t2072 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.07035 ps=0.755 w=0.42 l=0.15
X1549 a_22047_21859# a_21622_21903# dvss.t1100 dvss.t1099 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X1550 por_ana_0.comparator_1.vnn.t19 por_ana_0.comparator_1.vpp.t59 avdd.t415 avdd.t403 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1551 dvdd.t968 por_ana_0.sky130_fd_sc_hd__inv_4_4.Y por.t26 dvdd.t967 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1552 a_34026_24707# a_33926_24619# dvss.t512 dvss.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X1553 a_34098_30707# por_dig_0.clknet_0_osc_ck.t38 dvdd.t1457 dvdd.t1456 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1554 dvdd.t1699 dvss.t2299 dvdd.t1698 dvdd.t1522 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X1555 dvdd.t741 por_dig_0.net7.t13 a_33326_28263# dvdd.t740 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.135 ps=1.27 w=1 l=0.15
X1556 a_35958_31519# a_35740_31277# dvdd.t1094 dvdd.t1093 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X1557 avdd.t87 avdd.t86 avdd.t87 avdd.t33 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=8
X1558 a_35293_30189# a_34212_30189# a_34946_30431# dvdd.t1082 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X1559 dvss.t123 a_39510_31251# por_dig_0._044_ dvss.t122 sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X1560 avdd.t537 por_ana_0.comparator_1.n1.t12 por_ana_0.dcomp3v3 avdd.t536 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X1561 dvss.t479 a_29802_22973# a_31009_22637# dvss.t478 sky130_fd_pr__nfet_g5v0d10v5 ad=0.121875 pd=1.075 as=0.19875 ps=2.03 w=0.75 l=0.5
X1562 a_35859_36717# por_dig_0.net23.t15 dvss.t880 dvss.t879 sky130_fd_pr__nfet_01v8 ad=0.095875 pd=0.945 as=0.17225 ps=1.83 w=0.65 l=0.15
X1563 a_37789_31821# por_dig_0._032_ a_37616_32141# dvss.t299 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X1564 avdd.t383 por_ana_0.ibias_gen_0.vp.t9 por_ana_0.comparator_0.ibias.t2 avdd.t382 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X1565 a_35529_33819# a_35092_33427# dvdd.t329 dvdd.t328 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X1566 a_34486_33453# por_dig_0.net22.t14 dvss.t1175 dvss.t1174 sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112125 ps=0.995 w=0.65 l=0.15
X1567 a_36844_35463# a_36494_35091# a_36749_35451# dvdd.t874 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X1568 avdd.t85 avdd.t84 avdd.t85 avdd.t13 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=8
X1569 por_ana_0.rstring_mux_0.vtrip1.t7 por_ana_0.rstring_mux_0.vtrip2.t5 avss.t287 sky130_fd_pr__res_xhigh_po_1p41 l=35
X1570 dvss.t343 por_ana_0.sky130_fd_sc_hd__inv_4_1.Y porb.t9 dvss.t342 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1571 a_37062_35059# a_36844_35463# dvss.t749 dvss.t748 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X1572 por_ana_0.comparator_0.vm.t3 por_ana_0.comparator_0.vm.t2 avss.t349 avss.t100 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1573 dvdd.t1702 dvss.t2300 dvdd.t1701 dvdd.t1700 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1574 dvss.t1139 por_ana_0.sky130_fd_sc_hd__inv_4_4.Y por.t1 dvss.t1138 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1575 por_ana_0.rstring_mux_0.otrip_decoded_avdd[7] a_28897_24371# avdd.t319 avdd.t317 sky130_fd_pr__pfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.24375 ps=1.825 w=1.5 l=0.5
X1576 a_37580_34375# a_37064_34003# a_37485_34363# dvss.t1271 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X1577 avss.t403 por_ana_0.ibias_gen_0.vn1.t13 por_ana_0.ibias_gen_0.vp1.t6 avss.t396 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=8
X1578 por_ana_0.comparator_0.vinn.t31 por_ana_0.rstring_mux_0.vtrip_decoded_b_avdd[1] por_ana_0.rstring_mux_0.vtrip1.t6 avdd.t465 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X1579 por_ana_0.rstring_mux_0.vtrip1.t2 por_ana_0.rstring_mux_0.otrip_decoded_avdd[1] vin.t12 avss.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X1580 dvdd.t1704 dvss.t2301 dvdd.t1703 dvdd.t1561 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1581 por_ana_0.ibias_gen_0.vp.t6 por_ana_0.rstring_mux_0.ena.t8 avdd.t612 avdd.t611 sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=2
X1582 avss.t342 por_ana_0.ibias_gen_0.isrc_sel.t6 por_ana_0.ibias_gen_0.vn0.t18 avss.t341 sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=2
X1583 por_ana_0.comparator_0.vpp.t38 por_ana_0.comparator_0.vnn.t54 avdd.t369 avdd.t191 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1584 avdd.t299 a_21354_24707# a_22561_24371# avdd.t298 sky130_fd_pr__pfet_g5v0d10v5 ad=0.24375 pd=1.825 as=0.3975 ps=3.53 w=1.5 l=0.5
X1585 dvss.t81 a_36122_30341# por_dig_0.net29 dvss.t80 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X1586 dvss.t1615 dvss.t1613 a_29702_24619# dvss.t1614 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X1587 a_15886_35244# a_15508_27844# avss.t159 sky130_fd_pr__res_xhigh_po_1p41 l=35
X1588 a_34378_35629# por_dig_0.cnt_por\[2\] a_34282_35629# dvss.t1576 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1589 por_ana_0.comparator_0.vpp.t1 por_ana_0.comparator_0.vpp.t0 avdd.t192 avdd.t191 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1590 por_ana_0.rstring_mux_0.vtrip5.t1 por_ana_0.rstring_mux_0.vtrip4.t0 avss.t160 sky130_fd_pr__res_xhigh_po_1p41 l=35
X1591 a_36749_35451# por_dig_0._006_ dvss.t625 dvss.t624 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X1592 por_dig_0.cnt_por\[5\] a_33720_33213# dvss.t743 dvss.t742 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X1593 a_31717_30189# a_31651_30341# por_dig_0.net10 dvss.t1168 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1594 avdd.t83 avdd.t82 avdd.t83 avdd.t33 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=8
X1595 dvss.t1811 dvdd.t1865 dvss.t1810 dvss.t1797 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1596 a_33364_36173# por_dig_0.net24 dvdd.t343 dvdd.t342 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X1597 avdd.t81 avdd.t79 avdd.t80 avdd.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=8
X1598 dvss.t1809 dvdd.t1866 dvss.t1808 dvss.t1737 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X1599 por_ana_0.comparator_0.vnn.t27 por_ana_0.comparator_0.vinn.t57 por_ana_0.comparator_0.vt.t8 por_ana_0.comparator_0.vt.t3 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1600 a_36564_32339# por_dig_0.net20.t6 dvdd.t1427 dvdd.t1426 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.1625 ps=1.325 w=1 l=0.15
X1601 por_ana_0.comparator_0.vt.t29 avss.t426 por_ana_0.comparator_0.vnn.t19 por_ana_0.comparator_0.vt.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=8
X1602 dvdd.t811 por_dig_0.cnt_st\[3\] a_39579_30849# dvdd.t810 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X1603 a_38131_31099# por_dig_0.net25 dvss.t955 dvss.t954 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X1604 por_ana_0.comparator_1.vn.t2 por_ana_0.comparator_1.ena_b por_ana_0.ibias_gen_0.ibias0.t2 avdd.t460 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X1605 dvss.t2095 otrip[1].t3 a_33971_28557# dvss.t2094 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X1606 a_37751_31251# por_dig_0._045_ dvss.t1391 dvss.t1390 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.1359 ps=1.1 w=0.42 l=0.15
X1607 avdd.t78 avdd.t77 avdd.t78 avdd.t13 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=8
X1608 a_18920_13935# a_19298_6535# avss.t161 sky130_fd_pr__res_xhigh_po_1p41 l=35
X1609 por_dig_0._032_ por_dig_0._031_ dvss.t172 dvss.t171 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1610 dvdd.t555 por_ana_0.schmitt_trigger_0.m.t16 por_ana_0.schmitt_trigger_0.out.t2 dvdd.t554 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X1611 por_ana_0.comparator_0.vt.t44 vbg_1v2.t27 por_ana_0.comparator_0.vpp.t25 por_ana_0.comparator_0.vt.t36 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1612 avdd.t506 a_34719_23593# a_34026_24707# avdd.t505 sky130_fd_pr__pfet_g5v0d10v5 ad=0.2142 pd=1.99 as=0.2142 ps=1.99 w=0.42 l=1
X1613 a_21944_13935# a_22322_6535# avss.t162 sky130_fd_pr__res_xhigh_po_1p41 l=35
X1614 por_ana_0.rc_osc_0.n.t0 por_ana_0.rc_osc_0.m dvss.t530 dvss.t529 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X1615 por_ana_0.ibias_gen_0.ve.t4 por_ana_0.ibias_gen_0.vn0.t4 por_ana_0.ibias_gen_0.vn0.t5 avss.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X1616 a_24159_23593# a_23734_23637# dvss.t1129 dvss.t1128 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X1617 avdd.t659 a_25595_33708# a_26802_33372# avdd.t445 sky130_fd_pr__pfet_g5v0d10v5 ad=0.24375 pd=1.825 as=0.3975 ps=3.53 w=1.5 l=0.5
X1618 dvdd.t1706 dvss.t2302 dvdd.t1705 dvdd.t1522 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1619 dvdd.t189 por_ana_0.sky130_fd_sc_hd__inv_4_1.A por_ana_0.sky130_fd_sc_hd__inv_4_1.Y dvdd.t188 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1620 a_37409_35463# a_36328_35091# a_37062_35059# dvdd.t872 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X1621 dvdd.t778 osc_ck.t13 a_34387_32909# dvdd.t777 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1622 dvdd.t1125 por_dig_0.net3 por_dig_0.net9 dvdd.t1124 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1623 a_35122_33997# por_dig_0._022_ dvdd.t310 dvdd.t309 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X1624 dvdd.t117 a_34387_32909# por_dig_0.clknet_0_osc_ck.t23 dvdd.t116 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1625 a_35583_34541# por_dig_0.clknet_0_osc_ck.t39 dvss.t2133 dvss.t2132 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1626 por_dig_0._025_ por_dig_0.cnt_por\[6\] dvdd.t390 dvdd.t389 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X1627 por_dig_0._026_ por_dig_0.net22.t15 dvdd.t986 dvdd.t985 sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.39 as=0.182 ps=1.92 w=0.7 l=0.15
X1628 por_dig_0.clknet_1_1__leaf_osc_ck.t7 a_35583_34541# dvss.t580 dvss.t579 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.05775 ps=0.695 w=0.42 l=0.15
X1629 por_ana_0.comparator_0.vinn.t14 avss.t84 por_ana_0.comparator_0.vinn.t14 avss.t85 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=0.6
X1630 por_ana_0.rstring_mux_0.vtrip1.t0 por_ana_0.rstring_mux_0.otrip_decoded_b_avdd[1] vin.t10 avdd.t214 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X1631 a_35390_31277# a_35224_31277# dvdd.t1091 dvdd.t1090 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1632 por_dig_0.clknet_0_osc_ck.t7 a_34387_32909# dvss.t149 dvss.t148 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1633 dvdd.t265 por_dig_0.cnt_por\[8\] a_35000_31795# dvdd.t264 sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=1.61 as=0.2175 ps=1.435 w=1 l=0.15
X1634 dvdd.t1709 dvss.t2303 dvdd.t1708 dvdd.t1707 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1635 a_37504_33819# por_dig_0.net25 dvdd.t837 dvdd.t836 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X1636 por_ana_0.rstring_mux_0.otrip_decoded_b_avdd[2] por_ana_0.rstring_mux_0.otrip_decoded_avdd[2] avss.t4 avss.t3 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X1637 dvss.t1216 a_31776_29864# por_dig_0.net2 dvss.t1215 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X1638 a_39718_33605# por_dig_0.cnt_st\[1\] dvss.t600 dvss.t599 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.10025 ps=0.985 w=0.42 l=0.15
X1639 a_37614_32883# a_37396_33287# dvdd.t796 dvdd.t795 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X1640 dvss.t312 a_31914_22973# a_33121_22637# dvss.t311 sky130_fd_pr__nfet_g5v0d10v5 ad=0.121875 pd=1.075 as=0.19875 ps=2.03 w=0.75 l=0.5
X1641 a_37596_30555# por_dig_0.net25 dvdd.t835 dvdd.t834 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X1642 avdd.t76 avdd.t74 avdd.t75 avdd.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=8
X1643 dvdd.t419 por_dig_0.clknet_1_0__leaf_osc_ck.t40 a_36696_30739# dvdd.t418 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1644 a_35024_35629# por_dig_0.cnt_por\[1\] por_dig_0._034_.t5 dvss.t1401 sky130_fd_pr__nfet_01v8 ad=0.234 pd=2.02 as=0.08775 ps=0.92 w=0.65 l=0.15
X1645 dvss.t672 a_30070_21903# a_30495_21859# dvss.t671 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X1646 a_31776_29864# force_ena_rc_osc.t3 dvss.t2012 dvss.t177 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1647 por_dig_0._005_ a_35704_35124# dvdd.t1196 dvdd.t1195 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.15835 ps=1.395 w=1 l=0.15
X1648 dvdd.t998 por_ana_0.vl por_ana_0.sky130_fd_sc_hd__inv_4_3.Y dvdd.t997 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1649 a_25578_24707# a_25478_24619# dvss.t1482 dvss.t1481 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X1650 a_39354_32365# por_dig_0.cnt_st\[0\] a_39248_32365# dvss.t1331 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0798 ps=0.8 w=0.42 l=0.15
X1651 dvdd.t535 por_dig_0.cnt_por\[0\].t14 a_35918_35124# dvdd.t534 sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.07665 ps=0.785 w=0.42 l=0.15
X1652 pwup_filt.t5 por_ana_0.sky130_fd_sc_hd__inv_4_0.Y dvss.t238 dvss.t237 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1653 dvss.t1807 dvdd.t1867 dvss.t1806 dvss.t1805 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X1654 dvdd.t571 a_37409_35463# a_37584_35389# dvdd.t570 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X1655 dvdd.t481 a_35583_34541# por_dig_0.clknet_1_1__leaf_osc_ck.t21 dvdd.t480 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1656 por_ana_0.sky130_fd_sc_hvl__inv_1_0.A a_26802_33372# dvss.t1038 dvss.t1037 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.121875 ps=1.075 w=0.75 l=0.5
X1657 dvdd.t1516 a_32535_28013# a_32641_28013# dvdd.t1515 sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X1658 avdd.t514 a_23466_24707# a_24673_24371# avdd.t453 sky130_fd_pr__pfet_g5v0d10v5 ad=0.24375 pd=1.825 as=0.3975 ps=3.53 w=1.5 l=0.5
X1659 dvdd.t1004 a_39732_31829# startup_timed_out.t3 dvdd.t1003 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X1660 a_38957_32883# por_dig_0._029_ a_39177_33229# dvss.t2027 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X1661 avss.t83 avss.t80 avss.t82 avss.t81 sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0 ps=0 w=5 l=8
X1662 por_ana_0.dcomp3v3uv por_ana_0.comparator_0.n1.t11 avss.t275 avss.t274 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X1663 por_ana_0.rstring_mux_0.otrip_decoded_b_avdd[5] por_ana_0.rstring_mux_0.otrip_decoded_avdd[5] avdd.t467 avdd.t466 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X1664 dvss.t236 por_ana_0.sky130_fd_sc_hd__inv_4_0.Y pwup_filt.t4 dvss.t235 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1665 dvss.t147 a_34387_32909# por_dig_0.clknet_0_osc_ck.t6 dvss.t146 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X1666 dvdd.t864 a_38146_31429# por_dig_0.net34 dvdd.t863 sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.26 ps=2.52 w=1 l=0.15
X1667 dvdd.t1006 por_dig_0._040_ a_39094_32909# dvdd.t1005 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X1668 avss.t277 por_ana_0.comparator_0.n1.t12 por_ana_0.dcomp3v3uv avss.t276 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X1669 dvdd.t575 por_dig_0.net11 a_38444_28013# dvdd.t574 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X1670 a_34856_36493# por_dig_0.cnt_por\[0\].t15 a_34762_36493# dvss.t641 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X1671 por.t25 por_ana_0.sky130_fd_sc_hd__inv_4_4.Y dvdd.t966 dvdd.t965 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1672 por_ana_0.comparator_0.vinn.t2 avdd.t72 por_ana_0.comparator_0.vinn.t2 avdd.t73 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=0.6
X1673 dvss.t1804 dvdd.t1868 dvss.t1803 dvss.t1729 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1674 dvdd.t649 a_37062_35059# a_36952_35085# dvdd.t648 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X1675 dvss.t953 por_dig_0.net25 a_37750_30189# dvss.t952 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X1676 por_ana_0.comparator_0.vpp.t39 por_ana_0.comparator_0.vnn.t55 avdd.t370 avdd.t191 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1677 vin.t17 avss.t78 vin.t17 avss.t79 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=0.6
X1678 por_dig_0.force_pdnb a_31413_29075# dvdd.t1518 dvdd.t668 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X1679 dvdd.t327 a_35092_33427# por_dig_0.cnt_por\[4\] dvdd.t309 sky130_fd_pr__pfet_01v8_hvt ad=0.3012 pd=2.66 as=0.26 ps=2.52 w=1 l=0.15
X1680 a_26271_23593# a_25846_23637# dvss.t366 dvss.t365 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X1681 a_36006_33453# por_dig_0.net24 dvss.t431 dvss.t430 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1346 ps=1.15 w=0.42 l=0.15
X1682 por_ana_0.comparator_0.vnn.t46 por_ana_0.comparator_0.vnn.t45 avdd.t361 avdd.t182 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1683 avdd.t71 avdd.t70 avdd.t71 avdd.t33 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=8
X1684 por_dig_0.otrip_decoded[1] a_32701_28531# dvdd.t3 dvdd.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X1685 a_36659_31277# por_dig_0.net25 dvss.t951 dvss.t950 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X1686 dvss.t1325 otrip[0].t2 a_32039_28013# dvss.t677 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X1687 a_33804_31251# por_dig_0.cnt_por\[8\] a_34235_31277# dvss.t316 sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.11375 ps=1 w=0.65 l=0.15
X1688 por_dig_0._035_ por_dig_0.cnt_por\[5\] a_34738_32141# dvss.t2083 sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.10725 ps=0.98 w=0.65 l=0.15
X1689 a_39728_31527# por_dig_0._030_ a_39510_31251# dvdd.t1504 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.26 ps=2.52 w=1 l=0.15
X1690 por_ana_0.rstring_mux_0.otrip_decoded_avdd[1] a_22561_24371# dvss.t1306 dvss.t1305 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.121875 ps=1.075 w=0.75 l=0.5
X1691 avdd.t640 por_ana_0.comparator_1.vnn.t54 por_ana_0.comparator_1.vpp.t24 avdd.t392 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1692 por_dig_0.net11 por_dig_0.net5.t9 a_35770_29351# dvdd.t668 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1693 a_15140_13935# a_15518_6535# avss.t163 sky130_fd_pr__res_xhigh_po_1p41 l=35
X1694 a_33269_31111# a_32188_30739# a_32922_30707# dvdd.t817 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X1695 dvdd.t1060 a_40247_23627# por_ana_0.vl dvdd.t1058 sky130_fd_pr__pfet_01v8_hvt ad=0.1568 pd=1.4 as=0.2968 ps=2.77 w=1.12 l=0.15
X1696 a_37611_31277# por_dig_0._042_ dvss.t306 dvss.t305 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.258375 ps=1.445 w=0.65 l=0.15
X1697 avdd.t69 avdd.t68 avdd.t69 avdd.t13 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=8
X1698 a_36376_28789# por_dig_0.net7.t14 dvdd.t743 dvdd.t742 sky130_fd_pr__pfet_01v8_hvt ad=0.074375 pd=0.815 as=0.142225 ps=1.335 w=0.42 l=0.15
X1699 dvss.t358 a_34026_22973# a_35233_22637# dvss.t357 sky130_fd_pr__nfet_g5v0d10v5 ad=0.121875 pd=1.075 as=0.19875 ps=2.03 w=0.75 l=0.5
X1700 a_38162_30189# a_36972_30189# a_38053_30189# dvss.t26 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1701 dvss.t678 por_dig_0.net11 a_38444_28013# dvss.t677 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X1702 dvss.t1118 a_32182_21903# a_32607_21859# dvss.t1117 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X1703 a_14374_35244# a_14752_27844# avss.t164 sky130_fd_pr__res_xhigh_po_1p41 l=35
X1704 dvss.t1802 dvdd.t1869 dvss.t1801 dvss.t1800 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1705 a_33550_32141# por_dig_0.cnt_por\[8\] a_33466_32141# dvss.t315 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X1706 por_ana_0.sky130_fd_sc_hd__inv_4_4.Y por_dig_0.por_unbuf.t14 dvss.t810 dvss.t809 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1707 a_16652_13935# a_16274_6535# avss.t165 sky130_fd_pr__res_xhigh_po_1p41 l=35
X1708 por_dig_0.clknet_1_0__leaf_osc_ck.t24 a_34098_30707# dvdd.t165 dvdd.t164 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1709 a_34098_30707# por_dig_0.clknet_0_osc_ck.t40 dvdd.t1459 dvdd.t1458 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1710 avdd.t551 por_ana_0.ibias_gen_0.vp0.t3 por_ana_0.ibias_gen_0.vp0.t4 avdd.t550 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X1711 por_ana_0.ibias_gen_0.vstart.t1 vbg_1v2.t28 por_ana_0.ibias_gen_0.vn0.t14 avss.t150 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=0.6
X1712 dvss.t1799 dvdd.t1870 dvss.t1798 dvss.t1797 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1713 dvss.t933 por_dig_0.cnt_st\[3\] a_39497_30849# dvss.t932 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X1714 avss.t17 por_ana_0.comparator_1.n1.t13 por_ana_0.dcomp3v3 avss.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X1715 a_33326_28263# por_dig_0.net6 a_33242_28263# dvdd.t675 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1716 dvss.t1796 dvdd.t1871 dvss.t1795 dvss.t1794 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X1717 dvdd.t1443 por_dig_0.net5.t10 a_32358_28013# dvdd.t1442 sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X1718 dvss.t812 por_dig_0.por_unbuf.t15 por_ana_0.sky130_fd_sc_hd__inv_4_4.Y dvss.t811 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1719 vin.t5 avdd.t66 vin.t5 avdd.t67 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=0.6
X1720 dvss.t1612 dvss.t1610 a_31814_22885# dvss.t1611 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X1721 avdd.t303 a_25578_24707# a_26785_24371# avdd.t302 sky130_fd_pr__pfet_g5v0d10v5 ad=0.24375 pd=1.825 as=0.3975 ps=3.53 w=1.5 l=0.5
X1722 avdd.t65 avdd.t63 avdd.t64 avdd.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=8
X1723 a_34175_36539# por_dig_0.net24 dvss.t429 dvss.t428 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X1724 a_36278_35629# a_36234_35871# a_36112_35629# dvss.t1985 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X1725 dvss.t1964 por_dig_0._025_ a_33097_34317# dvss.t1963 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X1726 dvdd.t745 por_dig_0.net7.t15 a_34934_28013# dvdd.t744 sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X1727 dvdd.t13 a_31932_31419# a_31893_31545# dvdd.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1728 a_37504_32909# por_dig_0.net24 dvdd.t341 dvdd.t340 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X1729 a_38956_32339# por_dig_0.cnt_st\[0\] dvdd.t1112 dvdd.t1111 sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.0777 ps=0.79 w=0.42 l=0.15
X1730 por_dig_0.net18 a_35776_28013# dvdd.t1214 dvdd.t632 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X1731 por_dig_0.otrip_decoded[4] a_34265_27987# dvdd.t1133 dvdd.t1132 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X1732 a_31413_29619# por_dig_0.net10 dvdd.t523 dvdd.t522 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X1733 a_35390_31277# a_35224_31277# dvss.t1287 dvss.t1286 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1734 por_dig_0.cnt_por\[0\].t7 a_36756_35603# dvdd.t469 dvdd.t468 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1735 a_34842_35451# por_dig_0.cnt_por\[0\].t16 a_34754_35451# dvss.t642 sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
X1736 avss.t167 a_38954_6535# avss.t166 sky130_fd_pr__res_xhigh_po_1p41 l=35
X1737 por_dig_0._011_ por_dig_0._023_ a_35122_33997# dvdd.t805 sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.39 as=0.105 ps=1.21 w=1 l=0.15
X1738 por_ana_0.comparator_0.vpp.t26 vbg_1v2.t29 por_ana_0.comparator_0.vt.t43 por_ana_0.comparator_0.vt.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1739 a_33242_33275# a_33198_32883# a_33076_33287# dvss.t1392 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X1740 porb_h.t27 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.t25 avss.t187 avss.t186 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X1741 a_33256_36551# a_32906_36179# a_33161_36539# dvdd.t614 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X1742 por_dig_0._015_ a_34496_29645# a_34746_29645# dvdd.t70 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.26 ps=2.52 w=1 l=0.15
X1743 a_37392_31251# a_37751_31251# a_37528_31527# dvdd.t1053 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X1744 a_20422_35244# a_20800_27844# avss.t168 sky130_fd_pr__res_xhigh_po_1p41 l=35
X1745 dvdd.t1201 a_37952_31037# a_37939_30733# dvdd.t1200 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X1746 dvdd.t891 por_dig_0.force_pdnb a_38150_22885# dvdd.t890 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X1747 por_ana_0.rstring_mux_0.otrip_decoded_avdd[5] a_26785_24371# dvss.t1320 dvss.t1319 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.121875 ps=1.075 w=0.75 l=0.5
X1748 a_37106_35451# a_37062_35059# a_36940_35463# dvss.t750 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X1749 avdd.t624 por_ana_0.ibias_gen_0.vp1.t12 por_ana_0.ibias_gen_0.vp1.t13 avdd.t623 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X1750 a_34357_33427# por_dig_0.cnt_por\[4\] a_34580_33453# dvss.t1548 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1751 a_21354_22973# a_21254_22885# dvss.t1069 dvss.t1068 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X1752 dvdd.t1467 isrc_sel.t3 a_38150_24619# dvdd.t1466 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X1753 por_ana_0.schmitt_trigger_0.out.t1 por_ana_0.schmitt_trigger_0.m.t17 dvdd.t557 dvdd.t556 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X1754 por_dig_0.net32 a_34116_31821# dvss.t775 dvss.t774 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X1755 por_dig_0.cnt_por\[10\] a_36480_31251# dvss.t1508 dvss.t1507 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X1756 a_32885_33275# por_dig_0._010_ dvdd.t1328 dvdd.t1327 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X1757 a_34175_35451# por_dig_0.net24 dvss.t427 dvss.t426 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X1758 por_ana_0.ibias_gen_0.vp0.t6 por_ana_0.ibias_gen_0.vn0.t20 por_ana_0.ibias_gen_0.vr.t2 avss.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X1759 dvdd.t1712 dvss.t2304 dvdd.t1711 dvdd.t1710 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1760 a_32088_33690# a_31893_33721# a_32398_33453# dvss.t476 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.1401 ps=1.1 w=0.36 l=0.15
X1761 dvss.t133 a_36138_22973# a_37345_22637# dvss.t132 sky130_fd_pr__nfet_g5v0d10v5 ad=0.121875 pd=1.075 as=0.19875 ps=2.03 w=0.75 l=0.5
X1762 dvdd.t780 osc_ck.t14 a_34387_32909# dvdd.t779 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1763 por_ana_0.rstring_mux_0.otrip_decoded_b_avdd[7] por_ana_0.rstring_mux_0.otrip_decoded_avdd[7] avss.t228 avss.t227 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X1764 dvdd.t1715 dvss.t2305 dvdd.t1714 dvdd.t1713 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1765 a_35583_34541# por_dig_0.clknet_0_osc_ck.t41 dvss.t2135 dvss.t2134 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X1766 avdd.t428 a_22047_21859# a_21354_22973# avdd.t427 sky130_fd_pr__pfet_g5v0d10v5 ad=0.2142 pd=1.99 as=0.2142 ps=1.99 w=0.42 l=1
X1767 por_ana_0.schmitt_trigger_0.m.t10 por_ana_0.schmitt_trigger_0.out.t10 dvss.t820 dvss.t819 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X1768 dvdd.t988 por_dig_0.net22.t16 por_dig_0._025_ dvdd.t987 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1769 por_dig_0.clknet_0_osc_ck.t5 a_34387_32909# dvss.t145 dvss.t144 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1770 dvdd.t421 por_dig_0.clknet_1_0__leaf_osc_ck.t41 a_35224_31277# dvdd.t420 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1771 avdd.t416 por_ana_0.comparator_1.vpp.t60 por_ana_0.comparator_1.vnn.t18 avdd.t401 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1772 dvss.t1793 dvdd.t1872 dvss.t1792 dvss.t1787 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1773 dvdd.t1218 a_37800_28013# por_dig_0.otrip_decoded[3].t3 dvdd.t1217 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X1774 a_38936_32159# por_dig_0.cnt_st\[4\] dvdd.t1242 dvdd.t1241 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X1775 a_7079_22912# a_6701_15512# avss.t27 sky130_fd_pr__res_xhigh_po_1p41 l=35
X1776 avdd.t589 a_31914_24707# a_32607_23593# avdd.t588 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.1365 ps=1.49 w=0.42 l=1
X1777 a_31526_31827# a_31360_31827# dvdd.t22 dvdd.t21 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1778 por_ana_0.comparator_0.vpp.t40 por_ana_0.comparator_0.vnn.t56 avdd.t371 avdd.t191 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1779 dvss.t1609 dvss.t1607 a_33926_22885# dvss.t1608 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X1780 dvdd.t1717 dvss.t2306 dvdd.t1716 dvdd.t1522 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X1781 por_ana_0.comparator_1.vpp.t39 vin.t58 por_ana_0.comparator_1.vt.t27 por_ana_0.comparator_1.vt.t18 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1782 avss.t77 avss.t76 avss.t77 avss.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=8
X1783 a_31615_31529# a_31932_31419# a_31890_31277# dvss.t24 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0669 ps=0.75 w=0.36 l=0.15
X1784 por_dig_0._034_.t4 por_dig_0.cnt_por\[1\] a_35024_35629# dvss.t1400 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1785 por_ana_0.ibias_gen_0.ve.t0 avss.t74 avss.t75 avss.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=4
X1786 a_34762_36493# por_dig_0.net23.t16 dvss.t882 dvss.t881 sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112125 ps=0.995 w=0.65 l=0.15
X1787 dvdd.t1461 por_dig_0.clknet_0_osc_ck.t42 a_35583_34541# dvdd.t1460 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1788 por_dig_0.por_unbuf.t3 a_36381_36691# dvdd.t1475 dvdd.t1474 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X1789 dvdd.t479 a_35583_34541# por_dig_0.clknet_1_1__leaf_osc_ck.t20 dvdd.t478 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1790 por_ana_0.dcomp3v3uv por_ana_0.comparator_0.n1.t13 avdd.t486 avdd.t485 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X1791 por_ana_0.comparator_1.vpp.t40 vin.t59 por_ana_0.comparator_1.vt.t26 por_ana_0.comparator_1.vt.t18 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1792 a_33465_35629# por_dig_0._053_ a_33162_35603# dvss.t1998 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.089375 ps=0.925 w=0.65 l=0.15
X1793 dvdd.t537 por_dig_0.cnt_por\[0\].t17 a_35450_35124# dvdd.t536 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.1176 ps=1.4 w=0.42 l=0.15
X1794 a_36831_21859# a_36406_21903# dvss.t1312 dvss.t1311 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X1795 a_38053_30189# a_37138_30189# a_37706_30431# dvss.t2036 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X1796 por_ana_0.comparator_0.vt.t28 avss.t427 por_ana_0.comparator_0.vnn.t18 por_ana_0.comparator_0.vt.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=8
X1797 por_dig_0.net22.t1 a_36380_33971# dvss.t1021 dvss.t1020 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1798 a_35330_33453# a_35295_33705# a_35092_33427# dvss.t1393 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.1092 ps=1.36 w=0.42 l=0.15
X1799 dvss.t2118 por_dig_0.net5.t11 a_35933_28917# dvss.t2117 sky130_fd_pr__nfet_01v8 ad=0.122275 pd=1.08 as=0.05355 ps=0.675 w=0.42 l=0.15
X1800 dvdd.t307 por_dig_0.net30 a_33934_29645# dvdd.t70 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1801 por_ana_0.comparator_1.vn.t4 por_ana_0.comparator_1.vn.t3 avss.t289 avss.t288 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1802 dvdd.t477 a_35583_34541# por_dig_0.clknet_1_1__leaf_osc_ck.t19 dvdd.t476 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X1803 avdd.t62 avdd.t61 avdd.t62 avdd.t13 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=8
X1804 a_36308_13935# a_36686_6535# avss.t169 sky130_fd_pr__res_xhigh_po_1p41 l=35
X1805 dvdd.t1357 por_ana_0.rc_osc_0.n.t9 osc_ck.t4 dvdd.t1356 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X1806 dvdd.t371 a_33821_36551# a_33996_36477# dvdd.t370 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X1807 a_32616_32125# a_32441_32199# a_32795_32187# dvss.t1304 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X1808 startup_timed_out.t2 a_39732_31829# dvdd.t1002 dvdd.t1001 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X1809 a_34633_30189# por_dig_0._014_ dvss.t2172 dvss.t2171 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X1810 por_dig_0.net13 por_dig_0.net7.t16 dvss.t858 dvss.t857 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10025 ps=0.985 w=0.65 l=0.15
X1811 por_ana_0.ibias_gen_0.vr.t4 a_8969_15512# avss.t27 sky130_fd_pr__res_xhigh_po_1p41 l=35
X1812 a_37961_33453# a_36880_33453# a_37614_33695# dvdd.t650 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X1813 avdd.t60 avdd.t59 avdd.t60 avdd.t13 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=8
X1814 a_25578_22973# a_25478_22885# dvss.t1562 dvss.t1561 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X1815 dvdd.t1388 a_38957_32883# por_dig_0._001_ dvdd.t1387 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.15
X1816 por_dig_0._006_ por_dig_0._048_ a_36328_36493# dvss.t1110 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1817 por_ana_0.comparator_0.vt.t27 avss.t428 por_ana_0.comparator_0.vnn.t17 por_ana_0.comparator_0.vt.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=8
X1818 por_ana_0.rstring_mux_0.otrip_decoded_avdd[7] a_28897_24371# dvss.t767 dvss.t766 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.121875 ps=1.075 w=0.75 l=0.5
X1819 a_37117_31099# por_dig_0._004_ dvdd.t1008 dvdd.t1007 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X1820 a_36112_35629# a_35666_35629# a_36016_35629# dvss.t619 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X1821 por_dig_0._015_ por_dig_0._028_ a_34746_29965# dvss.t369 sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.08775 ps=0.92 w=0.65 l=0.15
X1822 dvss.t661 a_21354_24707# a_22561_24371# dvss.t660 sky130_fd_pr__nfet_g5v0d10v5 ad=0.121875 pd=1.075 as=0.19875 ps=2.03 w=0.75 l=0.5
X1823 por_ana_0.comparator_1.vpp.t41 vin.t60 por_ana_0.comparator_1.vt.t25 por_ana_0.comparator_1.vt.t18 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1824 dvdd.t933 por_dig_0.cnt_por\[7\] por_dig_0._035_ dvdd.t932 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1825 dvdd.t674 por_dig_0.net6 a_34290_28557# dvdd.t673 sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X1826 por_ana_0.rstring_mux_0.vtrip1.t8 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[1] por_ana_0.comparator_0.vinn.t38 avss.t315 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X1827 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[4].t1 a_35233_22637# dvss.t2035 dvss.t2034 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.121875 ps=1.075 w=0.75 l=0.5
X1828 por.t24 por_ana_0.sky130_fd_sc_hd__inv_4_4.Y dvdd.t964 dvdd.t963 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1829 avdd.t360 por_ana_0.comparator_0.vnn.t43 por_ana_0.comparator_0.vnn.t44 avdd.t180 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1830 a_31016_13935# a_30638_6535# avss.t170 sky130_fd_pr__res_xhigh_po_1p41 l=35
X1831 dvdd.t163 a_34098_30707# por_dig_0.clknet_1_0__leaf_osc_ck.t23 dvdd.t162 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1832 a_25863_32638# a_25495_33620# dvdd.t1205 dvdd.t1204 sky130_fd_pr__pfet_01v8_hvt ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X1833 dvss.t266 a_38518_21903# a_38943_21859# dvss.t265 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X1834 por_ana_0.comparator_1.vpp.t42 vin.t61 por_ana_0.comparator_1.vt.t24 por_ana_0.comparator_1.vt.t18 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1835 dvss.t23 a_31932_31419# a_31893_31545# dvss.t22 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1836 dvdd.t1186 a_31802_32909# a_31908_32909# dvdd.t1185 sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.5
X1837 a_31413_29619# por_dig_0.net10 dvss.t623 dvss.t622 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X1838 a_36016_35629# a_35500_35629# a_35921_35629# dvss.t525 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X1839 a_37230_34003# a_37064_34003# dvss.t1270 dvss.t1269 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1840 a_31772_13935# a_32150_6535# avss.t171 sky130_fd_pr__res_xhigh_po_1p41 l=35
X1841 avdd.t305 a_24159_21859# a_23466_22973# avdd.t304 sky130_fd_pr__pfet_g5v0d10v5 ad=0.2142 pd=1.99 as=0.2142 ps=1.99 w=0.42 l=1
X1842 a_36952_35085# por_dig_0.net24 dvdd.t339 dvdd.t338 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X1843 dvdd.t1320 a_35768_33690# a_35699_33819# dvdd.t1319 sky130_fd_pr__pfet_01v8_hvt ad=0.2184 pd=2.2 as=0.12915 ps=1.185 w=0.84 l=0.15
X1844 a_38123_33819# a_37046_33453# a_37961_33453# dvdd.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X1845 por_ana_0.rc_osc_0.in dvss.t289 sky130_fd_pr__cap_mim_m3_2 l=30 w=30
X1846 a_38215_30555# a_37138_30189# a_38053_30189# dvdd.t1210 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X1847 avdd.t58 avdd.t56 avdd.t57 avdd.t3 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=8
X1848 por_ana_0.comparator_0.vpp.t46 avss.t429 avdd.t521 avdd.t520 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X1849 dvss.t2225 a_25595_33708# a_26802_33372# dvss.t2224 sky130_fd_pr__nfet_g5v0d10v5 ad=0.121875 pd=1.075 as=0.19875 ps=2.03 w=0.75 l=0.5
X1850 dvdd.t565 por_ana_0.schmitt_trigger_0.in.t9 por_ana_0.schmitt_trigger_0.m.t4 dvdd.t564 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X1851 dvss.t1791 dvdd.t1873 dvss.t1790 dvss.t1706 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1852 por_dig_0.clknet_1_0__leaf_osc_ck.t22 a_34098_30707# dvdd.t161 dvdd.t160 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1853 a_34295_34317# por_dig_0._019_ dvss.t2180 dvss.t2179 sky130_fd_pr__nfet_01v8 ad=0.095875 pd=0.945 as=0.17225 ps=1.83 w=0.65 l=0.15
X1854 avss.t189 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.t26 porb_h.t26 avss.t188 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X1855 a_39162_33453# a_38926_33453# dvdd.t623 dvdd.t622 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.5
X1856 dvss.t548 a_39417_31795# por_dig_0.net4 dvss.t547 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X1857 a_23734_21903# a_23366_22885# dvdd.t788 dvdd.t787 sky130_fd_pr__pfet_01v8_hvt ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X1858 a_31822_30849# por_dig_0.net19 a_31727_30849# dvdd.t1010 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.06825 ps=0.745 w=0.42 l=0.15
X1859 a_32918_32365# a_31728_32365# a_32809_32365# dvss.t692 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1860 a_33934_32365# por_dig_0._019_ dvss.t2178 dvss.t2177 sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112125 ps=0.995 w=0.65 l=0.15
X1861 a_33466_32141# por_dig_0.cnt_por\[10\] dvss.t1512 dvss.t1511 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1862 a_39077_31527# por_dig_0._032_ a_38986_31527# dvdd.t246 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.1525 ps=1.305 w=1 l=0.15
X1863 dvdd.t1445 por_dig_0.net5.t12 a_36376_28789# dvdd.t1444 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.074375 ps=0.815 w=0.42 l=0.15
X1864 dvss.t341 por_ana_0.sky130_fd_sc_hd__inv_4_1.Y porb.t8 dvss.t340 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1865 por_dig_0.cnt_por\[1\] a_37584_35389# dvss.t1015 dvss.t1014 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.2087 ps=2.02 w=0.65 l=0.15
X1866 a_23734_23637# a_23366_24619# dvdd.t1232 dvdd.t1231 sky130_fd_pr__pfet_01v8_hvt ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X1867 a_39497_30849# por_dig_0.net4 dvss.t90 dvss.t89 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1868 por_dig_0._033_ a_34672_35451# dvdd.t1026 dvdd.t1025 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.31245 ps=1.68 w=1 l=0.15
X1869 dvss.t425 por_dig_0.net24 a_37106_35451# dvss.t424 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X1870 a_32607_23593# a_32182_23637# dvss.t7 dvss.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X1871 dvdd.t595 por_dig_0.clknet_1_1__leaf_osc_ck.t37 a_32740_36179# dvdd.t594 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1872 por_ana_0.rstring_mux_0.vtrip1.t5 por_ana_0.rstring_mux_0.vtrip_decoded_b_avdd[1] por_ana_0.comparator_0.vinn.t30 avdd.t464 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X1873 vin.t16 avss.t72 vin.t16 avss.t73 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=0.6
X1874 a_38943_21859# a_38518_21903# dvss.t264 dvss.t263 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X1875 dvss.t753 a_37156_28013# por_dig_0.otrip_decoded[7].t1 dvss.t523 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X1876 dvdd.t1720 dvss.t2307 dvdd.t1719 dvdd.t1718 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1877 dvss.t314 a_36382_31795# por_dig_0.net20.t0 dvss.t313 sky130_fd_pr__nfet_01v8 ad=0.203125 pd=1.275 as=0.169 ps=1.82 w=0.65 l=0.15
X1878 dvdd.t1723 dvss.t2308 dvdd.t1722 dvdd.t1721 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1879 por_dig_0.net27 a_34852_31277# dvdd.t1394 dvdd.t1393 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X1880 porb.t7 por_ana_0.sky130_fd_sc_hd__inv_4_1.Y dvss.t339 dvss.t338 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1881 avdd.t553 por_ana_0.ibias_gen_0.vp0.t13 por_ana_0.ibias_gen_0.vn0.t0 avdd.t552 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X1882 a_27690_22973# a_27590_22885# dvss.t1373 dvss.t1372 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X1883 dvss.t2137 por_dig_0.clknet_0_osc_ck.t43 a_34098_30707# dvss.t2136 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1884 por_ana_0.comparator_0.vnn avss.t430 por_ana_0.comparator_0.vt.t26 por_ana_0.comparator_0.vt.t18 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=8
X1885 dvss.t212 a_32088_31514# a_32019_31643# dvss.t211 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0999 ps=0.985 w=0.64 l=0.15
X1886 avdd.t641 por_ana_0.comparator_1.vnn.t55 por_ana_0.comparator_1.vm.t1 avdd.t392 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1887 dvss.t503 por_dig_0.clknet_1_0__leaf_osc_ck.t42 a_35224_31277# dvss.t502 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1888 dvdd.t1160 por_dig_0.cnt_por\[1\] a_35592_36286# dvdd.t1159 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1889 dvdd.t115 a_34387_32909# por_dig_0.clknet_0_osc_ck.t22 dvdd.t114 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X1890 a_27690_22973# a_27590_22885# dvss.t1371 dvss.t1370 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X1891 a_32528_13935# a_32906_6535# avss.t172 sky130_fd_pr__res_xhigh_po_1p41 l=35
X1892 dvss.t1447 a_23466_24707# a_24673_24371# dvss.t1446 sky130_fd_pr__nfet_g5v0d10v5 ad=0.121875 pd=1.075 as=0.19875 ps=2.03 w=0.75 l=0.5
X1893 dvdd.t1446 por_dig_0.net5.t13 a_35774_28673# dvdd.t1438 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.074375 ps=0.815 w=0.42 l=0.15
X1894 dvdd.t1726 dvss.t2309 dvdd.t1725 dvdd.t1724 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
R1 dvss por_dig_0._137__26.LO sky130_fd_pr__res_generic_po w=0.48 l=0.045
X1895 por_dig_0.clknet_1_1__leaf_osc_ck.t6 a_35583_34541# dvss.t578 dvss.t577 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1896 a_32149_32365# por_dig_0._012_ dvss.t1436 dvss.t1435 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X1897 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[6].t1 a_37345_22637# dvss.t2086 dvss.t2085 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.121875 ps=1.075 w=0.75 l=0.5
X1898 avdd.t55 avdd.t54 avdd.t55 avdd.t13 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=8
X1899 dvss.t1789 dvdd.t1874 dvss.t1788 dvss.t1787 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1900 dvdd.t467 a_36756_35603# a_36743_35995# dvdd.t466 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X1901 dvdd.t71 a_35202_29877# por_dig_0.net30 dvdd.t70 sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.26 ps=2.52 w=1 l=0.15
X1902 dvss.t2106 por_dig_0.net20.t7 a_34378_35629# dvss.t1265 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X1903 por_ana_0.rstring_mux_0.vtrip_decoded_b_avdd[5] por_ana_0.rstring_mux_0.vtrip_decoded_avdd[5].t3 avdd.t504 avdd.t503 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X1904 dvdd.t907 por_dig_0._027_ a_34102_29645# dvdd.t70 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1905 a_37528_31527# por_dig_0.net34 dvdd.t868 dvdd.t867 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X1906 pwup_filt.t25 por_ana_0.sky130_fd_sc_hd__inv_4_0.Y dvdd.t213 dvdd.t212 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1907 a_21354_24707# a_21254_24619# dvss.t1083 dvss.t1082 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X1908 por_dig_0.cnt_por\[9\] a_35468_30163# dvdd.t450 dvdd.t449 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X1909 a_35000_31795# por_dig_0.net23.t17 dvdd.t765 dvdd.t764 sky130_fd_pr__pfet_01v8_hvt ad=0.2125 pd=1.425 as=0.305 ps=1.61 w=1 l=0.15
X1910 por_ana_0.comparator_0.vpp.t41 por_ana_0.comparator_0.vnn.t57 avdd.t372 avdd.t191 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1911 dvdd.t597 por_dig_0.clknet_1_1__leaf_osc_ck.t38 a_32740_35091# dvdd.t596 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1912 avss.t386 por_ana_0.rstring_mux_0.ena.t9 por_ana_0.rstring_mux_0.ena_b avss.t385 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X1913 vin.t4 avdd.t52 vin.t4 avdd.t53 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=0.6
X1914 dvdd.t1729 dvss.t2310 dvdd.t1728 dvdd.t1727 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X1915 a_37961_33287# a_36880_32915# a_37614_32883# dvdd.t431 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X1916 a_32812_30733# por_dig_0.net24 dvdd.t337 dvdd.t336 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X1917 dvdd.t1732 dvss.t2311 dvdd.t1731 dvdd.t1730 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X1918 dvss.t1369 a_27590_22885# a_27690_22973# dvss.t1368 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X1919 a_24968_13935# a_25346_6535# avss.t173 sky130_fd_pr__res_xhigh_po_1p41 l=35
X1920 dvss.t423 por_dig_0.net24 a_32966_31099# dvss.t422 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X1921 por_ana_0.sky130_fd_sc_hd__inv_4_1.A por_dig_0.por_unbuf.t16 dvss.t814 dvss.t813 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1922 a_32913_35629# por_dig_0._051_ a_32610_35603# dvss.t773 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.089375 ps=0.925 w=0.65 l=0.15
X1923 itest.t1 por_ana_0.ibias_gen_0.vp.t10 avdd.t385 avdd.t384 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X1924 a_7835_22912# a_8213_15512# avss.t27 sky130_fd_pr__res_xhigh_po_1p41 l=35
X1925 dvdd.t39 por_ana_0.sky130_fd_sc_hd__inv_4_3.Y dcomp.t17 dvdd.t38 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1926 a_25846_21903# a_25478_22885# dvdd.t1262 dvdd.t1261 sky130_fd_pr__pfet_01v8_hvt ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X1927 avdd.t283 a_29802_22973# a_30495_21859# avdd.t282 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.1365 ps=1.49 w=0.42 l=1
X1928 por_dig_0.clknet_0_osc_ck.t4 a_34387_32909# dvss.t143 dvss.t142 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1929 pwup_filt.t3 por_ana_0.sky130_fd_sc_hd__inv_4_0.Y dvss.t234 dvss.t233 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1930 por_dig_0.clknet_0_osc_ck.t3 a_34387_32909# dvss.t141 dvss.t140 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1931 a_25846_23637# a_25478_24619# dvdd.t1213 dvdd.t1212 sky130_fd_pr__pfet_01v8_hvt ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X1932 a_33482_31527# por_dig_0._036_.t6 por_dig_0._026_ dvdd.t1349 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.174 ps=1.39 w=1 l=0.15
X1933 por_ana_0.comparator_1.vt.t23 vin.t62 por_ana_0.comparator_1.vpp.t43 por_ana_0.comparator_1.vt.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1934 avdd.t387 por_ana_0.ibias_gen_0.vp.t11 itest.t0 avdd.t386 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X1935 por_ana_0.rstring_mux_0.vtrip1.t4 por_ana_0.rstring_mux_0.vtrip0.t0 avss.t214 sky130_fd_pr__res_xhigh_po_1p41 l=35
X1936 a_34719_23593# a_34294_23637# dvss.t1341 dvss.t1340 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X1937 por_timed_out.t2 a_31413_32339# dvdd.t722 dvdd.t721 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X1938 dvss.t816 por_dig_0.por_unbuf.t17 por_ana_0.sky130_fd_sc_hd__inv_4_1.A dvss.t815 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1939 dvdd.t962 por_ana_0.sky130_fd_sc_hd__inv_4_4.Y por.t23 dvdd.t961 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1940 por_ana_0.comparator_0.vpp.t27 vbg_1v2.t30 por_ana_0.comparator_0.vt.t42 por_ana_0.comparator_0.vt.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1941 dvss.t1033 a_35111_28013# a_35217_28013# dvss.t677 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X1942 a_37301_33453# por_dig_0._001_ dvss.t1088 dvss.t1087 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X1943 por_ana_0.comparator_0.ena_b.t0 avss.t431 avdd.t523 avdd.t522 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X1944 a_38123_32909# a_37046_32915# a_37961_33287# dvdd.t435 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X1945 por_ana_0.comparator_0.vn.t4 por_ana_0.comparator_0.vn.t3 avss.t389 avss.t45 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1946 dvdd.t790 a_34946_30431# a_34836_30555# dvdd.t789 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X1947 por_ana_0.comparator_0.vpp.t28 vbg_1v2.t31 por_ana_0.comparator_0.vt.t41 por_ana_0.comparator_0.vt.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1948 a_24159_23593# a_23734_23637# dvss.t1127 dvss.t1126 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X1949 por.t22 por_ana_0.sky130_fd_sc_hd__inv_4_4.Y dvdd.t960 dvdd.t959 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1950 a_34235_31277# por_dig_0.net22.t17 a_33940_31277# dvss.t1176 sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.143 ps=1.09 w=0.65 l=0.15
X1951 isrc_sel.t0 dvss.t1604 dvss.t1606 dvss.t1605 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X1952 dvss.t676 a_25578_24707# a_26785_24371# dvss.t675 sky130_fd_pr__nfet_g5v0d10v5 ad=0.121875 pd=1.075 as=0.19875 ps=2.03 w=0.75 l=0.5
X1953 por_ana_0.ibias_gen_0.vn0.t15 vbg_1v2.t32 por_ana_0.ibias_gen_0.vstart.t0 avss.t150 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X1954 por_dig_0.net15 por_dig_0.net5.t14 dvss.t2120 dvss.t2119 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1955 por_dig_0.net17 a_35130_28673# dvss.t723 dvss.t722 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.122275 ps=1.08 w=0.65 l=0.15
X1956 a_31802_32909# a_31566_32909# dvdd.t1199 dvdd.t1198 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.5
X1957 a_35802_32365# por_dig_0.net23.t18 dvss.t884 dvss.t883 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.13165 ps=1.14 w=0.42 l=0.15
X1958 por_ana_0.sky130_fd_sc_hvl__lsbuflv2hv_1_0[0|8].X a_39457_22637# dvss.t1041 dvss.t1040 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.121875 ps=1.075 w=0.75 l=0.5
X1959 dvss.t797 por_dig_0.net6 por_dig_0.net11 dvss.t796 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1960 a_32809_32365# a_31894_32365# a_32462_32607# dvss.t1971 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X1961 vin.t31 por_ana_0.rstring_mux_0.otrip_decoded_avdd[5] por_ana_0.rstring_mux_0.vtrip5.t5 avss.t260 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X1962 por_ana_0.rstring_mux_0.vtrip6.t1 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[6].t4 por_ana_0.comparator_0.vinn.t20 avss.t211 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X1963 a_32630_32915# a_32464_32915# dvdd.t402 dvdd.t401 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1964 por_ana_0.rstring_mux_0.vtop.t5 por_ana_0.rstring_mux_0.ena_b avdd.t229 avdd.t228 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X1965 a_25578_24707# a_25478_24619# dvss.t1480 dvss.t1479 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X1966 dvss.t689 a_36564_32339# por_dig_0.net23.t0 dvss.t688 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.0567 ps=0.69 w=0.42 l=0.15
X1967 a_32609_31099# por_dig_0._013_ dvdd.t1016 dvdd.t1015 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X1968 por_ana_0.comparator_1.n0.t4 por_ana_0.comparator_1.vm.t8 avss.t347 avss.t294 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1969 por_ana_0.ibias_gen_0.vp.t1 avss.t70 por_ana_0.ibias_gen_0.vp.t1 avss.t71 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=0.6
X1970 por_ana_0.rc_osc_0.n.t5 dvdd.t1287 por_ana_0.rc_osc_0.m dvdd.t1288 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X1971 a_36328_36493# por_dig_0._050_ dvss.t1010 dvss.t1009 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X1972 dvss.t670 a_30070_21903# a_30495_21859# dvss.t669 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X1973 a_33380_35879# por_dig_0._016_ dvdd.t1155 dvdd.t1154 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X1974 porb.t6 por_ana_0.sky130_fd_sc_hd__inv_4_1.Y dvss.t337 dvss.t336 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1975 a_34633_36147# por_dig_0.cnt_por\[1\] a_34856_36493# dvss.t1399 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1976 dvss.t1603 dvss.t1601 a_36038_24619# dvss.t1602 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X1977 a_34746_29965# por_dig_0.net29 dvss.t214 dvss.t213 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1978 a_31592_30965# a_31864_30823# a_31822_30849# dvdd.t1009 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X1979 a_31592_30965# a_31864_30823# dvss.t1198 dvss.t1197 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1980 avdd.t51 avdd.t49 avdd.t50 avdd.t3 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=8
X1981 dvdd.t159 a_34098_30707# por_dig_0.clknet_1_0__leaf_osc_ck.t21 dvdd.t158 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1982 a_31932_31419# por_dig_0.clknet_1_0__leaf_osc_ck.t43 dvdd.t422 dvdd.t396 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1983 a_34212_33997# por_dig_0.net22.t18 dvdd.t605 dvdd.t604 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1475 ps=1.295 w=1 l=0.15
X1984 a_37751_31251# por_dig_0._045_ dvdd.t1147 dvdd.t1146 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X1985 dvdd.t1342 a_31412_31251# por_dig_0.cnt_rsb_stg1 dvdd.t425 sky130_fd_pr__pfet_01v8_hvt ad=0.3012 pd=2.66 as=0.26 ps=2.52 w=1 l=0.15
X1986 dvss.t1786 dvdd.t1875 dvss.t1785 dvss.t1784 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X1987 dvdd.t958 por_ana_0.sky130_fd_sc_hd__inv_4_4.Y por.t21 dvdd.t957 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1988 dvss.t867 por_dig_0._034_.t14 por_dig_0.net19 dvss.t866 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1989 dvss.t550 por_dig_0._018_ a_35582_34317# dvss.t549 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X1990 a_38506_32365# por_dig_0.cnt_st\[0\] a_38434_32365# dvss.t1330 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X1991 dvdd.t1383 por_dig_0.net21 a_39732_31829# dvdd.t1382 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X1992 por_ana_0.rstring_mux_0.otrip_decoded_avdd[2] a_24673_22637# avdd.t650 avdd.t596 sky130_fd_pr__pfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.24375 ps=1.825 w=1.5 l=0.5
X1993 dvss.t1499 a_35960_29101# por_dig_0.otrip_decoded[6].t0 dvss.t1498 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X1994 dvss.t335 por_ana_0.sky130_fd_sc_hd__inv_4_1.Y porb.t5 dvss.t334 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1995 avdd.t373 por_ana_0.comparator_0.vnn.t58 por_ana_0.comparator_0.vpp.t42 avdd.t195 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1996 a_37886_31111# a_36696_30739# a_37777_31111# dvss.t1262 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1997 a_27958_21903# a_27590_22885# dvdd.t1139 dvdd.t1138 sky130_fd_pr__pfet_01v8_hvt ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X1998 dvss.t705 por_dig_0.clknet_1_1__leaf_osc_ck.t39 a_37064_34003# dvss.t704 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1999 por_ana_0.comparator_1.vpp.t9 por_ana_0.comparator_1.vpp.t8 avdd.t397 avdd.t395 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X2000 a_27958_23637# a_27590_24619# dvdd.t1141 dvdd.t1140 sky130_fd_pr__pfet_01v8_hvt ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X2001 a_37584_35389# a_37409_35463# a_37763_35451# dvss.t662 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X2002 a_30495_21859# a_30070_21903# dvss.t668 dvss.t667 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X2003 avdd.t488 por_ana_0.comparator_0.n1.t14 por_ana_0.dcomp3v3uv avdd.t487 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X2004 vin.t33 por_ana_0.rstring_mux_0.otrip_decoded_b_avdd[5] por_ana_0.rstring_mux_0.vtrip5.t7 avdd.t469 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X2005 por_dig_0.clknet_1_0__leaf_osc_ck.t20 a_34098_30707# dvdd.t157 dvdd.t156 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2006 por_dig_0.net24 a_35100_32339# dvdd.t1046 dvdd.t1045 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.3 ps=2.6 w=1 l=0.15
X2007 por_ana_0.rstring_mux_0.vtrip6.t3 por_ana_0.rstring_mux_0.vtrip_decoded_b_avdd[6] por_ana_0.comparator_0.vinn.t40 avdd.t558 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X2008 avdd.t48 avdd.t47 avdd.t48 avdd.t13 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=8
X2009 dvss.t1961 por_dig_0._039_ a_38986_34317# dvss.t1960 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2010 a_30495_21859# a_30070_21903# dvss.t666 dvss.t665 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X2011 dcomp.t6 por_ana_0.sky130_fd_sc_hd__inv_4_3.Y dvss.t61 dvss.t60 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2012 por_dig_0.net4 a_39417_31795# dvss.t546 dvss.t545 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X2013 dvss.t576 a_35583_34541# por_dig_0.clknet_1_1__leaf_osc_ck.t5 dvss.t575 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2014 dvss.t1045 por_dig_0._041_ a_39630_33229# dvss.t1044 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X2015 a_19676_13935# a_19298_6535# avss.t215 sky130_fd_pr__res_xhigh_po_1p41 l=35
X2016 a_26271_23593# a_25846_23637# dvss.t364 dvss.t363 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X2017 a_31984_31821# a_31360_31827# a_31876_32199# dvdd.t20 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X2018 a_33172_28165# por_dig_0.net5.t15 dvdd.t1448 dvdd.t1447 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14575 ps=1.335 w=0.42 l=0.15
X2019 dvss.t1783 dvdd.t1876 dvss.t1782 dvss.t1781 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X2020 a_22700_13935# a_22322_6535# avss.t216 sky130_fd_pr__res_xhigh_po_1p41 l=35
X2021 dvdd.t1055 a_37392_31251# por_dig_0._004_ dvdd.t1054 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2022 porb.t4 por_ana_0.sky130_fd_sc_hd__inv_4_1.Y dvss.t333 dvss.t332 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2023 por_ana_0.rstring_mux_0.vtrip0.t1 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[0] por_ana_0.comparator_0.vinn.t22 avss.t221 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X2024 dvss.t1780 dvdd.t1877 dvss.t1779 dvss.t1723 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X2025 por_ana_0.schmitt_trigger_0.in.t10 dvss.t657 sky130_fd_pr__cap_mim_m3_2 l=30 w=30
X2026 a_33172_28165# por_dig_0.net5.t16 dvss.t2122 dvss.t2121 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.10025 ps=0.985 w=0.42 l=0.15
X2027 dvss.t1778 dvdd.t1878 dvss.t1777 dvss.t1776 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X2028 por_ana_0.rstring_mux_0.otrip_decoded_b_avdd[3] por_ana_0.rstring_mux_0.otrip_decoded_avdd[3] avdd.t450 avdd.t449 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X2029 dvdd.t335 por_dig_0.net24 a_31412_33427# dvdd.t334 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X2030 a_38146_31429# a_38242_31251# dvdd.t1100 dvdd.t1099 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14075 ps=1.325 w=0.42 l=0.5
X2031 dvdd.t607 por_dig_0.net22.t19 por_dig_0._020_ dvdd.t606 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2032 avdd.t213 a_26271_23593# a_25578_24707# avdd.t212 sky130_fd_pr__pfet_g5v0d10v5 ad=0.2142 pd=1.99 as=0.2142 ps=1.99 w=0.42 l=1
X2033 dvss.t192 a_34098_30707# por_dig_0.clknet_1_0__leaf_osc_ck.t6 dvss.t191 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2034 avdd.t374 por_ana_0.comparator_0.vnn.t59 por_ana_0.comparator_0.vpp.t43 avdd.t195 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X2035 dvss.t190 a_34098_30707# por_dig_0.clknet_1_0__leaf_osc_ck.t5 dvss.t189 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2036 por_ana_0.ibias_gen_0.vp0.t2 por_ana_0.ibias_gen_0.vp0.t1 avdd.t549 avdd.t548 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X2037 a_27690_24707# a_27590_24619# dvss.t1383 dvss.t1382 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X2038 a_38145_34375# a_37064_34003# a_37798_33971# dvdd.t1073 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X2039 a_32354_30739# a_32188_30739# dvdd.t816 dvdd.t815 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2040 avss.t191 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.t27 porb_h.t25 avss.t190 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X2041 a_39738_32909# por_dig_0._041_ por_dig_0._002_ dvdd.t904 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.174 ps=1.39 w=1 l=0.15
X2042 dvdd.t143 por_dig_0._031_ a_38936_32159# dvdd.t142 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X2043 a_35704_35451# a_35450_35124# dvss.t727 dvss.t726 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1449 ps=1.11 w=0.42 l=0.15
X2044 a_13628_13935# a_14006_6535# avss.t217 sky130_fd_pr__res_xhigh_po_1p41 l=35
X2045 dvdd.t113 a_34387_32909# por_dig_0.clknet_0_osc_ck.t21 dvdd.t112 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2046 dvss.t1116 a_32182_21903# a_32607_21859# dvss.t1115 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X2047 por_dig_0.cnt_st\[1\] a_38136_33427# dvdd.t233 dvdd.t232 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X2048 a_27690_24707# a_27590_24619# dvss.t1381 dvss.t1380 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X2049 por_dig_0.otrip_decoded[0].t3 a_38444_28013# dvdd.t1316 dvdd.t1315 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X2050 avdd.t420 a_29802_24707# a_31009_24371# avdd.t419 sky130_fd_pr__pfet_g5v0d10v5 ad=0.24375 pd=1.825 as=0.3975 ps=3.53 w=1.5 l=0.5
X2051 dvdd.t1735 dvss.t2312 dvdd.t1734 dvdd.t1733 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X2052 a_35776_36967# por_dig_0.cnt_por\[0\].t18 dvdd.t539 dvdd.t538 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1475 ps=1.295 w=1 l=0.15
X2053 por_dig_0.clknet_1_1__leaf_osc_ck.t4 a_35583_34541# dvss.t574 dvss.t573 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2054 a_39248_32365# por_dig_0.cnt_st\[3\] a_39152_32365# dvss.t931 sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0693 ps=0.75 w=0.42 l=0.15
X2055 dvss.t785 a_27958_23637# a_28383_23593# dvss.t784 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X2056 dvdd.t187 por_ana_0.sky130_fd_sc_hd__inv_4_1.A por_ana_0.sky130_fd_sc_hd__inv_4_1.Y dvdd.t186 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2057 por_dig_0._050_ a_35592_36286# dvss.t1008 dvss.t1007 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X2058 dvss.t1575 por_dig_0.cnt_por\[2\] a_34948_35451# dvss.t1574 sky130_fd_pr__nfet_01v8 ad=0.196275 pd=1.33 as=0.0693 ps=0.75 w=0.42 l=0.15
X2059 por_dig_0._047_ a_33600_34335# dvss.t450 dvss.t449 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X2060 a_15140_13935# a_14762_6535# avss.t218 sky130_fd_pr__res_xhigh_po_1p41 l=35
X2061 dvdd.t79 por_dig_0.net4 a_33482_31527# dvdd.t78 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X2062 avss.t404 por_ana_0.ibias_gen_0.vn1.t14 por_ana_0.ibias_gen_0.vp1.t5 avss.t396 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=8
X2063 dvss.t1067 a_21254_22885# a_21354_22973# dvss.t1066 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X2064 por_ana_0.sky130_fd_sc_hd__inv_4_3.Y por_ana_0.vl dvdd.t996 dvdd.t995 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2065 por_ana_0.comparator_0.vnn.t14 avss.t432 avdd.t525 avdd.t524 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X2066 avdd.t209 a_36138_22973# a_36831_21859# avdd.t208 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.1365 ps=1.49 w=0.42 l=1
X2067 dvss.t218 por_dig_0.otrip_decoded[1] a_21254_24619# dvss.t217 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X2068 dvss.t1775 dvdd.t1879 dvss.t1774 dvss.t1773 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X2069 a_35913_33819# a_35699_33819# dvdd.t1153 dvdd.t1152 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07035 ps=0.755 w=0.42 l=0.15
X2070 a_36305_31277# a_35224_31277# a_35958_31519# dvdd.t1089 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X2071 dvdd.t1737 dvss.t2313 dvdd.t1736 dvdd.t1556 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X2072 avdd.t46 avdd.t43 avdd.t45 avdd.t44 sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.58 as=0 ps=0 w=5 l=4
X2073 por_ana_0.comparator_1.vt.t7 avss.t433 por_ana_0.comparator_1.vnn.t32 por_ana_0.comparator_1.vt.t3 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=8
X2074 por_ana_0.rstring_mux_0.vtrip0.t3 por_ana_0.rstring_mux_0.vtrip_decoded_b_avdd[0] por_ana_0.comparator_0.vinn.t24 avdd.t425 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X2075 dvdd.t792 a_38145_34375# a_38320_34301# dvdd.t791 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X2076 avdd.t375 por_ana_0.comparator_0.vnn.t60 por_ana_0.comparator_0.vpp.t44 avdd.t195 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X2077 dvdd.t1739 dvss.t2314 dvdd.t1738 dvdd.t1534 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X2078 dvss.t2082 por_dig_0.cnt_por\[5\] a_34357_33427# dvss.t2081 sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.10725 ps=0.98 w=0.65 l=0.15
X2079 porb_h.t2 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.t28 avdd.t349 avdd.t348 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X2080 dvdd.t994 por_ana_0.vl por_ana_0.sky130_fd_sc_hd__inv_4_3.Y dvdd.t993 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2081 a_34719_21859# a_34294_21903# dvss.t1491 dvss.t1490 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X2082 a_34948_35451# por_dig_0.cnt_por\[3\] a_34842_35451# dvss.t451 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X2083 por_ana_0.sky130_fd_sc_hd__inv_4_0.Y por_ana_0.schmitt_trigger_0.out.t11 dvss.t822 dvss.t821 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2084 a_36567_32141# por_dig_0._037_ dvss.t121 dvss.t120 sky130_fd_pr__nfet_01v8 ad=0.118625 pd=1.015 as=0.1365 ps=1.07 w=0.65 l=0.15
X2085 pwup_filt.t2 por_ana_0.sky130_fd_sc_hd__inv_4_0.Y dvss.t232 dvss.t231 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2086 por_ana_0.rc_osc_0.m por_ana_0.rc_osc_0.in dvdd.t237 dvdd.t236 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X2087 dvss.t1379 a_27590_24619# a_27690_24707# dvss.t1378 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X2088 dvdd.t990 otrip[0].t3 a_32039_28013# dvdd.t989 sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X2089 porb_h.t24 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.t29 avss.t193 avss.t192 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X2090 a_35874_32365# por_dig_0._033_ a_35802_32365# dvss.t34 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X2091 a_32651_33819# a_31932_33595# a_32088_33690# dvss.t2090 sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0594 ps=0.69 w=0.36 l=0.15
X2092 dvss.t1256 a_38956_32339# por_dig_0._031_ dvss.t1255 sky130_fd_pr__nfet_01v8 ad=0.196275 pd=1.33 as=0.169 ps=1.82 w=0.65 l=0.15
X2093 dvdd.t1286 dvdd.t1284 osc_ck.t2 dvdd.t1285 sky130_fd_pr__pfet_01v8 ad=0.1475 pd=1.295 as=0.15 ps=1.3 w=1 l=0.18
X2094 dvss.t131 a_39887_21959# a_40246_21893# dvss.t130 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.105 ps=1.03 w=0.75 l=0.5
X2095 dvdd.t1184 a_32922_30707# a_32812_30733# dvdd.t1183 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X2096 por_dig_0.clknet_1_1__leaf_osc_ck.t18 a_35583_34541# dvdd.t475 dvdd.t474 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2097 por_ana_0.schmitt_trigger_0.m.t3 por_ana_0.schmitt_trigger_0.in.t11 dvdd.t567 dvdd.t566 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X2098 a_33198_32883# a_32980_33287# dvdd.t527 dvdd.t526 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X2099 a_28383_23593# a_27958_23637# dvss.t783 dvss.t782 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X2100 dvss.t949 por_dig_0.net25 a_34990_30189# dvss.t948 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X2101 por_ana_0.comparator_0.vnn avss.t434 por_ana_0.comparator_0.vt.t25 por_ana_0.comparator_0.vt.t18 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=8
X2102 por_ana_0.rc_osc_0.vr dvdd.t1282 por_ana_0.rc_osc_0.ena_b dvdd.t1283 sky130_fd_pr__pfet_01v8 ad=0.1475 pd=1.295 as=0.145 ps=1.29 w=1 l=0.5
X2103 a_21622_23637# a_21254_24619# dvss.t1081 dvss.t1080 sky130_fd_pr__nfet_01v8 ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X2104 dvss.t230 por_ana_0.sky130_fd_sc_hd__inv_4_0.Y pwup_filt.t1 dvss.t229 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2105 dvdd.t29 por_dig_0._033_ a_34486_33703# dvdd.t28 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X2106 dvdd.t1412 a_36305_31277# a_36480_31251# dvdd.t1411 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X2107 a_31932_31419# por_dig_0.clknet_1_0__leaf_osc_ck.t44 dvss.t505 dvss.t504 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2108 dvss.t818 por_dig_0.por_unbuf.t18 a_25495_33620# dvss.t817 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X2109 por_ana_0.rstring_mux_0.vtrip5.t8 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[5].t4 por_ana_0.comparator_0.vinn.t36 avss.t302 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X2110 a_35958_31519# a_35740_31277# dvss.t1290 dvss.t1289 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X2111 por_ana_0.comparator_1.vpp.t7 por_ana_0.comparator_1.vpp.t6 avdd.t396 avdd.t395 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X2112 a_37301_33453# por_dig_0._001_ dvdd.t924 dvdd.t923 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X2113 a_21354_22973# a_21254_22885# dvss.t1065 dvss.t1064 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X2114 dvss.t1238 a_32984_32339# a_32918_32365# dvss.t1237 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X2115 a_37393_30189# por_dig_0._003_ dvdd.t663 dvdd.t662 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X2116 a_34302_34541# por_dig_0.cnt_por\[1\] por_dig_0._051_ dvss.t1398 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.195 ps=1.9 w=0.65 l=0.15
X2117 a_33934_32615# por_dig_0.cnt_por\[6\] dvdd.t388 dvdd.t387 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X2118 por.t20 por_ana_0.sky130_fd_sc_hd__inv_4_4.Y dvdd.t956 dvdd.t955 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2119 dvss.t298 a_38250_22973# a_39457_22637# dvss.t297 sky130_fd_pr__nfet_g5v0d10v5 ad=0.121875 pd=1.075 as=0.19875 ps=2.03 w=0.75 l=0.5
X2120 a_37777_31111# a_36862_30739# a_37430_30707# dvss.t1275 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X2121 avdd.t321 a_28383_23593# a_27690_24707# avdd.t320 sky130_fd_pr__pfet_g5v0d10v5 ad=0.2142 pd=1.99 as=0.2142 ps=1.99 w=0.42 l=1
X2122 por_ana_0.comparator_0.vnn avss.t435 por_ana_0.comparator_0.vt.t24 por_ana_0.comparator_0.vt.t18 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=8
X2123 a_33162_35603# por_dig_0._047_ dvss.t841 dvss.t840 sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.25675 ps=1.44 w=0.65 l=0.15
X2124 avss.t69 avss.t67 avss.t69 avss.t68 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=8
X2125 dvdd.t1742 dvss.t2315 dvdd.t1741 dvdd.t1740 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X2126 a_36410_36173# por_dig_0._049_ dvdd.t1014 dvdd.t1013 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X2127 dvss.t1772 dvdd.t1880 dvss.t1771 dvss.t1770 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X2128 por_ana_0.comparator_0.vm.t6 por_ana_0.comparator_0.ena_b.t3 avss.t333 avss.t100 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X2129 por_ana_0.comparator_1.vnn avss.t436 por_ana_0.comparator_1.vt.t6 por_ana_0.comparator_1.vt.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=8
X2130 dvss.t2031 por_dig_0.cnt_st\[2\] a_38506_32365# dvss.t2030 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X2131 a_36886_32141# por_dig_0._031_ a_36567_32141# dvss.t170 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.118625 ps=1.015 w=0.65 l=0.15
X2132 a_19094_870# a_41694_1248# dvss.t895 sky130_fd_pr__res_xhigh_po_1p41 l=111
X2133 dvss.t1489 a_34294_21903# a_34719_21859# dvss.t1488 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X2134 a_32828_35879# por_dig_0._047_ a_32610_35603# dvdd.t725 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.26 ps=2.52 w=1 l=0.15
X2135 dvdd.t954 por_ana_0.sky130_fd_sc_hd__inv_4_4.Y por.t19 dvdd.t953 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2136 avdd.t587 a_31914_24707# a_33121_24371# avdd.t556 sky130_fd_pr__pfet_g5v0d10v5 ad=0.24375 pd=1.825 as=0.3975 ps=3.53 w=1.5 l=0.5
X2137 a_33821_36551# a_32740_36179# a_33474_36147# dvdd.t375 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X2138 dvss.t706 por_dig_0.clknet_1_1__leaf_osc_ck.t40 a_36880_33453# dvss.t702 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2139 a_35632_35124# a_35450_35124# dvdd.t621 dvdd.t620 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X2140 dvdd.t609 por_dig_0.net22.t20 a_33934_32615# dvdd.t608 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X2141 dvss.t777 a_34828_29253# por_dig_0.net15 dvss.t776 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.221 ps=1.98 w=0.65 l=0.15
X2142 por_ana_0.comparator_1.vt.t22 vin.t63 por_ana_0.comparator_1.vpp.t44 por_ana_0.comparator_1.vt.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X2143 a_39888_23693# a_39888_24823# avdd.t312 avdd.t311 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.1197 ps=1.41 w=0.42 l=0.5
X2144 dvdd.t1344 por_dig_0.cnt_rsb_stg1 a_31566_32909# dvdd.t1343 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2145 por_dig_0.net11 por_dig_0.net7.t17 dvss.t860 dvss.t859 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2146 a_40246_21893# a_39887_21959# dvss.t129 dvss.t128 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.178875 ps=1.26 w=0.75 l=0.5
X2147 dvss.t910 a_23366_22885# a_23466_22973# dvss.t909 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X2148 dvss.t1258 a_40247_23627# por_ana_0.vl dvss.t1257 sky130_fd_pr__nfet_01v8 ad=0.1961 pd=2.01 as=0.1961 ps=2.01 w=0.74 l=0.15
X2149 dvss.t2231 a_31413_29075# por_dig_0.force_pdnb dvss.t2230 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X2150 avss.t15 por_ana_0.comparator_1.n1.t14 por_ana_0.dcomp3v3 avss.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.6
X2151 dvdd.t424 por_dig_0.clknet_1_0__leaf_osc_ck.t45 a_32464_32915# dvdd.t423 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X2152 dvss.t1242 a_35100_32339# por_dig_0.net24 dvss.t1241 sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.0588 ps=0.7 w=0.42 l=0.15
X2153 por_ana_0.schmitt_trigger_0.m.t11 por_ana_0.schmitt_trigger_0.out.t12 dvdd.t714 dvdd.t713 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X2154 avdd.t251 a_38250_22973# a_38943_21859# avdd.t250 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.1365 ps=1.49 w=0.42 l=1
X2155 dvss.t1302 por_dig_0.otrip_decoded[3].t5 a_23366_24619# dvss.t1301 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X2156 por_ana_0.comparator_1.vt.t21 vin.t64 por_ana_0.comparator_1.vpp.t45 por_ana_0.comparator_1.vt.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X2157 dvss.t1769 dvdd.t1881 dvss.t1768 dvss.t1682 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X2158 a_33242_28263# a_33172_28165# por_dig_0.net12 dvdd.t944 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.32 ps=2.64 w=1 l=0.15
X2159 por_dig_0.cnt_por\[8\] a_33444_31037# dvss.t380 dvss.t379 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X2160 por_ana_0.rstring_mux_0.vtrip5.t3 por_ana_0.rstring_mux_0.vtrip_decoded_b_avdd[5] por_ana_0.comparator_0.vinn.t29 avdd.t459 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X2161 a_35612_33595# por_dig_0.clknet_1_1__leaf_osc_ck.t41 dvdd.t599 dvdd.t598 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2162 dvdd.t27 por_dig_0._033_ a_36414_32909# dvdd.t26 sky130_fd_pr__pfet_01v8_hvt ad=0.1475 pd=1.295 as=0.14 ps=1.28 w=1 l=0.15
X2163 avdd.t42 avdd.t41 avdd.t42 avdd.t13 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=8
X2164 a_34836_30555# a_34212_30189# a_34728_30189# dvdd.t1081 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X2165 dvdd.t541 por_dig_0.cnt_por\[0\].t19 por_dig_0._034_.t2 dvdd.t540 sky130_fd_pr__pfet_01v8_hvt ad=0.335 pd=1.67 as=0.135 ps=1.27 w=1 l=0.15
X2166 por_dig_0._051_ por_dig_0.cnt_por\[2\] dvdd.t1270 dvdd.t1269 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2167 a_35925_35451# por_dig_0._046_ a_35704_35124# dvss.t2152 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X2168 por_ana_0.rstring_mux_0.vtop.t4 por_ana_0.rstring_mux_0.ena_b avdd.t227 avdd.t226 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X2169 dvss.t1767 dvdd.t1882 dvss.t1766 dvss.t1765 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X2170 a_32966_31099# a_32922_30707# a_32800_31111# dvss.t1428 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X2171 avss.t66 avss.t63 avss.t65 avss.t64 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=8
X2172 a_35674_28557# por_dig_0.net7.t18 dvdd.t747 dvdd.t746 sky130_fd_pr__pfet_01v8_hvt ad=0.1087 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X2173 dvss.t1036 a_40246_21893# por_ana_0.sky130_fd_sc_hvl__lsbufhv2lv_1_1.X dvss.t1035 sky130_fd_pr__nfet_01v8 ad=0.1961 pd=2.01 as=0.1961 ps=2.01 w=0.74 l=0.15
X2174 a_33806_33427# por_dig_0._047_ dvss.t839 dvss.t838 sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.25675 ps=1.44 w=0.65 l=0.15
X2175 por_ana_0.rstring_mux_0.otrip_decoded_b_avdd[2] por_ana_0.rstring_mux_0.otrip_decoded_avdd[2] avdd.t1 avdd.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X2176 vin.t38 dvss.t1598 dvss.t1600 dvss.t1599 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X2177 a_34796_13935# a_35174_6535# avss.t154 sky130_fd_pr__res_xhigh_po_1p41 l=35
X2178 dvss.t1764 dvdd.t1883 dvss.t1763 dvss.t1688 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X2179 por_dig_0.clknet_1_0__leaf_osc_ck.t4 a_34098_30707# dvss.t188 dvss.t187 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2180 dvss.t1762 dvdd.t1884 dvss.t1761 dvss.t1760 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X2181 a_38136_33213# a_37961_33287# a_38315_33275# dvss.t621 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X2182 a_23466_22973# a_23366_22885# dvss.t908 dvss.t907 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X2183 porb_h.t23 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.t30 avss.t195 avss.t194 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X2184 a_37485_34363# por_dig_0._000_ dvss.t897 dvss.t896 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X2185 osc_ck.t5 por_ana_0.rc_osc_0.n.t10 dvss.t2022 dvss.t2021 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X2186 por_dig_0.cnt_por\[0\].t6 a_36756_35603# dvdd.t465 dvdd.t464 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2187 a_33899_33275# por_dig_0.net24 dvss.t421 dvss.t420 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X2188 por_dig_0.net6 a_33971_28557# dvdd.t1143 dvdd.t1142 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X2189 dvdd.t897 a_33474_36147# a_33364_36173# dvdd.t896 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X2190 por_ana_0.dcomp3v3uv por_ana_0.comparator_0.n1.t15 avdd.t490 avdd.t489 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X2191 por_dig_0._029_ por_dig_0.cnt_st\[1\] dvdd.t503 dvdd.t502 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2192 dvss.t1310 a_36406_21903# a_36831_21859# dvss.t1309 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X2193 a_36476_30163# por_dig_0.cnt_por\[10\] dvss.t1510 dvss.t1509 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2194 por_ana_0.ibias_gen_0.vp1.t4 por_ana_0.ibias_gen_0.vn1.t15 avss.t405 avss.t398 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=8
X2195 avdd.t287 a_34026_24707# a_35233_24371# avdd.t286 sky130_fd_pr__pfet_g5v0d10v5 ad=0.24375 pd=1.825 as=0.3975 ps=3.53 w=1.5 l=0.5
X2196 a_39162_33453# a_38926_33453# dvss.t729 dvss.t728 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.5
X2197 a_32149_32365# por_dig_0._012_ dvdd.t1190 dvdd.t1189 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X2198 dvdd.t235 por_ana_0.rc_osc_0.in por_ana_0.rc_osc_0.m dvdd.t234 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X2199 dvss.t1024 por_dig_0.force_pdnb a_38150_22885# dvss.t1023 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X2200 dvss.t186 a_34098_30707# por_dig_0.clknet_1_0__leaf_osc_ck.t3 dvss.t185 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2201 a_33821_36551# a_32906_36179# a_33474_36147# dvss.t720 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X2202 a_31412_33427# a_31615_33705# dvdd.t720 dvdd.t719 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1134 ps=1.38 w=0.42 l=0.15
X2203 por_dig_0._020_ por_dig_0._019_ dvdd.t1488 dvdd.t1487 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2204 dvss.t2176 por_dig_0._019_ a_34734_34363# dvss.t2175 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X2205 dvss.t1560 a_25478_22885# a_25578_22973# dvss.t1559 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X2206 a_36952_35085# a_36328_35091# a_36844_35463# dvdd.t871 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X2207 a_37301_33275# por_dig_0._002_ dvdd.t1300 dvdd.t1299 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X2208 por_ana_0.comparator_1.vn.t0 por_ana_0.rstring_mux_0.ena.t10 por_ana_0.ibias_gen_0.ibias0.t3 avss.t387 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X2209 por_dig_0.clknet_1_1__leaf_osc_ck.t17 a_35583_34541# dvdd.t473 dvdd.t472 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2210 dvss.t1759 dvdd.t1885 dvss.t1758 dvss.t1757 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X2211 avss.t197 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.t31 porb_h.t22 avss.t196 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X2212 a_35640_32517# por_dig_0.cnt_por\[4\] a_35874_32365# dvss.t1547 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X2213 dvdd.t1744 dvss.t2316 dvdd.t1743 dvdd.t1578 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X2214 a_34114_35879# por_dig_0.cnt_por\[3\] a_33896_35603# dvdd.t380 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2215 dvdd.t305 a_37614_33695# a_37504_33819# dvdd.t304 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X2216 dvss.t1339 a_39718_33605# por_dig_0._040_ dvss.t1338 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.169 ps=1.82 w=0.65 l=0.15
X2217 dvdd.t426 por_dig_0.clknet_1_0__leaf_osc_ck.t46 a_31360_31827# dvdd.t425 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X2218 dvdd.t786 a_37706_30431# a_37596_30555# dvdd.t785 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X2219 a_3299_22912# a_3677_15512# avss.t27 sky130_fd_pr__res_xhigh_po_1p41 l=35
X2220 avdd.t513 a_23466_24707# a_24159_23593# avdd.t512 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.1365 ps=1.49 w=0.42 l=1
X2221 dvss.t1079 a_21254_24619# a_21354_24707# dvss.t1078 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X2222 a_35111_28013# a_34934_28013# dvss.t1032 dvss.t523 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X2223 dvss.t1756 dvdd.t1886 dvss.t1755 dvss.t1754 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X2224 dvss.t1753 dvdd.t1887 dvss.t1752 dvss.t1703 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X2225 a_35774_28673# por_dig_0.net6 dvdd.t672 dvdd.t671 sky130_fd_pr__pfet_01v8_hvt ad=0.074375 pd=0.815 as=0.0567 ps=0.69 w=0.42 l=0.15
X2226 dvss.t795 por_dig_0.net6 por_dig_0.net15 dvss.t794 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.08775 ps=0.92 w=0.65 l=0.15
X2227 a_39813_31277# por_dig_0._042_ a_39510_31251# dvss.t304 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.089375 ps=0.925 w=0.65 l=0.15
X2228 por_dig_0._023_ a_34580_34110# dvss.t1218 dvss.t1217 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X2229 por_ana_0.rstring_mux_0.vtrip3.t6 por_ana_0.rstring_mux_0.otrip_decoded_avdd[3] vin.t27 avss.t238 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X2230 dvss.t1329 por_dig_0.cnt_st\[0\] a_39718_33605# dvss.t1328 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2231 a_38228_30163# a_38053_30189# a_38407_30189# dvss.t117 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X2232 por_dig_0._006_ por_dig_0._050_ a_36410_36173# dvdd.t877 sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.39 as=0.105 ps=1.21 w=1 l=0.15
X2233 a_33161_35451# por_dig_0._008_ dvdd.t324 dvdd.t323 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X2234 por_ana_0.comparator_0.vnn.t28 por_ana_0.comparator_0.vinn.t58 por_ana_0.comparator_0.vt.t7 por_ana_0.comparator_0.vt.t3 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X2235 a_38320_34301# por_dig_0.net25 dvdd.t833 dvdd.t832 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X2236 a_33934_29645# por_dig_0._027_ a_33852_29645# dvdd.t70 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2237 a_36382_31795# por_dig_0.cnt_st\[4\] a_36886_32141# dvss.t1527 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.06825 ps=0.86 w=0.65 l=0.15
X2238 a_39579_30849# por_dig_0.net4 a_39497_30849# dvdd.t77 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X2239 dvdd.t1747 dvss.t2317 dvdd.t1746 dvdd.t1745 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X2240 dvss.t824 por_ana_0.schmitt_trigger_0.out.t13 por_ana_0.sky130_fd_sc_hd__inv_4_0.Y dvss.t823 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2241 dvdd.t569 por_ana_0.schmitt_trigger_0.in.t12 por_ana_0.schmitt_trigger_0.m.t2 dvdd.t568 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X2242 force_ena_rc_osc.t0 dvss.t1595 dvss.t1597 dvss.t1596 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X2243 dvss.t1751 dvdd.t1888 dvss.t1750 dvss.t1749 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X2244 a_34444_32517# por_dig_0._026_ a_34842_32365# dvss.t1994 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.06825 ps=0.86 w=0.65 l=0.15
X2245 por_ana_0.comparator_0.vt.t39 vbg_1v2.t33 por_ana_0.comparator_0.vpp.t29 por_ana_0.comparator_0.vt.t36 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X2246 por_ana_0.schmitt_trigger_0.in.t13 dvss.t658 sky130_fd_pr__cap_mim_m3_2 l=30 w=30
X2247 dvdd.t1749 dvss.t2318 dvdd.t1748 dvdd.t1646 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X2248 a_5567_22912# a_5945_15512# avss.t27 sky130_fd_pr__res_xhigh_po_1p41 l=35
X2249 a_39417_31795# force_short_oneshot.t3 dvss.t847 dvss.t846 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X2250 por_ana_0.ibias_gen_0.vp0.t11 por_ana_0.rstring_mux_0.ena.t11 avdd.t614 avdd.t613 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X2251 dvss.t1463 a_25495_33620# a_25595_33708# dvss.t1462 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X2252 dvss.t88 por_dig_0.net4 a_33940_31277# dvss.t87 sky130_fd_pr__nfet_01v8 ad=0.105625 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X2253 por_dig_0.cnt_st\[4\] a_37952_31037# dvss.t1453 dvss.t1452 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X2254 a_32233_31643# a_32019_31643# dvdd.t1088 dvdd.t1087 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07035 ps=0.755 w=0.42 l=0.15
X2255 dvss.t262 a_38518_21903# a_38943_21859# dvss.t261 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X2256 a_32795_32187# por_dig_0.net8 dvss.t1419 dvss.t1418 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X2257 a_21354_24707# a_21254_24619# dvss.t1077 dvss.t1076 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X2258 a_36480_31251# por_dig_0.net25 dvdd.t831 dvdd.t830 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X2259 por_ana_0.comparator_1.vt.t5 avss.t437 por_ana_0.comparator_1.vnn.t31 por_ana_0.comparator_1.vt.t3 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=8
X2260 a_33930_35463# a_32740_35091# a_33821_35463# dvss.t1221 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X2261 dvdd.t1469 a_36100_32517# por_dig_0._019_ dvdd.t1468 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.26 ps=2.52 w=1 l=0.15
X2262 avdd.t306 a_36138_24707# a_37345_24371# avdd.t292 sky130_fd_pr__pfet_g5v0d10v5 ad=0.24375 pd=1.825 as=0.3975 ps=3.53 w=1.5 l=0.5
X2263 dvdd.t513 a_33162_35603# por_dig_0._008_ dvdd.t512 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2264 a_30070_21903# a_29702_22885# dvdd.t411 dvdd.t410 sky130_fd_pr__pfet_01v8_hvt ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X2265 dvdd.t601 por_dig_0.clknet_1_1__leaf_osc_ck.t42 a_36328_35091# dvdd.t600 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X2266 por_ana_0.comparator_0.vinn.t13 avss.t61 por_ana_0.comparator_0.vinn.t13 avss.t62 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=0.6
X2267 dvdd.t1752 dvss.t2319 dvdd.t1751 dvdd.t1750 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X2268 por_ana_0.rstring_mux_0.vtrip3.t8 por_ana_0.rstring_mux_0.otrip_decoded_b_avdd[3] vin.t29 avdd.t452 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X2269 avdd.t566 a_27690_22973# a_28897_22637# avdd.t565 sky130_fd_pr__pfet_g5v0d10v5 ad=0.24375 pd=1.825 as=0.3975 ps=3.53 w=1.5 l=0.5
X2270 a_30070_23637# a_29702_24619# dvdd.t1251 dvdd.t1250 sky130_fd_pr__pfet_01v8_hvt ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X2271 dvss.t793 por_dig_0.net6 a_36649_28789# dvss.t792 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.10785 ps=1.36 w=0.42 l=0.15
X2272 por_ana_0.comparator_1.vt.t4 avss.t438 por_ana_0.comparator_1.vnn.t30 por_ana_0.comparator_1.vt.t3 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=8
X2273 dvss.t708 por_dig_0.clknet_1_1__leaf_osc_ck.t43 a_32740_36179# dvss.t707 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2274 por_ana_0.ibias_gen_0.vp.t3 por_ana_0.ibias_gen_0.isrc_sel_b.t7 por_ana_0.ibias_gen_0.vp0.t8 avss.t337 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X2275 dvss.t1748 dvdd.t1889 dvss.t1747 dvss.t1746 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X2276 dvss.t631 por_dig_0.net26 a_32651_31643# dvss.t630 sky130_fd_pr__nfet_01v8 ad=0.2205 pd=1.89 as=0.066 ps=0.745 w=0.42 l=0.15
X2277 avdd.t616 por_ana_0.rstring_mux_0.ena.t12 por_ana_0.rstring_mux_0.ena_b avdd.t615 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X2278 por_ana_0.rstring_mux_0.otrip_decoded_b_avdd[4] por_ana_0.rstring_mux_0.otrip_decoded_avdd[4] avss.t377 avss.t376 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X2279 dvss.t468 a_32616_32125# a_32550_32199# dvss.t467 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X2280 dvss.t2079 a_31413_29619# por_dig_0.osc_ena.t1 dvss.t2078 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X2281 a_32971_32731# a_31894_32365# a_32809_32365# dvdd.t1311 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X2282 por_dig_0._041_ por_dig_0.net33 dvss.t1043 dvss.t1042 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X2283 dvss.t2011 a_31412_33427# por_dig_0.cnt_por\[6\] dvss.t2010 sky130_fd_pr__nfet_01v8 ad=0.2087 pd=2.02 as=0.169 ps=1.82 w=0.65 l=0.15
X2284 avdd.t301 a_25578_24707# a_26271_23593# avdd.t300 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.1365 ps=1.49 w=0.42 l=1
X2285 dvss.t1520 a_23366_24619# a_23466_24707# dvss.t1519 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X2286 por_dig_0.otrip_decoded[3].t2 a_37800_28013# dvdd.t1216 dvdd.t1215 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X2287 dvss.t1240 a_35100_32339# por_dig_0.net24 dvss.t1239 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2288 por_ana_0.rc_osc_0.in dvss.t288 sky130_fd_pr__cap_mim_m3_2 l=30 w=30
X2289 a_33804_31251# por_dig_0._036_.t7 a_34022_31527# dvdd.t1350 sky130_fd_pr__pfet_01v8_hvt ad=0.22 pd=1.44 as=0.1625 ps=1.325 w=1 l=0.15
X2290 a_35394_28013# a_35217_28013# dvdd.t438 dvdd.t437 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X2291 dvss.t894 a_29802_24707# a_31009_24371# dvss.t517 sky130_fd_pr__nfet_g5v0d10v5 ad=0.121875 pd=1.075 as=0.19875 ps=2.03 w=0.75 l=0.5
X2292 por_ana_0.dcomp3v3 por_ana_0.comparator_1.n1.t15 avss.t13 avss.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X2293 a_35848_31643# por_dig_0.net25 dvdd.t829 dvdd.t828 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X2294 por_ana_0.comparator_1.vnn avss.t439 por_ana_0.comparator_1.vt.t2 por_ana_0.comparator_1.vt.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=8
X2295 por_ana_0.comparator_1.vpp.t25 por_ana_0.comparator_1.vnn.t56 avdd.t642 avdd.t395 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X2296 por_dig_0.otrip_decoded[7].t0 a_37156_28013# dvss.t752 dvss.t523 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X2297 por_ana_0.rstring_mux_0.otrip_decoded_b_avdd[7] por_ana_0.rstring_mux_0.otrip_decoded_avdd[7] avdd.t436 avdd.t435 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X2298 por_dig_0.otrip_decoded[6].t2 a_35960_29101# dvdd.t1219 dvdd.t668 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X2299 dvdd.t543 por_dig_0.cnt_por\[0\].t20 por_dig_0._051_ dvdd.t542 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.165 ps=1.33 w=1 l=0.15
X2300 a_23734_21903# a_23366_22885# dvss.t906 dvss.t905 sky130_fd_pr__nfet_01v8 ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X2301 por_ana_0.comparator_1.vnn avss.t440 por_ana_0.comparator_1.vt.t1 por_ana_0.comparator_1.vt.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=8
X2302 por_dig_0.cnt_st\[0\] a_38320_34301# dvdd.t716 dvdd.t715 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X2303 a_39720_32365# por_dig_0.cnt_st\[1\] por_dig_0._041_ dvss.t598 sky130_fd_pr__nfet_01v8 ad=0.095875 pd=0.945 as=0.091 ps=0.93 w=0.65 l=0.15
X2304 por_ana_0.comparator_0.vinn.t1 avdd.t39 por_ana_0.comparator_0.vinn.t1 avdd.t40 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=0.6
X2305 a_35582_34317# por_dig_0._017_ dvss.t769 dvss.t768 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X2306 dvss.t710 por_dig_0.clknet_1_1__leaf_osc_ck.t44 a_32740_35091# dvss.t709 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2307 a_34990_30189# a_34946_30431# a_34824_30189# dvss.t913 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X2308 a_37212_31111# a_36696_30739# a_37117_31099# dvss.t1261 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X2309 por_dig_0._016_ por_dig_0._033_ dvdd.t25 dvdd.t24 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2310 dvdd.t1135 a_37614_32883# a_37504_32909# dvdd.t1134 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X2311 dvdd.t1754 dvss.t2320 dvdd.t1753 dvdd.t1556 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X2312 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[5].t0 a_35233_24371# avdd.t291 avdd.t286 sky130_fd_pr__pfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.24375 ps=1.825 w=1.5 l=0.5
X2313 a_33983_35085# a_32906_35091# a_33821_35463# dvdd.t1017 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X2314 a_32984_32339# a_32809_32365# a_33163_32365# dvss.t929 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X2315 avss.t293 por_ana_0.comparator_1.vn.t7 por_ana_0.comparator_1.vt.t54 avss.t292 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X2316 por_ana_0.comparator_0.vinn.t19 avss.t59 vin.t14 avss.t60 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X2317 dvdd.t314 a_33444_31037# a_33431_30733# dvdd.t313 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X2318 avss.t58 avss.t57 avss.t58 avss.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=8
X2319 dvss.t1745 dvdd.t1890 dvss.t1744 dvss.t1743 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X2320 a_23466_24707# a_23366_24619# dvss.t1518 dvss.t1517 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X2321 a_33654_33287# a_32464_32915# a_33545_33287# dvss.t469 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X2322 a_36743_35995# a_35666_35629# a_36581_35629# dvdd.t518 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X2323 avdd.t394 por_ana_0.comparator_1.vpp.t4 por_ana_0.comparator_1.vpp.t5 avdd.t392 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X2324 a_37614_33695# a_37396_33453# dvss.t1084 dvss.t917 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X2325 dvdd.t1131 a_34265_27987# por_dig_0.otrip_decoded[4] dvdd.t1130 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X2326 a_32182_21903# a_31814_22885# dvdd.t1484 dvdd.t1483 sky130_fd_pr__pfet_01v8_hvt ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X2327 dvdd.t463 a_36756_35603# por_dig_0.cnt_por\[0\].t5 dvdd.t462 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2328 a_2543_22912# a_2165_15512# avss.t27 sky130_fd_pr__res_xhigh_po_1p41 l=35
X2329 avdd.t267 a_34026_22973# a_34719_21859# avdd.t266 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.1365 ps=1.49 w=0.42 l=1
X2330 a_32182_23637# a_31814_24619# dvdd.t1386 dvdd.t1385 sky130_fd_pr__pfet_01v8_hvt ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X2331 a_37518_35463# a_36328_35091# a_37409_35463# dvss.t991 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X2332 a_32326_33453# por_dig_0.net24 dvss.t419 dvss.t418 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1346 ps=1.15 w=0.42 l=0.15
X2333 avss.t56 avss.t54 por_ana_0.ibias_gen_0.vr.t0 avss.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=4
X2334 dvdd.t1322 a_36328_29645# por_dig_0.net25 dvdd.t70 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2335 a_31890_33453# a_31412_33427# dvss.t2009 dvss.t2008 sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.12495 ps=1.015 w=0.42 l=0.15
X2336 a_39630_33229# por_dig_0._030_ dvss.t2190 dvss.t2189 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X2337 a_25724_13935# a_25346_6535# avss.t155 sky130_fd_pr__res_xhigh_po_1p41 l=35
X2338 dvdd.t895 a_35111_28013# a_35217_28013# dvdd.t894 sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X2339 dvss.t554 a_32794_33971# por_dig_0._012_ dvss.t553 sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X2340 vin.t26 por_ana_0.rstring_mux_0.otrip_decoded_avdd[3] por_ana_0.rstring_mux_0.vtrip3.t5 avss.t237 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X2341 avss.t348 por_ana_0.comparator_0.vm.t0 por_ana_0.comparator_0.vm.t1 avss.t100 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X2342 dvss.t184 a_34098_30707# por_dig_0.clknet_1_0__leaf_osc_ck.t2 dvss.t183 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2343 pwup_filt.t24 por_ana_0.sky130_fd_sc_hd__inv_4_0.Y dvdd.t211 dvdd.t210 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2344 dvss.t1742 dvdd.t1891 dvss.t1741 dvss.t1740 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X2345 avdd.t316 a_27690_24707# a_28383_23593# avdd.t315 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.1365 ps=1.49 w=0.42 l=1
X2346 avdd.t541 por_ana_0.comparator_1.n1.t16 por_ana_0.dcomp3v3 avdd.t540 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.6
X2347 a_21188_13935# a_20810_6535# avss.t156 sky130_fd_pr__res_xhigh_po_1p41 l=35
X2348 dvss.t1478 a_25478_24619# a_25578_24707# dvss.t1477 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X2349 a_32818_28013# a_32641_28013# dvdd.t825 dvdd.t824 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X2350 dvdd.t1406 a_34357_33427# por_dig_0._021_ dvdd.t1405 sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.265 ps=2.53 w=1 l=0.15
X2351 por_dig_0.clknet_0_osc_ck.t20 a_34387_32909# dvdd.t111 dvdd.t110 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2352 a_35918_35124# por_dig_0.net23.t19 a_35704_35124# dvdd.t766 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.1932 ps=1.34 w=0.42 l=0.15
X2353 dvss.t417 por_dig_0.net24 a_31650_33453# dvss.t416 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.06405 ps=0.725 w=0.42 l=0.15
X2354 dvss.t2057 a_31914_24707# a_33121_24371# dvss.t517 sky130_fd_pr__nfet_g5v0d10v5 ad=0.121875 pd=1.075 as=0.19875 ps=2.03 w=0.75 l=0.5
X2355 dvss.t916 a_38500_31251# a_38242_31251# dvss.t915 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.5
X2356 dvdd.t854 a_38974_34693# por_dig_0.net31 dvdd.t853 sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.26 ps=2.52 w=1 l=0.15
X2357 a_4811_22912# a_4433_15512# avss.t27 sky130_fd_pr__res_xhigh_po_1p41 l=35
X2358 dvdd.t209 por_ana_0.sky130_fd_sc_hd__inv_4_0.Y pwup_filt.t23 dvdd.t208 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2359 dvdd.t1369 por_dig_0.cnt_st\[2\] a_38926_33453# dvdd.t1368 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2360 a_35704_35124# por_dig_0.net23.t20 a_35704_35451# dvss.t885 sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X2361 por_dig_0.cnt_st\[2\] a_38136_33213# dvss.t1248 dvss.t283 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X2362 por_ana_0.comparator_0.vinn.t7 avdd.t37 vin.t2 avdd.t38 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X2363 dvdd.t529 por_dig_0.net26 a_32651_31643# dvdd.t528 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X2364 por_ana_0.ibias_gen_0.vp.t4 por_ana_0.ibias_gen_0.isrc_sel.t7 por_ana_0.ibias_gen_0.vp0.t10 avdd.t583 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X2365 a_33364_36173# a_32740_36179# a_33256_36551# dvdd.t374 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X2366 a_26271_23593# a_25846_23637# dvss.t362 dvss.t361 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X2367 dvss.t2000 a_36376_28789# por_dig_0.net16 dvss.t1999 sky130_fd_pr__nfet_01v8 ad=0.122275 pd=1.08 as=0.169 ps=1.82 w=0.65 l=0.15
X2368 a_25846_21903# a_25478_22885# dvss.t1558 dvss.t1557 sky130_fd_pr__nfet_01v8 ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X2369 a_18164_13935# a_17786_6535# avss.t157 sky130_fd_pr__res_xhigh_po_1p41 l=35
X2370 dvss.t1739 dvdd.t1892 dvss.t1738 dvss.t1737 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X2371 dvss.t127 a_39887_21959# a_40246_21893# dvss.t126 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.19875 ps=2.03 w=0.75 l=0.5
X2372 dvdd.t629 a_35674_28557# a_35774_28673# dvdd.t628 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1085 ps=1.36 w=0.42 l=0.15
X2373 dvdd.t804 a_34633_36147# por_dig_0._052_ dvdd.t803 sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.265 ps=2.53 w=1 l=0.15
X2374 a_37046_33453# a_36880_33453# dvss.t751 dvss.t520 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2375 dvss.t1028 a_39888_23693# a_40247_23627# dvss.t1027 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.19875 ps=2.03 w=0.75 l=0.5
X2376 por_ana_0.ibias_gen_0.isrc_sel_b.t0 avdd.t35 por_ana_0.ibias_gen_0.ena_b.t0 avdd.t36 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X2377 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[7].t0 a_37345_24371# avdd.t293 avdd.t292 sky130_fd_pr__pfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.24375 ps=1.825 w=1.5 l=0.5
X2378 avss.t199 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.t32 porb_h.t21 avss.t198 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X2379 por_dig_0.net28 a_31908_32909# dvdd.t1188 dvdd.t1187 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X2380 dvdd.t109 a_34387_32909# por_dig_0.clknet_0_osc_ck.t19 dvdd.t108 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X2381 a_19094_2382# a_41694_2760# dvss.t632 sky130_fd_pr__res_xhigh_po_1p41 l=111
X2382 por_ana_0.comparator_1.vnn.t17 por_ana_0.comparator_1.vpp.t61 avdd.t417 avdd.t403 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X2383 por_ana_0.comparator_0.vt.t6 por_ana_0.comparator_0.vinn.t59 por_ana_0.comparator_0.vnn por_ana_0.comparator_0.vt.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X2384 vin.t28 por_ana_0.rstring_mux_0.otrip_decoded_b_avdd[3] por_ana_0.rstring_mux_0.vtrip3.t7 avdd.t451 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X2385 por.t18 por_ana_0.sky130_fd_sc_hd__inv_4_4.Y dvdd.t952 dvdd.t951 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2386 dvss.t791 por_dig_0.net6 a_33155_28640# dvss.t790 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X2387 dvdd.t1473 a_36381_36691# por_dig_0.por_unbuf.t2 dvdd.t1472 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X2388 por_dig_0._039_ por_dig_0.net21 a_39554_33997# dvdd.t1381 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X2389 a_34010_31821# a_33774_31821# dvdd.t926 dvdd.t925 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.5
X2390 por_ana_0.comparator_1.vt.t45 vbg_1v2.t34 por_ana_0.comparator_1.vnn por_ana_0.comparator_1.vt.t41 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X2391 a_35699_33819# a_35573_33721# a_35295_33705# dvss.t1977 sky130_fd_pr__special_nfet_01v8 ad=0.0999 pd=0.985 as=0.0711 ps=0.755 w=0.36 l=0.15
X2392 porb.t19 por_ana_0.sky130_fd_sc_hd__inv_4_1.Y dvdd.t279 dvdd.t278 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2393 dvdd.t1756 dvss.t2321 dvdd.t1755 dvdd.t1609 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X2394 a_32506_32365# a_32462_32607# a_32340_32365# dvss.t1970 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X2395 a_34294_21903# a_33926_22885# dvdd.t515 dvdd.t514 sky130_fd_pr__pfet_01v8_hvt ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X2396 a_36100_32517# por_dig_0.cnt_por\[5\] a_36334_32365# dvss.t2080 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X2397 dvss.t1063 a_21254_22885# a_21354_22973# dvss.t1062 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X2398 a_39077_31527# por_dig_0._044_ a_38904_31277# dvss.t475 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X2399 dvss.t1019 a_36380_33971# por_dig_0.net22.t0 dvss.t1018 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.0567 ps=0.69 w=0.42 l=0.15
X2400 a_32550_32199# a_31360_31827# a_32441_32199# dvss.t30 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X2401 a_34294_23637# a_33926_24619# dvdd.t430 dvdd.t429 sky130_fd_pr__pfet_01v8_hvt ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X2402 por_ana_0.comparator_1.vt.t44 vbg_1v2.t35 por_ana_0.comparator_1.vnn por_ana_0.comparator_1.vt.t41 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X2403 dvss.t1736 dvdd.t1893 dvss.t1735 dvss.t1734 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X2404 por_dig_0.net19 por_dig_0._035_ dvss.t2064 dvss.t2063 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2405 a_38957_32883# por_dig_0.net4 a_39349_32909# dvdd.t76 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.155 ps=1.31 w=1 l=0.15
X2406 porb.t3 por_ana_0.sky130_fd_sc_hd__inv_4_1.Y dvss.t331 dvss.t330 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2407 a_35861_28917# a_35674_28557# a_35774_28673# dvss.t732 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.107825 ps=1.36 w=0.42 l=0.15
X2408 avdd.t393 por_ana_0.comparator_1.vpp.t2 por_ana_0.comparator_1.vpp.t3 avdd.t392 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X2409 a_33805_32339# por_dig_0.cnt_por\[7\] a_33934_32615# dvdd.t931 sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X2410 a_32535_28013# a_32358_28013# dvdd.t1514 dvdd.t1513 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X2411 por_dig_0._035_ por_dig_0.cnt_por\[4\] dvdd.t1253 dvdd.t1252 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X2412 a_36935_35629# por_dig_0.net24 dvss.t415 dvss.t414 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X2413 a_35597_31821# por_dig_0._036_.t8 a_35000_31795# dvdd.t1351 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.2125 ps=1.425 w=1 l=0.15
X2414 porb_h.t20 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.t33 avss.t201 avss.t200 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X2415 dvdd.t613 a_39328_34515# a_39070_34515# dvdd.t612 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.5
X2416 dvss.t861 por_dig_0.net7.t19 por_dig_0.net12 dvss.t523 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.08775 ps=0.92 w=0.65 l=0.15
X2417 a_33545_33287# a_32630_32915# a_33198_32883# dvss.t983 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X2418 dvss.t518 a_34026_24707# a_35233_24371# dvss.t517 sky130_fd_pr__nfet_g5v0d10v5 ad=0.121875 pd=1.075 as=0.19875 ps=2.03 w=0.75 l=0.5
X2419 dvdd.t1758 dvss.t2322 dvdd.t1757 dvdd.t1522 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X2420 dvss.t542 a_35468_30163# a_35402_30189# dvss.t541 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X2421 a_39728_31527# por_dig_0._043_ dvdd.t1308 dvdd.t1307 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X2422 por_ana_0.comparator_1.vt.t43 vbg_1v2.t36 por_ana_0.comparator_1.vnn por_ana_0.comparator_1.vt.t41 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X2423 dvdd.t1760 dvss.t2323 dvdd.t1759 dvdd.t1666 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X2424 por_ana_0.comparator_0.vnn.t29 por_ana_0.comparator_0.vinn.t60 por_ana_0.comparator_0.vt.t5 por_ana_0.comparator_0.vt.t3 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X2425 a_28383_23593# a_27958_23637# dvss.t781 dvss.t780 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X2426 por_ana_0.ibias_gen_0.vp1.t15 por_ana_0.ibias_gen_0.isrc_sel.t8 por_ana_0.ibias_gen_0.vp.t5 avss.t343 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X2427 avdd.t225 por_ana_0.rstring_mux_0.ena_b por_ana_0.rstring_mux_0.vtop.t3 avdd.t224 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X2428 por_dig_0.net13 a_33155_28640# a_33418_28557# dvdd.t1197 sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.135 ps=1.27 w=1 l=0.15
X2429 dvss.t1733 dvdd.t1894 dvss.t1732 dvss.t1682 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X2430 a_27958_21903# a_27590_22885# dvss.t1367 dvss.t1366 sky130_fd_pr__nfet_01v8 ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X2431 a_35836_31277# a_35390_31277# a_35740_31277# dvss.t924 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X2432 avss.t53 avss.t52 avss.t53 avss.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=8
X2433 a_21354_22973# a_21254_22885# dvss.t1061 dvss.t1060 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X2434 a_37409_35463# a_36494_35091# a_37062_35059# dvss.t995 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X2435 dvdd.t231 a_38136_33427# a_38123_33819# dvdd.t230 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X2436 por_ana_0.comparator_1.vt.t42 vbg_1v2.t37 por_ana_0.comparator_1.vnn por_ana_0.comparator_1.vt.t41 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X2437 dvdd.t255 a_38228_30163# a_38215_30555# dvdd.t254 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X2438 a_39630_33229# por_dig_0._039_ por_dig_0._002_ dvss.t1959 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2439 dvss.t1731 dvdd.t1895 dvss.t1730 dvss.t1729 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X2440 dvdd.t1503 a_35000_31795# por_dig_0._028_ dvdd.t1502 sky130_fd_pr__pfet_01v8_hvt ad=0.3825 pd=1.765 as=0.26 ps=2.52 w=1 l=0.15
X2441 por_ana_0.comparator_0.vt.t38 vbg_1v2.t38 por_ana_0.comparator_0.vpp.t30 por_ana_0.comparator_0.vt.t36 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X2442 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[0] a_31009_22637# dvss.t2194 dvss.t2193 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.121875 ps=1.075 w=0.75 l=0.5
X2443 por_ana_0.comparator_0.vnn.t30 por_ana_0.comparator_0.vinn.t61 por_ana_0.comparator_0.vt.t4 por_ana_0.comparator_0.vt.t3 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X2444 avss.t279 por_ana_0.comparator_0.n1.t16 por_ana_0.dcomp3v3uv avss.t278 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.6
X2445 dvss.t1728 dvdd.t1896 dvss.t1727 dvss.t1726 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X2446 a_37763_35451# por_dig_0.net24 dvss.t413 dvss.t412 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X2447 dvdd.t902 por_dig_0._024_ a_33012_33997# dvdd.t901 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X2448 por_ana_0.ibias_gen_0.isrc_sel.t0 a_39457_24371# avdd.t295 avdd.t294 sky130_fd_pr__pfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.24375 ps=1.825 w=1.5 l=0.5
X2449 a_17398_35244# a_17776_27844# avss.t158 sky130_fd_pr__res_xhigh_po_1p41 l=35
X2450 dvdd.t1762 dvss.t2324 dvdd.t1761 dvdd.t1556 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X2451 por_dig_0._043_ a_39497_30849# dvss.t1967 dvss.t1966 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X2452 a_32398_33453# a_32019_33819# a_32326_33453# dvss.t1582 sky130_fd_pr__nfet_01v8 ad=0.1401 pd=1.1 as=0.0441 ps=0.63 w=0.42 l=0.15
X2453 dcomp.t5 por_ana_0.sky130_fd_sc_hd__inv_4_3.Y dvss.t59 dvss.t58 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2454 por_ana_0.comparator_0.vt.t37 vbg_1v2.t39 por_ana_0.comparator_0.vpp.t31 por_ana_0.comparator_0.vt.t36 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X2455 dvdd.t207 por_ana_0.sky130_fd_sc_hd__inv_4_0.Y pwup_filt.t22 dvdd.t206 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2456 dvss.t1 por_dig_0.cnt_rsb a_34510_31277# dvss.t0 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2457 dvss.t644 por_dig_0.cnt_por\[0\].t21 a_35925_35451# dvss.t643 sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.0693 ps=0.75 w=0.42 l=0.15
X2458 dvdd.t753 por_dig_0._034_.t15 a_36962_32615# dvdd.t752 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X2459 por_ana_0.comparator_0.vnn.t42 por_ana_0.comparator_0.vnn.t41 avdd.t359 avdd.t182 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X2460 dvdd.t670 por_dig_0.net6 a_33155_28640# dvdd.t669 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.1092 ps=1.36 w=0.42 l=0.15
X2461 por_ana_0.sky130_fd_sc_hd__inv_4_1.Y por_ana_0.sky130_fd_sc_hd__inv_4_1.A dvss.t222 dvss.t221 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2462 a_36376_28789# a_36649_28789# dvdd.t1392 dvdd.t1391 sky130_fd_pr__pfet_01v8_hvt ad=0.1085 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2463 porb.t2 por_ana_0.sky130_fd_sc_hd__inv_4_1.Y dvss.t329 dvss.t328 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2464 dvss.t1013 a_37584_35389# por_dig_0.cnt_por\[1\] dvss.t1012 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2465 avss.t203 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.t34 porb_h.t19 avss.t202 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X2466 a_36406_21903# a_36038_22885# dvdd.t229 dvdd.t228 sky130_fd_pr__pfet_01v8_hvt ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X2467 a_32906_36179# a_32740_36179# dvdd.t373 dvdd.t372 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2468 dvss.t57 por_ana_0.sky130_fd_sc_hd__inv_4_3.Y dcomp.t4 dvss.t56 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2469 dvss.t904 a_23366_22885# a_23466_22973# dvss.t903 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X2470 dvss.t1594 dvss.t1592 force_dis_rc_osc.t0 dvss.t1593 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X2471 por_dig_0._048_ por_dig_0.net22.t21 dvdd.t611 dvdd.t610 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2472 por_ana_0.rstring_mux_0.vtrip3.t0 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[3] por_ana_0.comparator_0.vinn.t8 avss.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X2473 a_36406_23637# a_36038_24619# dvdd.t577 dvdd.t576 sky130_fd_pr__pfet_01v8_hvt ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X2474 a_21178_35244# por_ana_0.schmitt_trigger_0.in.t0 avss.t352 sky130_fd_pr__res_xhigh_po_1p41 l=35
X2475 a_36669_31821# por_dig_0._035_ a_36567_31821# dvdd.t1389 sky130_fd_pr__pfet_01v8_hvt ad=0.21 pd=1.42 as=0.18 ps=1.36 w=1 l=0.15
X2476 a_37820_13935# a_38198_6535# avss.t353 sky130_fd_pr__res_xhigh_po_1p41 l=35
X2477 dvdd.t625 a_40246_23089# a_40246_21893# dvdd.t624 sky130_fd_pr__pfet_01v8_hvt ad=0.2968 pd=2.77 as=0.2968 ps=2.77 w=1.12 l=0.15
X2478 dvss.t327 por_ana_0.sky130_fd_sc_hd__inv_4_1.Y porb.t1 dvss.t326 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2479 osc_ck.t6 por_ana_0.rc_osc_0.n.t11 dvdd.t1359 dvdd.t1358 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X2480 dvdd.t155 a_34098_30707# por_dig_0.clknet_1_0__leaf_osc_ck.t19 dvdd.t154 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2481 dvdd.t1764 dvss.t2325 dvdd.t1763 dvdd.t1593 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X2482 dvss.t1725 dvdd.t1897 dvss.t1724 dvss.t1723 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X2483 por_ana_0.comparator_0.vt.t23 avss.t441 por_ana_0.comparator_0.vnn.t16 por_ana_0.comparator_0.vt.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=8
X2484 a_36381_36691# por_dig_0.net20.t8 dvdd.t1429 dvdd.t1428 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X2485 a_34754_35451# por_dig_0.cnt_por\[1\] a_34672_35451# dvss.t1397 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.1092 ps=1.36 w=0.42 l=0.15
X2486 por_ana_0.comparator_0.n0.t4 por_ana_0.comparator_0.ena_b.t4 avss.t334 avss.t45 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X2487 por_ana_0.rstring_mux_0.vtrip_decoded_b_avdd[6] por_ana_0.rstring_mux_0.vtrip_decoded_avdd[6].t5 avss.t213 avss.t212 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X2488 a_36831_21859# a_36406_21903# dvss.t1308 dvss.t1307 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X2489 a_35592_36286# por_dig_0.cnt_por\[0\].t22 dvdd.t545 dvdd.t544 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X2490 a_32603_31821# a_31526_31827# a_32441_32199# dvdd.t945 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X2491 por_ana_0.comparator_0.vm.t4 por_ana_0.comparator_0.vnn.t61 avdd.t376 avdd.t191 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X2492 dvss.t1984 a_36328_29645# por_dig_0.net25 dvss.t1983 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2493 avdd.t502 por_ana_0.comparator_0.n0.t7 por_ana_0.comparator_0.n1.t2 avdd.t501 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X2494 dvdd.t1767 dvss.t2326 dvdd.t1766 dvdd.t1765 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X2495 por_ana_0.comparator_0.vnn.t40 por_ana_0.comparator_0.vnn.t39 avdd.t358 avdd.t182 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X2496 por_dig_0.net25 a_36328_29645# dvdd.t1321 dvdd.t70 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X2497 por_ana_0.comparator_1.vm.t0 por_ana_0.comparator_1.vnn.t57 avdd.t643 avdd.t395 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X2498 dvss.t686 a_36138_24707# a_37345_24371# dvss.t517 sky130_fd_pr__nfet_g5v0d10v5 ad=0.121875 pd=1.075 as=0.19875 ps=2.03 w=0.75 l=0.5
X2499 dvdd.t768 por_dig_0.net23.t21 a_35592_36286# dvdd.t767 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X2500 por_dig_0.net8 a_32004_30189# dvss.t1417 dvss.t1416 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2501 a_35295_33705# a_35612_33595# a_35570_33453# dvss.t1470 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0669 ps=0.75 w=0.36 l=0.15
X2502 avss.t11 por_ana_0.comparator_1.n1.t17 por_ana_0.dcomp3v3 avss.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X2503 dvdd.t992 a_32088_33690# a_32019_33819# dvdd.t991 sky130_fd_pr__pfet_01v8_hvt ad=0.2184 pd=2.2 as=0.12915 ps=1.185 w=0.84 l=0.15
X2504 a_35556_29619# por_dig_0.cnt_por\[9\] dvdd.t1499 dvdd.t325 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2505 dvdd.t205 por_ana_0.sky130_fd_sc_hd__inv_4_0.Y pwup_filt.t21 dvdd.t204 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2506 dvdd.t1770 dvss.t2327 dvdd.t1769 dvdd.t1768 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X2507 a_32441_32199# a_31526_31827# a_32094_31795# dvss.t1134 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X2508 dvdd.t1339 por_dig_0.net16 a_36512_28013# dvdd.t1338 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X2509 a_23466_22973# a_23366_22885# dvss.t902 dvss.t901 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X2510 a_32906_35091# a_32740_35091# dvdd.t1032 dvdd.t1031 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2511 por_dig_0.clknet_0_osc_ck.t18 a_34387_32909# dvdd.t107 dvdd.t106 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2512 avdd.t626 por_ana_0.comparator_1.vnn.t2 por_ana_0.comparator_1.vnn.t3 avdd.t401 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X2513 a_38986_34317# por_dig_0.net31 por_dig_0._000_ dvss.t970 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2514 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[2] a_33121_22637# dvss.t1254 dvss.t1253 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.121875 ps=1.075 w=0.75 l=0.5
X2515 por_ana_0.rstring_mux_0.vtrip3.t2 por_ana_0.rstring_mux_0.vtrip_decoded_b_avdd[3] por_ana_0.comparator_0.vinn.t10 avdd.t260 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X2516 vin.t15 avss.t50 vin.t15 avss.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=0.6
X2517 dvss.t572 a_35583_34541# por_dig_0.clknet_1_1__leaf_osc_ck.t3 dvss.t571 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2518 dvss.t411 por_dig_0.net24 a_32506_32365# dvss.t410 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X2519 dvss.t1722 dvdd.t1898 dvss.t1721 dvss.t1720 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X2520 a_32701_28531# por_dig_0.net12 dvdd.t405 dvdd.t404 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X2521 avdd.t34 avdd.t32 avdd.t34 avdd.t33 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=8
X2522 dvdd.t603 por_dig_0.clknet_1_1__leaf_osc_ck.t45 a_35500_35629# dvdd.t602 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X2523 dvss.t485 a_29702_22885# a_29802_22973# dvss.t484 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X2524 dvdd.t1772 dvss.t2328 dvdd.t1771 dvdd.t1700 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X2525 por_ana_0.comparator_1.vpp.t46 vin.t65 por_ana_0.comparator_1.vt.t19 por_ana_0.comparator_1.vt.t18 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X2526 a_32922_30707# a_32704_31111# dvss.t940 dvss.t939 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X2527 dvss.t1719 dvdd.t1899 dvss.t1718 dvss.t1717 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X2528 avdd.t190 por_ana_0.comparator_0.vpp.t54 por_ana_0.comparator_0.vnn.t8 avdd.t180 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X2529 dvss.t228 por_ana_0.sky130_fd_sc_hd__inv_4_0.Y pwup_filt.t0 dvss.t227 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2530 dvdd.t939 por_dig_0._048_ por_dig_0._011_ dvdd.t938 sky130_fd_pr__pfet_01v8_hvt ad=0.182 pd=1.92 as=0.174 ps=1.39 w=0.7 l=0.15
X2531 por_ana_0.rstring_mux_0.otrip_decoded_b_avdd[0] por_ana_0.rstring_mux_0.otrip_decoded_avdd[0] avdd.t508 avdd.t507 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X2532 dvdd.t1038 a_32984_32339# a_32971_32731# dvdd.t1037 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X2533 por_ana_0.schmitt_trigger_0.in.t14 dvss.t659 sky130_fd_pr__cap_mim_m3_2 l=30 w=30
X2534 a_38518_21903# a_38150_22885# dvdd.t95 dvdd.t94 sky130_fd_pr__pfet_01v8_hvt ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X2535 por_ana_0.sky130_fd_sc_hd__inv_4_4.Y por_dig_0.por_unbuf.t19 dvdd.t696 dvdd.t695 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2536 por.t17 por_ana_0.sky130_fd_sc_hd__inv_4_4.Y dvdd.t950 dvdd.t949 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2537 dvss.t1556 a_25478_22885# a_25578_22973# dvss.t1555 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X2538 a_35933_28917# por_dig_0.net6 a_35861_28917# dvss.t789 sky130_fd_pr__nfet_01v8 ad=0.05355 pd=0.675 as=0.0441 ps=0.63 w=0.42 l=0.15
X2539 dvdd.t1414 a_31932_33595# a_31893_33721# dvdd.t1413 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X2540 dvdd.t1775 dvss.t2329 dvdd.t1774 dvdd.t1773 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X2541 por_ana_0.comparator_0.vnn.t7 por_ana_0.comparator_0.vpp.t55 avdd.t189 avdd.t182 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X2542 por_ana_0.rstring_mux_0.vtrip_decoded_b_avdd[0] por_ana_0.rstring_mux_0.vtrip_decoded_avdd[0] avss.t220 avss.t219 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X2543 a_38518_23637# a_38150_24619# dvdd.t35 dvdd.t34 sky130_fd_pr__pfet_01v8_hvt ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X2544 a_37614_33695# a_37396_33453# dvdd.t922 dvdd.t921 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X2545 porb.t18 por_ana_0.sky130_fd_sc_hd__inv_4_1.Y dvdd.t277 dvdd.t276 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2546 a_14374_35244# por_ana_0.vl avss.t354 sky130_fd_pr__res_xhigh_po_1p41 l=35
X2547 dvdd.t1050 a_38136_33213# a_38123_32909# dvdd.t1049 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X2548 dvdd.t75 por_dig_0.net4 a_35597_31821# dvdd.t74 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.105 ps=1.21 w=1 l=0.15
X2549 dvss.t2001 por_dig_0.net16 a_36512_28013# dvss.t677 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X2550 dvdd.t1777 dvss.t2330 dvdd.t1776 dvdd.t1522 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X2551 por_ana_0.rstring_mux_0.vtrip_decoded_b_avdd[7] por_ana_0.rstring_mux_0.vtrip_decoded_avdd[7].t5 avdd.t620 avdd.t619 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X2552 avss.t205 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.t35 porb_h.t18 avss.t204 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X2553 dvss.t1469 a_35612_33595# a_35573_33721# dvss.t1468 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2554 por.t0 por_ana_0.sky130_fd_sc_hd__inv_4_4.Y dvss.t1137 dvss.t1136 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2555 por_dig_0.force_pdnb a_31413_29075# dvss.t2229 dvss.t2228 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X2556 dvdd.t948 por_ana_0.sky130_fd_sc_hd__inv_4_4.Y por.t16 dvdd.t947 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2557 por_ana_0.comparator_0.vt.t22 avss.t442 por_ana_0.comparator_0.vnn.t15 por_ana_0.comparator_0.vt.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=8
X2558 dvdd.t263 por_dig_0.cnt_por\[8\] a_33774_31821# dvdd.t262 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2559 a_38943_21859# a_38518_21903# dvss.t260 dvss.t259 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X2560 dvdd.t275 por_ana_0.sky130_fd_sc_hd__inv_4_1.Y porb.t17 dvdd.t274 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2561 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[5].t1 a_35233_24371# dvss.t628 dvss.t517 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.121875 ps=1.075 w=0.75 l=0.5
X2562 dvss.t1075 a_21254_24619# a_21354_24707# dvss.t1074 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X2563 por_ana_0.comparator_0.vinn.t37 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[5].t5 por_ana_0.rstring_mux_0.vtrip5.t9 avss.t303 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X2564 dvss.t734 por_dig_0._021_ a_34109_33453# dvss.t733 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X2565 vin.t3 avdd.t30 vin.t3 avdd.t31 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=0.6
X2566 avdd.t29 avdd.t26 avdd.t28 avdd.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=8
X2567 a_34040_13935# a_34418_6535# avss.t355 sky130_fd_pr__res_xhigh_po_1p41 l=35
X2568 dvss.t139 a_34387_32909# por_dig_0.clknet_0_osc_ck.t2 dvss.t138 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2569 por_dig_0.net11 por_dig_0.net5.t17 dvss.t2124 dvss.t2123 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2570 por_dig_0.cnt_rsb a_32616_32125# dvss.t466 dvss.t465 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X2571 avdd.t188 por_ana_0.comparator_0.vpp.t56 por_ana_0.comparator_0.vnn.t6 avdd.t180 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X2572 por_dig_0._034_.t3 por_dig_0.cnt_por\[0\].t23 dvdd.t547 dvdd.t546 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.215 ps=1.43 w=1 l=0.15
X2573 a_33378_31111# a_32188_30739# a_33269_31111# dvss.t935 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X2574 dvss.t55 por_ana_0.sky130_fd_sc_hd__inv_4_3.Y dcomp.t3 dvss.t54 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2575 a_27690_22973# a_27590_22885# dvss.t1365 dvss.t1364 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X2576 a_16642_35244# a_16264_27844# avss.t356 sky130_fd_pr__res_xhigh_po_1p41 l=35
X2577 dvdd.t1070 a_33996_35389# a_33983_35085# dvdd.t1069 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X2578 a_32138_32187# a_32094_31795# a_31972_32199# dvss.t2211 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X2579 dvss.t119 por_dig_0._037_ por_dig_0.net19 dvss.t118 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2580 a_37750_30189# a_37706_30431# a_37584_30189# dvss.t900 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X2581 por_ana_0.comparator_0.vnn.t5 por_ana_0.comparator_0.vpp.t57 avdd.t187 avdd.t182 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X2582 a_35552_13935# a_35174_6535# avss.t357 sky130_fd_pr__res_xhigh_po_1p41 l=35
X2583 a_35921_35629# por_dig_0._005_ dvdd.t573 dvdd.t572 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X2584 dvss.t325 por_ana_0.sky130_fd_sc_hd__inv_4_1.Y porb.t0 dvss.t324 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2585 a_25578_22973# a_25478_22885# dvss.t1554 dvss.t1553 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X2586 dvss.t1716 dvdd.t1900 dvss.t1715 dvss.t1714 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X2587 por_dig_0.clknet_1_1__leaf_osc_ck.t16 a_35583_34541# dvdd.t471 dvdd.t470 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2588 a_38320_34301# a_38145_34375# a_38499_34363# dvss.t914 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X2589 avss.t406 por_ana_0.ibias_gen_0.vn1.t16 por_ana_0.ibias_gen_0.vp1.t3 avss.t396 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=8
X2590 por_dig_0.net12 por_dig_0.net6 dvss.t788 dvss.t523 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2591 dvss.t1713 dvdd.t1901 dvss.t1712 dvss.t1711 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X2592 avdd.t440 a_38250_24707# a_39457_24371# avdd.t439 sky130_fd_pr__pfet_g5v0d10v5 ad=0.24375 pd=1.825 as=0.3975 ps=3.53 w=1.5 l=0.5
X2593 porb_h.t17 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.t36 avss.t207 avss.t206 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.19875 ps=2.03 w=0.75 l=0.5
X2594 dvss.t1461 a_25495_33620# a_25595_33708# dvss.t1460 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X2595 dvdd.t898 a_40246_21893# por_ana_0.sky130_fd_sc_hvl__lsbufhv2lv_1_1.X dvdd.t624 sky130_fd_pr__pfet_01v8_hvt ad=0.1568 pd=1.4 as=0.2968 ps=2.77 w=1.12 l=0.15
X2596 dvss.t2125 por_dig_0.net5.t18 a_35930_28013# dvss.t677 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X2597 a_20422_35244# a_20044_27844# avss.t358 sky130_fd_pr__res_xhigh_po_1p41 l=35
X2598 avdd.t578 por_ana_0.ibias_gen_0.isrc_sel_b.t8 por_ana_0.ibias_gen_0.vp0.t9 avdd.t577 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X2599 dvdd.t182 por_dig_0.net29 a_34578_29645# dvdd.t70 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2600 dvss.t2160 a_31814_22885# a_31914_22973# dvss.t2159 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X2601 a_38070_33453# a_36880_33453# a_37961_33453# dvss.t519 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X2602 a_26288_32594# a_25863_32638# dvss.t536 dvss.t535 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X2603 a_33418_28557# por_dig_0.net5.t19 a_33334_28557# dvdd.t1449 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2604 a_34467_28557# a_34290_28557# dvss.t972 dvss.t971 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X2605 por_ana_0.comparator_0.vt.t2 por_ana_0.comparator_0.vinn.t62 por_ana_0.comparator_0.vnn por_ana_0.comparator_0.vt.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X2606 a_21354_24707# a_21254_24619# dvss.t1073 dvss.t1072 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X2607 dvss.t1710 dvdd.t1902 dvss.t1709 dvss.t1682 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X2608 dvss.t1591 dvss.t1589 a_31814_24619# dvss.t1590 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X2609 a_18910_35244# a_18532_27844# avss.t359 sky130_fd_pr__res_xhigh_po_1p41 l=35
X2610 por_ana_0.comparator_0.vinn.t28 por_ana_0.rstring_mux_0.vtrip_decoded_b_avdd[5] por_ana_0.rstring_mux_0.vtrip5.t2 avdd.t458 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X2611 dvss.t1230 a_21622_23637# a_22047_23593# dvss.t1229 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X2612 dvdd.t1463 por_dig_0.clknet_0_osc_ck.t44 a_34098_30707# dvdd.t1462 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X2613 por_ana_0.comparator_1.n1.t2 por_ana_0.comparator_1.n0.t8 avss.t146 avss.t145 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.6
X2614 por_ana_0.rstring_mux_0.vtrip5.t4 por_ana_0.rstring_mux_0.otrip_decoded_avdd[5] vin.t30 avss.t259 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X2615 por_ana_0.comparator_0.vpp.t45 por_ana_0.comparator_0.vnn.t62 avdd.t377 avdd.t191 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X2616 por_dig_0.net18 a_35776_28013# dvss.t1485 dvss.t523 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X2617 por_dig_0.otrip_decoded[4] a_34265_27987# dvss.t1360 dvss.t523 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X2618 dvdd.t1333 a_33806_33427# por_dig_0._010_ dvdd.t1332 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2619 dvss.t125 a_39887_21959# a_40246_21893# dvss.t124 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.19875 ps=2.03 w=0.75 l=0.5
X2620 avdd.t625 por_ana_0.comparator_1.vnn.t0 por_ana_0.comparator_1.vnn.t1 avdd.t401 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X2621 por_dig_0.cnt_por\[0\].t0 a_36756_35603# dvss.t556 dvss.t555 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2622 por_dig_0._045_ a_37789_31821# dvdd.t1145 dvdd.t1144 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.3275 ps=1.655 w=1 l=0.15
X2623 dvss.t1363 a_27590_22885# a_27690_22973# dvss.t1362 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X2624 a_35455_30555# a_34378_30189# a_35293_30189# dvdd.t1120 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X2625 a_38315_33275# por_dig_0.net24 dvss.t409 dvss.t408 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X2626 por_dig_0._013_ a_34444_32517# dvdd.t911 dvdd.t910 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.36 ps=2.72 w=1 l=0.15
X2627 por_ana_0.comparator_0.vt.t1 por_ana_0.comparator_0.vinn.t63 por_ana_0.comparator_0.vnn por_ana_0.comparator_0.vt.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X2628 a_37688_33997# por_dig_0.net25 dvdd.t827 dvdd.t826 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X2629 avdd.t357 por_ana_0.comparator_0.vnn.t37 por_ana_0.comparator_0.vnn.t38 avdd.t180 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X2630 avdd.t25 avdd.t23 avdd.t25 avdd.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=4
X2631 vin.t24 por_ana_0.rstring_mux_0.otrip_decoded_avdd[7] por_ana_0.rstring_mux_0.vtrip7.t2 avss.t226 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X2632 dvss.t53 por_ana_0.sky130_fd_sc_hd__inv_4_3.Y dcomp.t2 dvss.t52 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2633 a_31615_31529# a_31893_31545# a_31849_31643# dvdd.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0567 ps=0.69 w=0.42 l=0.15
X2634 por_ana_0.dcomp3v3uv por_ana_0.comparator_0.n1.t17 avss.t281 avss.t280 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X2635 pwup_filt.t20 por_ana_0.sky130_fd_sc_hd__inv_4_0.Y dvdd.t203 dvdd.t202 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2636 dvdd.t1779 dvss.t2331 dvdd.t1778 dvdd.t1522 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X2637 avdd.t644 por_ana_0.comparator_1.vnn.t58 por_ana_0.comparator_1.vpp.t26 avdd.t392 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X2638 a_25595_33708# a_25495_33620# dvss.t1459 dvss.t1458 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X2639 a_34026_22973# a_33926_22885# dvss.t610 dvss.t609 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X2640 a_38622_31053# por_dig_0.net4 dvss.t86 dvss.t85 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2641 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[7].t1 a_37345_24371# dvss.t629 dvss.t517 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.121875 ps=1.075 w=0.75 l=0.5
X2642 dvss.t1516 a_23366_24619# a_23466_24707# dvss.t1515 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X2643 dvss.t646 por_dig_0.cnt_por\[0\].t24 a_35450_35124# dvss.t645 sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.1092 ps=1.36 w=0.42 l=0.15
X2644 dvss.t1247 a_38136_33213# a_38070_33287# dvss.t285 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X2645 a_25595_33708# a_25495_33620# dvss.t1457 dvss.t1456 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X2646 dvss.t407 por_dig_0.net24 a_37658_33275# dvss.t406 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X2647 dvss.t712 por_dig_0.clknet_1_1__leaf_osc_ck.t46 a_35500_35629# dvss.t711 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2648 dvss.t716 por_dig_0.net22.t22 a_33686_34335# dvss.t715 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X2649 dvss.t534 a_25863_32638# a_26288_32594# dvss.t533 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X2650 dvss.t1566 a_35640_32517# por_dig_0._017_ dvss.t1565 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X2651 avdd.t22 avdd.t20 avdd.t21 avdd.t3 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=8
X2652 dvss.t1708 dvdd.t1903 dvss.t1707 dvss.t1706 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X2653 a_22047_23593# a_21622_23637# dvss.t1228 dvss.t1227 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X2654 avdd.t356 por_ana_0.comparator_0.vnn.t35 por_ana_0.comparator_0.vnn.t36 avdd.t180 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X2655 dvdd.t1314 a_38444_28013# por_dig_0.otrip_decoded[0].t2 dvdd.t1313 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X2656 por_dig_0.cnt_por\[5\] a_33720_33213# dvdd.t641 dvdd.t640 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X2657 dvdd.t1044 a_35100_32339# por_dig_0.net24 dvdd.t1043 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.14 ps=1.28 w=1 l=0.15
X2658 por_ana_0.rstring_mux_0.vtrip5.t6 por_ana_0.rstring_mux_0.otrip_decoded_b_avdd[5] vin.t32 avdd.t468 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X2659 a_34114_35879# por_dig_0.cnt_por\[0\].t25 dvdd.t549 dvdd.t548 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X2660 por_dig_0.net25 a_36328_29645# dvss.t1982 dvss.t1981 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06825 ps=0.745 w=0.42 l=0.15
X2661 a_38986_31527# por_dig_0.net34 dvdd.t866 dvdd.t865 sky130_fd_pr__pfet_01v8_hvt ad=0.1525 pd=1.305 as=0.26 ps=2.52 w=1 l=0.15
X2662 dvdd.t906 a_33805_32339# por_dig_0._024_ dvdd.t905 sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.265 ps=2.53 w=1 l=0.15
X2663 a_35000_31795# por_dig_0.cnt_por\[9\] dvdd.t1498 dvdd.t1497 sky130_fd_pr__pfet_01v8_hvt ad=0.2175 pd=1.435 as=0.3825 ps=1.765 w=1 l=0.15
X2664 a_37676_34375# a_37230_34003# a_37580_34375# dvss.t1055 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X2665 avdd.t462 a_22047_23593# a_21354_24707# avdd.t461 sky130_fd_pr__pfet_g5v0d10v5 ad=0.2142 pd=1.99 as=0.2142 ps=1.99 w=0.42 l=1
X2666 avdd.t645 por_ana_0.comparator_1.vnn.t59 por_ana_0.comparator_1.vpp.t27 avdd.t392 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X2667 por_ana_0.comparator_0.ibias.t1 por_ana_0.ibias_gen_0.vp.t12 avdd.t389 avdd.t388 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X2668 vin.t48 por_ana_0.rstring_mux_0.otrip_decoded_b_avdd[7] por_ana_0.rstring_mux_0.vtrip7.t8 avdd.t653 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X2669 dvss.t1486 a_37800_28013# por_dig_0.otrip_decoded[3].t0 dvss.t523 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X2670 a_35556_29619# por_dig_0.cnt_por\[9\] dvss.t2185 dvss.t2184 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2671 por_dig_0.clknet_1_0__leaf_osc_ck.t1 a_34098_30707# dvss.t182 dvss.t181 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2672 por_ana_0.rstring_mux_0.vtrip7.t7 por_ana_0.rstring_mux_0.vtrip6.t5 avss.t360 sky130_fd_pr__res_xhigh_po_1p41 l=35
X2673 por_ana_0.sky130_fd_sc_hd__inv_4_0.Y por_ana_0.schmitt_trigger_0.out.t14 dvss.t826 dvss.t825 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2674 avdd.t543 por_ana_0.comparator_1.n1.t18 por_ana_0.dcomp3v3 avdd.t542 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X2675 dvss.t714 por_dig_0.clknet_1_1__leaf_osc_ck.t47 a_36328_35091# dvss.t713 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2676 dvss.t608 a_33926_22885# a_34026_22973# dvss.t607 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X2677 dvdd.t407 por_dig_0._044_ a_39077_31527# dvdd.t406 sky130_fd_pr__pfet_01v8_hvt ad=0.3275 pd=1.655 as=0.195 ps=1.39 w=1 l=0.15
X2678 por_ana_0.ibias_gen_0.vp1.t2 por_ana_0.ibias_gen_0.vn1.t17 avss.t407 avss.t398 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=8
X2679 a_37571_35085# a_36494_35091# a_37409_35463# dvdd.t873 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X2680 por_dig_0.clknet_0_osc_ck.t17 a_34387_32909# dvdd.t105 dvdd.t104 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2681 a_23466_24707# a_23366_24619# dvss.t1514 dvss.t1513 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X2682 por_ana_0.dcomp3v3 por_ana_0.comparator_1.n1.t19 avdd.t539 avdd.t538 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X2683 por_dig_0.clknet_0_osc_ck.t16 a_34387_32909# dvdd.t103 dvdd.t102 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2684 avdd.t19 avdd.t17 avdd.t18 avdd.t3 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=8
X2685 dvss.t1588 dvss.t1586 a_33926_24619# dvss.t1587 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X2686 dvss.t2139 por_dig_0.clknet_0_osc_ck.t45 a_35583_34541# dvss.t2138 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2687 a_38407_30189# por_dig_0.net25 dvss.t947 dvss.t946 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X2688 por_ana_0.rc_osc_0.vr a_41694_3516# dvss.t2025 sky130_fd_pr__res_xhigh_po_1p41 l=111
X2689 dvss.t1125 a_23734_23637# a_24159_23593# dvss.t1124 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X2690 a_33269_31111# a_32354_30739# a_32922_30707# dvss.t2232 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X2691 por_dig_0.por_unbuf.t0 a_36381_36691# dvss.t2148 dvss.t2147 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X2692 dvss.t570 a_35583_34541# por_dig_0.clknet_1_1__leaf_osc_ck.t2 dvss.t569 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2693 a_29504_13935# a_29882_6535# avss.t361 sky130_fd_pr__res_xhigh_po_1p41 l=35
X2694 dvss.t1705 dvdd.t1904 dvss.t1704 dvss.t1703 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X2695 dvss.t828 por_ana_0.schmitt_trigger_0.out.t15 por_ana_0.sky130_fd_sc_hd__inv_4_0.Y dvss.t827 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2696 dvss.t483 a_29702_22885# a_29802_22973# dvss.t482 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X2697 dvss.t1585 dvss.t1583 por_ana_0.schmitt_trigger_0.m.t12 dvss.t1584 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X2698 dvss.t568 a_35583_34541# por_dig_0.clknet_1_1__leaf_osc_ck.t1 dvss.t567 sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X2699 por_ana_0.rstring_mux_0.otrip_decoded_avdd[0] a_22561_22637# avdd.t310 avdd.t309 sky130_fd_pr__pfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.24375 ps=1.825 w=1.5 l=0.5
X2700 dvss.t1538 a_29702_24619# a_29802_24707# dvss.t1537 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X2701 por_ana_0.comparator_1.vm.t6 por_ana_0.comparator_1.ena_b avss.t253 avss.t252 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X2702 a_36962_32615# por_dig_0._035_ por_dig_0._036_.t1 dvdd.t1235 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X2703 dvdd.t1782 dvss.t2332 dvdd.t1781 dvdd.t1780 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X2704 dvss.t2029 por_dig_0.cnt_st\[2\] a_38926_33453# dvss.t2028 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2705 dvdd.t928 a_34010_31821# a_34116_31821# dvdd.t927 sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.5
X2706 a_19094_870# a_41694_492# dvss.t2026 sky130_fd_pr__res_xhigh_po_1p41 l=111
X2707 dvss.t310 a_38228_30163# a_38162_30189# dvss.t309 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X2708 a_36138_22973# a_36038_22885# dvss.t274 dvss.t273 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X2709 a_24212_13935# a_23834_6535# avss.t362 sky130_fd_pr__res_xhigh_po_1p41 l=35
X2710 a_30495_21859# a_30070_21903# dvss.t664 dvss.t663 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X2711 dvdd.t930 por_dig_0.cnt_por\[7\] por_dig_0._025_ dvdd.t929 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.165 ps=1.33 w=1 l=0.15
X2712 dvdd.t698 por_dig_0.por_unbuf.t20 por_ana_0.sky130_fd_sc_hd__inv_4_4.Y dvdd.t697 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2713 por_ana_0.ibias_gen_0.isrc_sel.t1 a_39457_24371# dvss.t633 dvss.t517 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.121875 ps=1.075 w=0.75 l=0.5
X2714 dvss.t1476 a_25478_24619# a_25578_24707# dvss.t1475 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X2715 por_ana_0.ibias_gen_0.vn0.t3 por_ana_0.ibias_gen_0.vn0.t2 por_ana_0.ibias_gen_0.ve.t3 avss.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X2716 por_ana_0.comparator_0.vnn.t4 por_ana_0.comparator_0.vpp.t58 avdd.t186 avdd.t182 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X2717 por_dig_0.osc_ena.t0 a_31413_29619# dvss.t2077 dvss.t2076 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X2718 dvdd.t91 a_33804_31251# por_dig_0._027_ dvdd.t90 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2719 a_30070_21903# a_29702_22885# dvss.t481 dvss.t480 sky130_fd_pr__nfet_01v8 ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X2720 a_36414_31277# a_35224_31277# a_36305_31277# dvss.t1285 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X2721 por_ana_0.comparator_0.vnn.t34 por_ana_0.comparator_0.vnn.t33 avdd.t355 avdd.t182 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X2722 dvdd.t1465 por_dig_0.clknet_0_osc_ck.t46 a_35583_34541# dvdd.t1464 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2723 avss.t397 por_ana_0.ibias_gen_0.vn1.t2 por_ana_0.ibias_gen_0.vn1.t3 avss.t396 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=8
X2724 a_39094_32909# por_dig_0._029_ dvdd.t1367 dvdd.t1366 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2725 dvss.t1702 dvdd.t1905 dvss.t1701 dvss.t1700 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X2726 avdd.t495 a_36831_21859# a_36138_22973# avdd.t494 sky130_fd_pr__pfet_g5v0d10v5 ad=0.2142 pd=1.99 as=0.2142 ps=1.99 w=0.42 l=1
X2727 avdd.t646 por_ana_0.comparator_1.vnn.t60 por_ana_0.comparator_1.vpp.t28 avdd.t392 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X2728 a_37430_30707# a_37212_31111# dvss.t1264 dvss.t1263 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X2729 por_dig_0._005_ a_35704_35124# dvss.t1445 dvss.t1444 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.11285 ps=1.045 w=0.65 l=0.15
X2730 dvss.t507 por_dig_0.clknet_1_0__leaf_osc_ck.t47 a_32188_30739# dvss.t506 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2731 dvss.t1573 por_dig_0.cnt_por\[2\] a_34633_36147# dvss.t1572 sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.10725 ps=0.98 w=0.65 l=0.15
X2732 dvdd.t1784 dvss.t2333 dvdd.t1783 dvdd.t1710 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X2733 dvss.t137 a_34387_32909# por_dig_0.clknet_0_osc_ck.t1 dvss.t136 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2734 a_33545_33287# a_32464_32915# a_33198_32883# dvdd.t400 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X2735 dvss.t1303 otrip[2].t3 a_34615_28013# dvss.t677 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X2736 avss.t388 por_ana_0.comparator_0.vn.t1 por_ana_0.comparator_0.vn.t2 avss.t45 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X2737 avdd.t265 a_24159_23593# a_23466_24707# avdd.t264 sky130_fd_pr__pfet_g5v0d10v5 ad=0.2142 pd=1.99 as=0.2142 ps=1.99 w=0.42 l=1
X2738 a_27690_24707# a_27590_24619# dvss.t1377 dvss.t1376 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X2739 dvdd.t1786 dvss.t2334 dvdd.t1785 dvdd.t1522 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X2740 a_37117_31099# por_dig_0._004_ dvss.t1196 dvss.t1195 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X2741 dcomp.t1 por_ana_0.sky130_fd_sc_hd__inv_4_3.Y dvss.t51 dvss.t50 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2742 dvdd.t73 por_dig_0.net4 por_dig_0._048_ dvdd.t72 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2743 por_ana_0.comparator_0.vinn.t12 avss.t48 por_ana_0.comparator_0.vinn.t12 avss.t49 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=0.6
X2744 a_37212_31111# a_36862_30739# a_37117_31099# dvdd.t1080 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X2745 dvdd.t1788 dvss.t2335 dvdd.t1787 dvdd.t1600 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X2746 a_25578_24707# a_25478_24619# dvss.t1474 dvss.t1473 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X2747 a_33374_31277# por_dig_0.net22.t23 por_dig_0._026_ dvss.t717 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2748 dvss.t1699 dvdd.t1906 dvss.t1698 dvss.t1697 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X2749 dvdd.t770 por_dig_0.net23.t22 por_dig_0._051_ dvdd.t769 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2750 a_31781_32187# por_dig_0.net28 dvdd.t1020 dvdd.t1019 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X2751 dvss.t360 a_25846_23637# a_26271_23593# dvss.t359 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X2752 dvdd.t1401 por_dig_0.cnt_por\[5\] por_dig_0._035_ dvdd.t1400 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.165 ps=1.33 w=1 l=0.15
X2753 a_33431_30733# a_32354_30739# a_33269_31111# dvdd.t1520 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X2754 a_36862_30739# a_36696_30739# dvss.t1260 dvss.t1259 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2755 por_ana_0.rstring_mux_0.otrip_decoded_avdd[4] a_26785_22637# avdd.t314 avdd.t313 sky130_fd_pr__pfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.24375 ps=1.825 w=1.5 l=0.5
X2756 por_ana_0.rstring_mux_0.vtrip_decoded_b_avdd[2] por_ana_0.rstring_mux_0.vtrip_decoded_avdd[2] avdd.t474 avdd.t473 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X2757 avdd.t647 por_ana_0.comparator_1.vnn.t61 por_ana_0.comparator_1.vpp.t29 avdd.t392 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X2758 dvdd.t639 a_33545_33287# a_33720_33213# dvdd.t638 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X2759 osc_ck.t0 por_ana_0.rc_osc_0.ena_b por_ana_0.rc_osc_0.vr dvdd.t823 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.1475 ps=1.295 w=1 l=0.18
X2760 dvss.t552 por_ana_0.dcomp3v3uv a_39887_23089# dvss.t551 sky130_fd_pr__nfet_g5v0d10v5 ad=0.178875 pd=1.26 as=0.1197 ps=1.41 w=0.42 l=0.5
X2761 por_dig_0.cnt_st\[3\] a_38228_30163# dvss.t308 dvss.t307 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X2762 dvss.t1278 por_ana_0.dcomp3v3 a_39888_24823# dvss.t1277 sky130_fd_pr__nfet_g5v0d10v5 ad=0.178875 pd=1.26 as=0.1197 ps=1.41 w=0.42 l=0.5
X2763 dvss.t2050 a_31814_24619# a_31914_24707# dvss.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X2764 por_dig_0.net14 a_35774_28673# dvss.t736 dvss.t735 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.122275 ps=1.08 w=0.65 l=0.15
X2765 a_34578_29645# por_dig_0._028_ a_34496_29645# dvdd.t70 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2766 dvss.t719 a_39328_34515# a_39070_34515# dvss.t718 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.5
X2767 a_36476_30163# por_dig_0.cnt_por\[10\] dvdd.t1230 dvdd.t1229 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2768 dvdd.t1791 dvss.t2336 dvdd.t1790 dvdd.t1789 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X2769 a_37580_34375# a_37230_34003# a_37485_34363# dvdd.t914 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X2770 dvdd.t153 a_34098_30707# por_dig_0.clknet_1_0__leaf_osc_ck.t18 dvdd.t152 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X2771 porb_h.t1 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.t37 avdd.t351 avdd.t350 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X2772 dvss.t1026 a_39888_23693# a_40247_23627# dvss.t1025 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.19875 ps=2.03 w=0.75 l=0.5
X2773 dvdd.t271 a_39162_33453# a_39268_33453# dvdd.t270 sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.5
X2774 a_38070_33287# a_36880_32915# a_37961_33287# dvss.t519 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X2775 a_38250_22973# a_38150_22885# dvss.t106 dvss.t105 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X2776 por_dig_0._049_ por_dig_0.cnt_por\[1\] a_35776_36967# dvdd.t1158 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X2777 a_33163_32365# por_dig_0.net24 dvss.t405 dvss.t404 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X2778 dvdd.t261 por_dig_0.cnt_por\[8\] por_dig_0._037_ dvdd.t260 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X2779 avss.t283 por_ana_0.comparator_0.n1.t18 por_ana_0.dcomp3v3uv avss.t282 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X2780 a_32607_21859# a_32182_21903# dvss.t1114 dvss.t1113 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X2781 dvss.t1375 a_27590_24619# a_27690_24707# dvss.t1374 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X2782 a_21188_13935# a_21566_6535# avss.t363 sky130_fd_pr__res_xhigh_po_1p41 l=35
X2783 a_28383_23593# a_27958_23637# dvss.t779 dvss.t778 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X2784 dvdd.t461 a_36756_35603# por_dig_0.cnt_por\[0\].t4 dvdd.t460 sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=2.61 as=0.135 ps=1.27 w=1 l=0.15
X2785 porb_h.t16 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.t38 avss.t209 avss.t208 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X2786 por_ana_0.comparator_0.vnn avss.t443 por_ana_0.comparator_0.vt.t20 por_ana_0.comparator_0.vt.t18 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=8
X2787 a_32182_21903# a_31814_22885# dvss.t2158 dvss.t2157 sky130_fd_pr__nfet_01v8 ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X2788 por_ana_0.comparator_0.vinn.t0 avdd.t15 por_ana_0.comparator_0.vinn.t0 avdd.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=0.6
X2789 dvdd.t1110 por_dig_0.cnt_st\[0\] por_dig_0._029_ dvdd.t1109 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2790 a_31849_31643# a_31412_31251# dvdd.t1341 dvdd.t1340 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X2791 a_17408_13935# a_17030_6535# avss.t364 sky130_fd_pr__res_xhigh_po_1p41 l=35
X2792 a_22047_21859# a_21622_21903# dvss.t1098 dvss.t1097 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X2793 dvdd.t784 a_34467_28557# a_34573_28557# dvdd.t783 sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X2794 a_33282_33453# por_dig_0._019_ dvss.t2174 dvss.t2173 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2795 por_dig_0._037_ por_dig_0.cnt_por\[9\] a_33550_32141# dvss.t2183 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X2796 a_34026_24707# a_33926_24619# dvss.t511 dvss.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X2797 a_35740_31277# a_35390_31277# a_35645_31277# dvdd.t801 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X2798 avdd.t498 a_38943_21859# a_38250_22973# avdd.t497 sky130_fd_pr__pfet_g5v0d10v5 ad=0.2142 pd=1.99 as=0.2142 ps=1.99 w=0.42 l=1
X2799 pwup_filt.t19 por_ana_0.sky130_fd_sc_hd__inv_4_0.Y dvdd.t201 dvdd.t200 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2800 dvss.t945 por_dig_0.net25 a_37842_34363# dvss.t944 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X2801 por_dig_0.net5.t1 a_32039_28013# dvdd.t1024 dvdd.t1023 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X2802 por_ana_0.rstring_mux_0.vtop.t2 por_ana_0.rstring_mux_0.ena_b avdd.t223 avdd.t222 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X2803 por_ana_0.comparator_0.vnn.t3 por_ana_0.comparator_0.vpp.t59 avdd.t185 avdd.t182 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X2804 avdd.t353 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.t39 porb_h.t0 avdd.t352 sky130_fd_pr__pfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X2805 a_18164_13935# a_18542_6535# avss.t243 sky130_fd_pr__res_xhigh_po_1p41 l=35
X2806 a_34750_28557# a_34573_28557# dvss.t747 dvss.t746 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X2807 por_dig_0.net23.t2 a_36564_32339# dvdd.t581 dvdd.t580 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2808 a_33686_34335# por_dig_0.net4 a_33600_34335# dvss.t84 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X2809 a_35921_35629# por_dig_0._005_ dvss.t674 dvss.t673 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X2810 a_31932_33595# por_dig_0.clknet_1_1__leaf_osc_ck.t48 dvdd.t1234 dvdd.t1233 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2811 dvdd.t1042 a_35100_32339# por_dig_0.net24 dvdd.t1041 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2812 por_ana_0.rstring_mux_0.otrip_decoded_b_avdd[4] por_ana_0.rstring_mux_0.otrip_decoded_avdd[4] avdd.t601 avdd.t600 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X2813 a_31650_33453# a_31615_33705# a_31412_33427# dvss.t833 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.1092 ps=1.36 w=0.42 l=0.15
X2814 dvdd.t1211 a_37777_31111# a_37952_31037# dvdd.t1210 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X2815 a_33474_36147# a_33256_36551# dvss.t1442 dvss.t1441 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X2816 dvdd.t428 por_dig_0.clknet_1_0__leaf_osc_ck.t48 a_34212_30189# dvdd.t427 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X2817 avdd.t418 por_ana_0.comparator_1.vpp.t62 por_ana_0.comparator_1.vnn.t16 avdd.t401 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X2818 a_36305_31277# a_35390_31277# a_35958_31519# dvss.t923 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X2819 dvdd.t1157 por_dig_0.cnt_por\[1\] a_34114_35879# dvdd.t1156 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2820 vin.t0 por_ana_0.rstring_mux_0.otrip_decoded_avdd[2] por_ana_0.rstring_mux_0.vtrip2.t0 avss.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X2821 dvss.t920 a_31592_30965# por_dig_0._038_ dvss.t919 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.17875 ps=1.85 w=0.65 l=0.15
X2822 por_ana_0.rstring_mux_0.otrip_decoded_avdd[6] a_28897_22637# avdd.t569 avdd.t565 sky130_fd_pr__pfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.24375 ps=1.825 w=1.5 l=0.5
X2823 por_dig_0.clknet_1_0__leaf_osc_ck.t0 a_34098_30707# dvss.t180 dvss.t179 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.05775 ps=0.695 w=0.42 l=0.15
X2824 dvdd.t1793 dvss.t2337 dvdd.t1792 dvdd.t1707 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X2825 avdd.t221 por_ana_0.rstring_mux_0.ena_b por_ana_0.rstring_mux_0.vtop.t1 avdd.t220 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X2826 avdd.t509 a_21354_22973# a_22561_22637# avdd.t309 sky130_fd_pr__pfet_g5v0d10v5 ad=0.24375 pd=1.825 as=0.3975 ps=3.53 w=1.5 l=0.5
X2827 por_dig_0.net32 a_34116_31821# dvdd.t667 dvdd.t666 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X2828 por_ana_0.rc_osc_0.m por_ana_0.rc_osc_0.n.t12 dvdd.t1361 dvdd.t1360 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2829 dvss.t510 a_33926_24619# a_34026_24707# dvss.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X2830 a_36380_33971# por_dig_0.net23.t23 dvdd.t772 dvdd.t771 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.1625 ps=1.325 w=1 l=0.15
X2831 por_dig_0.net9 por_dig_0.net3 dvss.t1355 dvss.t1354 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2832 por_ana_0.rc_osc_0.in dvss.t287 sky130_fd_pr__cap_mim_m3_2 l=30 w=30
X2833 a_39634_32615# por_dig_0.cnt_st\[0\] dvdd.t1108 dvdd.t1107 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.1475 ps=1.295 w=1 l=0.15
X2834 avdd.t14 avdd.t12 avdd.t14 avdd.t13 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=8
X2835 dvss.t1011 a_38250_24707# a_39457_24371# dvss.t517 sky130_fd_pr__nfet_g5v0d10v5 ad=0.121875 pd=1.075 as=0.19875 ps=2.03 w=0.75 l=0.5
X2836 por_ana_0.sky130_fd_sc_hvl__inv_4_0.A por_ana_0.sky130_fd_sc_hvl__inv_1_0.A avdd.t444 avdd.t443 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X2837 dvdd.t141 por_dig_0._031_ a_36382_31795# dvdd.t140 sky130_fd_pr__pfet_01v8_hvt ad=0.15 pd=1.3 as=0.1375 ps=1.275 w=1 l=0.15
X2838 dvdd.t1795 dvss.t2338 dvdd.t1794 dvdd.t1721 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X2839 dvss.t1536 a_29702_24619# a_29802_24707# dvss.t1535 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X2840 dvdd.t1174 por_dig_0.net8 a_32233_31643# dvdd.t1173 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1092 ps=1.36 w=0.42 l=0.15
X2841 avdd.t648 por_ana_0.comparator_1.vnn.t62 por_ana_0.comparator_1.vpp.t30 avdd.t392 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X2842 a_36234_35871# a_36016_35629# dvss.t942 dvss.t941 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X2843 avss.t350 por_ana_0.comparator_0.vm.t7 por_ana_0.comparator_0.n0.t3 avss.t100 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X2844 a_34294_21903# a_33926_22885# dvss.t606 dvss.t605 sky130_fd_pr__nfet_01v8 ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X2845 por_dig_0.cnt_por\[7\] a_32984_32339# dvss.t1236 dvss.t1235 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X2846 por_ana_0.comparator_0.vnn avss.t444 por_ana_0.comparator_0.vt.t19 por_ana_0.comparator_0.vt.t18 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=8
X2847 dvdd.t1798 dvss.t2339 dvdd.t1797 dvdd.t1796 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X2848 por_ana_0.ibias_gen_0.vp1.t11 por_ana_0.ibias_gen_0.vp1.t10 avdd.t622 avdd.t621 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X2849 a_34387_32909# osc_ck.t15 dvss.t893 dvss.t892 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2850 dvdd.t800 por_dig_0._038_ por_dig_0.net10 dvdd.t799 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.135 ps=1.27 w=1 l=0.15
X2851 por_dig_0.clknet_0_osc_ck.t0 a_34387_32909# dvss.t135 dvss.t134 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.05775 ps=0.695 w=0.42 l=0.15
X2852 avdd.t184 por_ana_0.comparator_0.vpp.t60 por_ana_0.comparator_0.vnn.t2 avdd.t180 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X2853 a_24159_21859# a_23734_21903# dvss.t1407 dvss.t1406 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X2854 por_ana_0.ibias_gen_0.ena_b.t2 por_ana_0.rstring_mux_0.ena.t13 avdd.t618 avdd.t617 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=1
X2855 a_36138_24707# a_36038_24619# dvss.t679 dvss.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X2856 dvss.t376 por_dig_0._022_ a_35040_34317# dvss.t100 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X2857 a_19094_3138# a_41694_3516# dvss.t1177 sky130_fd_pr__res_xhigh_po_1p41 l=111
X2858 a_34728_30189# a_34212_30189# a_34633_30189# dvss.t1279 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X2859 por_ana_0.comparator_0.n0.t2 por_ana_0.comparator_0.vm.t8 avss.t351 avss.t100 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X2860 dvdd.t273 por_ana_0.sky130_fd_sc_hd__inv_4_1.Y porb.t16 dvdd.t272 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2861 dvss.t1396 por_dig_0._016_ a_33465_35629# dvss.t1395 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X2862 dvdd.t1801 dvss.t2340 dvdd.t1800 dvdd.t1799 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X2863 avdd.t354 por_ana_0.comparator_0.vnn.t31 por_ana_0.comparator_0.vnn.t32 avdd.t180 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X2864 vin.t36 por_ana_0.rstring_mux_0.otrip_decoded_b_avdd[2] por_ana_0.rstring_mux_0.vtrip2.t6 avdd.t526 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X2865 a_35202_29877# a_35298_29619# dvdd.t326 dvdd.t325 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14075 ps=1.325 w=0.42 l=0.5
X2866 a_34633_30189# por_dig_0._014_ dvdd.t1486 dvdd.t1485 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X2867 a_36494_35091# a_36328_35091# dvdd.t870 dvdd.t869 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2868 por_dig_0._030_ a_38352_32365# dvdd.t627 dvdd.t626 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X2869 a_32828_35879# por_dig_0._052_ dvdd.t913 dvdd.t912 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X2870 por_ana_0.rstring_mux_0.vtrip_decoded_b_avdd[4] por_ana_0.rstring_mux_0.vtrip_decoded_avdd[4].t5 avss.t330 avss.t329 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X2871 dvdd.t139 por_dig_0._031_ por_dig_0._032_ dvdd.t138 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2872 a_15896_13935# a_15518_6535# avss.t244 sky130_fd_pr__res_xhigh_po_1p41 l=35
X2873 a_32906_36179# a_32740_36179# dvss.t446 dvss.t445 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2874 avdd.t11 avdd.t9 avdd.t10 avdd.t3 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=8
X2875 dvdd.t551 por_dig_0.cnt_por\[0\].t26 a_34762_36173# dvdd.t550 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X2876 avdd.t8 avdd.t6 avdd.t7 avdd.t3 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=8
X2877 por_ana_0.comparator_0.vn.t6 por_ana_0.comparator_0.ena_b.t5 por_ana_0.comparator_0.ibias.t3 avdd.t574 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X2878 dvdd.t1363 por_ana_0.rc_osc_0.n.t13 por_ana_0.rc_osc_0.m dvdd.t1362 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2879 por_dig_0.clknet_1_0__leaf_osc_ck.t17 a_34098_30707# dvdd.t151 dvdd.t150 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2880 por_dig_0.net1 a_31360_33997# dvdd.t1480 dvdd.t1479 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X2881 avdd.t597 a_23466_22973# a_24673_22637# avdd.t596 sky130_fd_pr__pfet_g5v0d10v5 ad=0.24375 pd=1.825 as=0.3975 ps=3.53 w=1.5 l=0.5
X2882 a_38576_13935# a_38198_6535# avss.t245 sky130_fd_pr__res_xhigh_po_1p41 l=35
X2883 dvdd.t1804 dvss.t2341 dvdd.t1803 dvdd.t1802 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X2884 a_38434_32365# por_dig_0.cnt_st\[1\] a_38352_32365# dvss.t597 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X2885 dcomp.t0 por_ana_0.sky130_fd_sc_hd__inv_4_3.Y dvss.t49 dvss.t48 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2886 a_35768_33690# a_35612_33595# a_35913_33819# dvdd.t1206 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.1155 ps=0.97 w=0.42 l=0.15
X2887 dvdd.t199 por_ana_0.sky130_fd_sc_hd__inv_4_0.Y pwup_filt.t18 dvdd.t198 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2888 por_ana_0.comparator_0.ena_b.t1 avss.t41 avss.t43 avss.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X2889 avdd.t297 a_21354_24707# a_22047_23593# avdd.t296 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.1365 ps=1.49 w=0.42 l=1
X2890 por_ana_0.sky130_fd_sc_hd__inv_4_1.Y por_ana_0.sky130_fd_sc_hd__inv_4_1.A dvss.t220 dvss.t219 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2891 por_ana_0.ibias_gen_0.vp0.t5 avss.t39 por_ana_0.ibias_gen_0.vn0.t16 avss.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X2892 dvss.t509 por_dig_0.clknet_1_0__leaf_osc_ck.t49 a_36696_30739# dvss.t508 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2893 dcomp.t16 por_ana_0.sky130_fd_sc_hd__inv_4_3.Y dvdd.t37 dvdd.t36 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2894 por_ana_0.comparator_0.vnn.t1 por_ana_0.comparator_0.vpp.t61 avdd.t183 avdd.t182 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X2895 por_ana_0.comparator_1.vnn.t41 vbg_1v2.t40 por_ana_0.comparator_1.vt.t40 por_ana_0.comparator_1.vt.t36 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X2896 a_33720_33213# por_dig_0.net24 dvdd.t333 dvdd.t332 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X2897 dvdd.t1236 por_dig_0.clknet_1_1__leaf_osc_ck.t49 a_36880_32915# dvdd.t1235 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X2898 por_ana_0.ibias_gen_0.vp1.t16 por_ana_0.ibias_gen_0.isrc_sel.t9 avdd.t585 avdd.t584 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=2
X2899 a_36406_21903# a_36038_22885# dvss.t272 dvss.t271 sky130_fd_pr__nfet_01v8 ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X2900 a_32906_35091# a_32740_35091# dvss.t1220 dvss.t1219 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2901 por_ana_0.sky130_fd_sc_hd__inv_4_1.A por_dig_0.por_unbuf.t21 dvdd.t700 dvdd.t699 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2902 dvdd.t1431 por_dig_0.net20.t9 por_dig_0._016_ dvdd.t1430 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2903 avdd.t219 por_ana_0.rstring_mux_0.ena_b por_ana_0.rstring_mux_0.vtop.t0 avdd.t218 sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=0.6
X2904 pwup_filt.t17 por_ana_0.sky130_fd_sc_hd__inv_4_0.Y dvdd.t197 dvdd.t196 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2905 a_37616_32141# por_dig_0._042_ dvss.t303 dvss.t302 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.08775 ps=0.92 w=0.65 l=0.15
X2906 a_26271_21859# a_25846_21903# dvss.t998 dvss.t997 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X2907 a_36749_35451# por_dig_0._006_ dvdd.t525 dvdd.t524 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X2908 a_38250_24707# a_38150_24619# dvss.t41 dvss.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X2909 por_ana_0.comparator_1.vnn.t40 vbg_1v2.t41 por_ana_0.comparator_1.vt.t39 por_ana_0.comparator_1.vt.t36 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X2910 dvss.t1696 dvdd.t1907 dvss.t1695 dvss.t1694 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X2911 dvdd.t454 a_39417_31795# por_dig_0.net4 dvdd.t453 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X2912 por_ana_0.rstring_mux_0.otrip_decoded_b_avdd[6] por_ana_0.rstring_mux_0.otrip_decoded_avdd[6] avss.t372 avss.t371 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X2913 por_dig_0._037_ por_dig_0.cnt_por\[10\] dvdd.t1228 dvdd.t1227 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2914 avss.t38 avss.t36 avss.t38 avss.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=8
X2915 por_dig_0.otrip_decoded[0].t0 a_38444_28013# dvss.t1975 dvss.t523 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X2916 por_dig_0._049_ por_dig_0.cnt_por\[0\].t27 a_35859_36717# dvss.t647 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.095875 ps=0.945 w=0.65 l=0.15
X2917 por_dig_0.clknet_1_0__leaf_osc_ck.t16 a_34098_30707# dvdd.t149 dvdd.t148 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2918 por_ana_0.comparator_1.vt.t55 por_ana_0.comparator_1.vn.t8 avss.t295 avss.t294 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X2919 dvdd.t1471 por_dig_0._020_ a_34024_33703# dvdd.t1470 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X2920 dvdd.t1806 dvss.t2342 dvdd.t1805 dvdd.t1628 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X2921 a_34594_32615# por_dig_0._026_ por_dig_0._013_ dvdd.t1329 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.165 ps=1.33 w=1 l=0.15
X2922 por_ana_0.comparator_0.n1.t3 por_ana_0.comparator_0.n0.t8 avss.t299 avss.t298 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.6
X2923 a_34040_13935# a_33662_6535# avss.t246 sky130_fd_pr__res_xhigh_po_1p41 l=35
X2924 a_37939_30733# a_36862_30739# a_37777_31111# dvdd.t1079 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X2925 dvdd.t794 a_38500_31251# a_38242_31251# dvdd.t793 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.5
X2926 avdd.t658 a_25595_33708# a_26288_32594# avdd.t657 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.1365 ps=1.49 w=0.42 l=1
X2927 por_ana_0.ibias_gen_0.isrc_sel_b.t1 avss.t34 por_ana_0.ibias_gen_0.ena_b.t1 avss.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X2928 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[1] a_31009_24371# avdd.t517 avdd.t419 sky130_fd_pr__pfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.24375 ps=1.825 w=1.5 l=0.5
X2929 a_34098_30707# por_dig_0.clknet_0_osc_ck.t47 dvss.t2141 dvss.t2140 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2930 por_ana_0.comparator_1.vpp.t1 por_ana_0.comparator_1.vpp.t0 avdd.t455 avdd.t395 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X2931 dvdd.t259 a_36382_31795# por_dig_0.net20.t1 dvdd.t258 sky130_fd_pr__pfet_01v8_hvt ad=0.3125 pd=1.625 as=0.26 ps=2.52 w=1 l=0.15
X2932 dvss.t1693 dvdd.t1908 dvss.t1692 dvss.t1691 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X2933 avdd.t181 por_ana_0.comparator_0.vpp.t62 por_ana_0.comparator_0.vnn.t0 avdd.t180 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X2934 dvss.t1506 a_36480_31251# a_36414_31277# dvss.t1505 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X2935 a_26288_32594# a_25863_32638# dvss.t532 dvss.t531 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X2936 dvss.t1690 dvdd.t1909 dvss.t1689 dvss.t1688 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X2937 dvss.t1980 a_35768_33690# a_35699_33819# dvss.t1979 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0999 ps=0.985 w=0.64 l=0.15
X2938 por_ana_0.comparator_1.vnn.t39 vbg_1v2.t42 por_ana_0.comparator_1.vt.t38 por_ana_0.comparator_1.vt.t36 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X2939 dvdd.t195 por_ana_0.sky130_fd_sc_hd__inv_4_0.Y pwup_filt.t16 dvdd.t194 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2940 dvdd.t1809 dvss.t2343 dvdd.t1808 dvdd.t1807 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X2941 dvss.t1226 a_21622_23637# a_22047_23593# dvss.t1225 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X2942 a_33088_32909# por_dig_0.net24 dvdd.t331 dvdd.t330 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X2943 por_dig_0.net33 a_39268_33453# dvss.t167 dvss.t166 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X2944 dvss.t1687 dvdd.t1910 dvss.t1686 dvss.t1685 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X2945 por_dig_0._033_ a_34672_35451# dvss.t1214 dvss.t1213 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.196275 ps=1.33 w=0.65 l=0.15
X2946 a_34672_35451# por_dig_0.cnt_por\[3\] dvdd.t379 dvdd.t378 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X2947 por_ana_0.comparator_1.vnn.t38 vbg_1v2.t43 por_ana_0.comparator_1.vt.t37 por_ana_0.comparator_1.vt.t36 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X2948 avdd.t562 a_25578_22973# a_26785_22637# avdd.t313 sky130_fd_pr__pfet_g5v0d10v5 ad=0.24375 pd=1.825 as=0.3975 ps=3.53 w=1.5 l=0.5
X2949 dvdd.t386 por_dig_0.cnt_por\[6\] a_34580_34110# dvdd.t385 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2950 dvss.t1684 dvdd.t1911 dvss.t1683 dvss.t1682 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X2951 por_dig_0.clknet_1_1__leaf_osc_ck.t0 a_35583_34541# dvss.t566 dvss.t565 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2952 avdd.t5 avdd.t2 avdd.t4 avdd.t3 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=8
X2953 a_35100_32339# por_dig_0.net27 dvdd.t1396 dvdd.t1395 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.165 ps=1.33 w=1 l=0.15
X2954 por_ana_0.dcomp3v3uv por_ana_0.comparator_0.n1.t19 avdd.t492 avdd.t491 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
R2 por_ana_0.comparator_0.vpp.t46 por_ana_0.comparator_0.vpp.n2 241.742
R3 por_ana_0.comparator_0.vpp.n2 por_ana_0.comparator_0.vpp.n9 204.284
R4 por_ana_0.comparator_0.vpp.n2 por_ana_0.comparator_0.vpp.n23 204.284
R5 por_ana_0.comparator_0.vpp.n2 por_ana_0.comparator_0.vpp.n22 204.284
R6 por_ana_0.comparator_0.vpp.n2 por_ana_0.comparator_0.vpp.n21 204.284
R7 por_ana_0.comparator_0.vpp.n2 por_ana_0.comparator_0.vpp.n20 204.284
R8 por_ana_0.comparator_0.vpp.n2 por_ana_0.comparator_0.vpp.n19 204.284
R9 por_ana_0.comparator_0.vpp.n2 por_ana_0.comparator_0.vpp.n18 204.284
R10 por_ana_0.comparator_0.vpp.n2 por_ana_0.comparator_0.vpp.n6 199.786
R11 por_ana_0.comparator_0.vpp.n2 por_ana_0.comparator_0.vpp.n5 199.65
R12 por_ana_0.comparator_0.vpp.n2 por_ana_0.comparator_0.vpp.n7 199.65
R13 por_ana_0.comparator_0.vpp.n2 por_ana_0.comparator_0.vpp.n8 199.65
R14 por_ana_0.comparator_0.vpp.n1 por_ana_0.comparator_0.vpp.n10 71.9371
R15 por_ana_0.comparator_0.vpp.n1 por_ana_0.comparator_0.vpp.n17 70.9612
R16 por_ana_0.comparator_0.vpp.n1 por_ana_0.comparator_0.vpp.n16 70.9612
R17 por_ana_0.comparator_0.vpp.n1 por_ana_0.comparator_0.vpp.n15 70.9612
R18 por_ana_0.comparator_0.vpp.n1 por_ana_0.comparator_0.vpp.n14 70.9612
R19 por_ana_0.comparator_0.vpp.n1 por_ana_0.comparator_0.vpp.n13 70.9612
R20 por_ana_0.comparator_0.vpp.n1 por_ana_0.comparator_0.vpp.n12 70.9612
R21 por_ana_0.comparator_0.vpp.n1 por_ana_0.comparator_0.vpp.n11 70.9612
R22 por_ana_0.comparator_0.vpp.n6 por_ana_0.comparator_0.vpp.t15 27.6955
R23 por_ana_0.comparator_0.vpp.n6 por_ana_0.comparator_0.vpp.t13 27.6955
R24 por_ana_0.comparator_0.vpp.n5 por_ana_0.comparator_0.vpp.t11 27.6955
R25 por_ana_0.comparator_0.vpp.n5 por_ana_0.comparator_0.vpp.t5 27.6955
R26 por_ana_0.comparator_0.vpp.n7 por_ana_0.comparator_0.vpp.t9 27.6955
R27 por_ana_0.comparator_0.vpp.n7 por_ana_0.comparator_0.vpp.t3 27.6955
R28 por_ana_0.comparator_0.vpp.n8 por_ana_0.comparator_0.vpp.t7 27.6955
R29 por_ana_0.comparator_0.vpp.n8 por_ana_0.comparator_0.vpp.t1 27.6955
R30 por_ana_0.comparator_0.vpp.n9 por_ana_0.comparator_0.vpp.t32 27.6955
R31 por_ana_0.comparator_0.vpp.n9 por_ana_0.comparator_0.vpp.t38 27.6955
R32 por_ana_0.comparator_0.vpp.n23 por_ana_0.comparator_0.vpp.t34 27.6955
R33 por_ana_0.comparator_0.vpp.n23 por_ana_0.comparator_0.vpp.t40 27.6955
R34 por_ana_0.comparator_0.vpp.n22 por_ana_0.comparator_0.vpp.t33 27.6955
R35 por_ana_0.comparator_0.vpp.n22 por_ana_0.comparator_0.vpp.t39 27.6955
R36 por_ana_0.comparator_0.vpp.n21 por_ana_0.comparator_0.vpp.t42 27.6955
R37 por_ana_0.comparator_0.vpp.n21 por_ana_0.comparator_0.vpp.t45 27.6955
R38 por_ana_0.comparator_0.vpp.n20 por_ana_0.comparator_0.vpp.t37 27.6955
R39 por_ana_0.comparator_0.vpp.n20 por_ana_0.comparator_0.vpp.t41 27.6955
R40 por_ana_0.comparator_0.vpp.n19 por_ana_0.comparator_0.vpp.t43 27.6955
R41 por_ana_0.comparator_0.vpp.n19 por_ana_0.comparator_0.vpp.t35 27.6955
R42 por_ana_0.comparator_0.vpp.n18 por_ana_0.comparator_0.vpp.t44 27.6955
R43 por_ana_0.comparator_0.vpp.n18 por_ana_0.comparator_0.vpp.t36 27.6955
R44 por_ana_0.comparator_0.vpp.n1 por_ana_0.comparator_0.vpp.t57 23.5879
R45 por_ana_0.comparator_0.vpp.n2 por_ana_0.comparator_0.vpp.n1 18.1658
R46 por_ana_0.comparator_0.vpp.n1 por_ana_0.comparator_0.vpp.n0 18.106
R47 por_ana_0.comparator_0.vpp.n1 por_ana_0.comparator_0.vpp.n3 16.9748
R48 por_ana_0.comparator_0.vpp.n17 por_ana_0.comparator_0.vpp.t19 16.5305
R49 por_ana_0.comparator_0.vpp.n17 por_ana_0.comparator_0.vpp.t16 16.5305
R50 por_ana_0.comparator_0.vpp.n16 por_ana_0.comparator_0.vpp.t29 16.5305
R51 por_ana_0.comparator_0.vpp.n16 por_ana_0.comparator_0.vpp.t26 16.5305
R52 por_ana_0.comparator_0.vpp.n15 por_ana_0.comparator_0.vpp.t24 16.5305
R53 por_ana_0.comparator_0.vpp.n15 por_ana_0.comparator_0.vpp.t22 16.5305
R54 por_ana_0.comparator_0.vpp.n14 por_ana_0.comparator_0.vpp.t20 16.5305
R55 por_ana_0.comparator_0.vpp.n14 por_ana_0.comparator_0.vpp.t17 16.5305
R56 por_ana_0.comparator_0.vpp.n13 por_ana_0.comparator_0.vpp.t30 16.5305
R57 por_ana_0.comparator_0.vpp.n13 por_ana_0.comparator_0.vpp.t27 16.5305
R58 por_ana_0.comparator_0.vpp.n12 por_ana_0.comparator_0.vpp.t21 16.5305
R59 por_ana_0.comparator_0.vpp.n12 por_ana_0.comparator_0.vpp.t18 16.5305
R60 por_ana_0.comparator_0.vpp.n11 por_ana_0.comparator_0.vpp.t31 16.5305
R61 por_ana_0.comparator_0.vpp.n11 por_ana_0.comparator_0.vpp.t28 16.5305
R62 por_ana_0.comparator_0.vpp.n10 por_ana_0.comparator_0.vpp.t25 16.5305
R63 por_ana_0.comparator_0.vpp.n10 por_ana_0.comparator_0.vpp.t23 16.5305
R64 por_ana_0.comparator_0.vpp.n0 por_ana_0.comparator_0.vpp.t60 16.3148
R65 por_ana_0.comparator_0.vpp.n0 por_ana_0.comparator_0.vpp.t48 16.3148
R66 por_ana_0.comparator_0.vpp.n4 por_ana_0.comparator_0.vpp.t62 16.3148
R67 por_ana_0.comparator_0.vpp.n0 por_ana_0.comparator_0.vpp.t53 16.3148
R68 por_ana_0.comparator_0.vpp.n0 por_ana_0.comparator_0.vpp.t49 16.3148
R69 por_ana_0.comparator_0.vpp.n1 por_ana_0.comparator_0.vpp.t54 16.3148
R70 por_ana_0.comparator_0.vpp.n1 por_ana_0.comparator_0.vpp.t56 16.3148
R71 por_ana_0.comparator_0.vpp.n3 por_ana_0.comparator_0.vpp.t51 16.3148
R72 por_ana_0.comparator_0.vpp.n2 por_ana_0.comparator_0.vpp.t0 14.2251
R73 por_ana_0.comparator_0.vpp.n2 por_ana_0.comparator_0.vpp.t6 14.2251
R74 por_ana_0.comparator_0.vpp.n2 por_ana_0.comparator_0.vpp.t2 14.2251
R75 por_ana_0.comparator_0.vpp.n2 por_ana_0.comparator_0.vpp.t8 14.2251
R76 por_ana_0.comparator_0.vpp.n2 por_ana_0.comparator_0.vpp.t4 14.2251
R77 por_ana_0.comparator_0.vpp.n2 por_ana_0.comparator_0.vpp.t10 14.2251
R78 por_ana_0.comparator_0.vpp.n2 por_ana_0.comparator_0.vpp.t14 14.2251
R79 por_ana_0.comparator_0.vpp.n2 por_ana_0.comparator_0.vpp.t12 14.2251
R80 por_ana_0.comparator_0.vpp.n0 por_ana_0.comparator_0.vpp.n4 14.2134
R81 por_ana_0.comparator_0.vpp.n0 por_ana_0.comparator_0.vpp.t58 12.0866
R82 por_ana_0.comparator_0.vpp.n0 por_ana_0.comparator_0.vpp.t61 12.0866
R83 por_ana_0.comparator_0.vpp.n4 por_ana_0.comparator_0.vpp.t59 12.0866
R84 por_ana_0.comparator_0.vpp.n0 por_ana_0.comparator_0.vpp.t50 12.0866
R85 por_ana_0.comparator_0.vpp.n0 por_ana_0.comparator_0.vpp.t47 12.0866
R86 por_ana_0.comparator_0.vpp.n1 por_ana_0.comparator_0.vpp.t55 12.0866
R87 por_ana_0.comparator_0.vpp.n3 por_ana_0.comparator_0.vpp.t52 12.0866
R88 avdd.n1720 avdd.n954 99969.2
R89 avdd.n1720 avdd.n1719 83663.1
R90 avdd.n1704 avdd.n955 66867
R91 avdd.n1705 avdd.n956 60783.5
R92 avdd.n1704 avdd.n1703 60384.8
R93 avdd.n971 avdd.n954 58787
R94 avdd.n1717 avdd.n956 52810.3
R95 avdd.n1718 avdd.n955 50831
R96 avdd.n1721 avdd.n952 49200
R97 avdd.n1703 avdd.n1702 47131.3
R98 avdd.n1721 avdd.n953 41239.5
R99 avdd.n1705 avdd.n961 29875.1
R100 avdd.n972 avdd.n952 29132.4
R101 avdd.n1719 avdd.n1718 27601.7
R102 avdd.n971 avdd.n962 27058.6
R103 avdd.n470 avdd.n343 25108.6
R104 avdd.n468 avdd.n343 25108.6
R105 avdd.n894 avdd.n591 25108.6
R106 avdd.n892 avdd.n591 25108.6
R107 avdd.n470 avdd.n469 25105.2
R108 avdd.n469 avdd.n468 25105.2
R109 avdd.n894 avdd.n893 25105.2
R110 avdd.n893 avdd.n892 25105.2
R111 avdd.n1701 avdd.n961 22957.3
R112 avdd.n1702 avdd.n962 17438.8
R113 avdd.n1773 avdd.n1766 15077.5
R114 avdd.n1773 avdd.n1767 15077.5
R115 avdd.n1810 avdd.n1767 15077.5
R116 avdd.n1810 avdd.n1766 15077.5
R117 avdd.n1717 avdd.n953 13877.8
R118 avdd.n972 avdd.n963 13642.7
R119 avdd.n471 avdd.n341 12653.5
R120 avdd.n467 avdd.n341 12653.5
R121 avdd.n895 avdd.n589 12653.5
R122 avdd.n891 avdd.n589 12653.5
R123 avdd.n471 avdd.n342 12651.9
R124 avdd.n467 avdd.n342 12651.9
R125 avdd.n895 avdd.n590 12651.9
R126 avdd.n891 avdd.n590 12651.9
R127 avdd.n491 avdd.n288 11582.8
R128 avdd.n451 avdd.n288 11582.8
R129 avdd.n915 avdd.n536 11582.8
R130 avdd.n875 avdd.n536 11582.8
R131 avdd.n493 avdd.n285 10507.7
R132 avdd.n453 avdd.n285 10507.7
R133 avdd.n917 avdd.n533 10507.7
R134 avdd.n877 avdd.n533 10507.7
R135 avdd.n485 avdd.n305 10039.9
R136 avdd.n485 avdd.n284 10039.9
R137 avdd.n487 avdd.n304 10039.9
R138 avdd.n487 avdd.n289 10039.9
R139 avdd.n909 avdd.n553 10039.9
R140 avdd.n909 avdd.n532 10039.9
R141 avdd.n911 avdd.n552 10039.9
R142 avdd.n911 avdd.n537 10039.9
R143 avdd.n1874 avdd.n18 9739.14
R144 avdd.n1874 avdd.n19 9739.14
R145 avdd.n1873 avdd.n19 9739.14
R146 avdd.n1873 avdd.n18 9739.14
R147 avdd.n1701 avdd.n963 8461.62
R148 avdd.n1707 avdd.n957 8070.02
R149 avdd.n1706 avdd.n960 6943.25
R150 avdd.n970 avdd.n969 6761.04
R151 avdd.n1716 avdd.n957 6168.09
R152 avdd.n1699 avdd.n965 5303.72
R153 avdd.n1712 avdd.n1711 4892.23
R154 avdd.n1723 avdd.n950 4681.79
R155 avdd.n967 avdd.n950 4335.44
R156 avdd.n1858 avdd.n1857 4316.28
R157 avdd.n1860 avdd.n1857 4316.28
R158 avdd.n1858 avdd.n1854 4316.28
R159 avdd.n1860 avdd.n1854 4316.28
R160 avdd.n1715 avdd.n958 3225.22
R161 avdd.n974 avdd.n973 3163.48
R162 avdd.n1825 avdd.n1738 3160.55
R163 avdd.n1826 avdd.n1738 3160.55
R164 avdd.n472 avdd.n340 2933.46
R165 avdd.n896 avdd.n588 2933.46
R166 avdd.n466 avdd.n344 2922.54
R167 avdd.n890 avdd.n592 2922.54
R168 avdd.n1809 avdd.n1768 2890.84
R169 avdd.n1774 avdd.n1768 2890.84
R170 avdd.n465 avdd.n345 2865.69
R171 avdd.n889 avdd.n593 2865.69
R172 avdd.n1775 avdd.n1769 2860.42
R173 avdd.n1808 avdd.n1769 2860.42
R174 avdd.n473 avdd.n339 2841.22
R175 avdd.n897 avdd.n587 2841.22
R176 avdd.n449 avdd.n304 2620.03
R177 avdd.n449 avdd.n305 2620.03
R178 avdd.n289 avdd.n286 2620.03
R179 avdd.n286 avdd.n284 2620.03
R180 avdd.n873 avdd.n552 2620.03
R181 avdd.n873 avdd.n553 2620.03
R182 avdd.n537 avdd.n534 2620.03
R183 avdd.n534 avdd.n532 2620.03
R184 avdd.n1819 avdd.n1745 2513.9
R185 avdd.n1819 avdd.n1737 2513.9
R186 avdd.n1820 avdd.n1742 2513.9
R187 avdd.n1820 avdd.n1739 2513.9
R188 avdd.n1711 avdd.n951 2495.62
R189 avdd.n447 avdd.n362 2480.48
R190 avdd.n447 avdd.n363 2480.48
R191 avdd.n362 avdd.n361 2480.48
R192 avdd.n363 avdd.n361 2480.48
R193 avdd.n871 avdd.n610 2480.48
R194 avdd.n871 avdd.n611 2480.48
R195 avdd.n610 avdd.n609 2480.48
R196 avdd.n611 avdd.n609 2480.48
R197 avdd.n1723 avdd.n1722 2412.42
R198 avdd.n1814 avdd.n1762 2346.83
R199 avdd.n1813 avdd.n1762 2346.83
R200 avdd.n450 avdd.n290 2223.06
R201 avdd.n490 avdd.n290 2223.06
R202 avdd.n874 avdd.n538 2223.06
R203 avdd.n914 avdd.n538 2223.06
R204 avdd.n1722 avdd.n951 2115.76
R205 avdd.n298 avdd.n297 2059.86
R206 avdd.n297 avdd.n296 2059.86
R207 avdd.n296 avdd.n293 2059.86
R208 avdd.n298 avdd.n293 2059.86
R209 avdd.n546 avdd.n545 2059.86
R210 avdd.n545 avdd.n544 2059.86
R211 avdd.n544 avdd.n541 2059.86
R212 avdd.n546 avdd.n541 2059.86
R213 avdd.n494 avdd.n283 2000.19
R214 avdd.n454 avdd.n283 2000.19
R215 avdd.n918 avdd.n531 2000.19
R216 avdd.n878 avdd.n531 2000.19
R217 avdd.n1700 avdd.n964 1971.95
R218 avdd.n488 avdd.n302 1923.01
R219 avdd.n489 avdd.n488 1923.01
R220 avdd.n912 avdd.n550 1923.01
R221 avdd.n913 avdd.n912 1923.01
R222 avdd.n1826 avdd.n1737 1837.76
R223 avdd.n1825 avdd.n1739 1837.76
R224 avdd.n20 avdd.n16 1616.56
R225 avdd.n21 avdd.n17 1616.56
R226 avdd.n1871 avdd.n21 1616.56
R227 avdd.n1876 avdd.n16 1615.06
R228 avdd.n491 avdd.n289 1542.93
R229 avdd.n451 avdd.n304 1542.93
R230 avdd.n915 avdd.n537 1542.93
R231 avdd.n875 avdd.n552 1542.93
R232 avdd.n1764 avdd.n1742 1322.79
R233 avdd.n1764 avdd.n1745 1322.79
R234 avdd.n1743 avdd.n1739 1322.79
R235 avdd.n1743 avdd.n1737 1322.79
R236 avdd.n484 avdd.n306 1237.08
R237 avdd.n484 avdd.n281 1237.08
R238 avdd.n908 avdd.n554 1237.08
R239 avdd.n908 avdd.n529 1237.08
R240 avdd.n1814 avdd.n1745 1024.03
R241 avdd.n1813 avdd.n1742 1024.03
R242 avdd.n1862 avdd.n1861 831.247
R243 avdd.n1862 avdd.n1853 831.247
R244 avdd.n982 avdd.t312 692.692
R245 avdd.n1355 avdd.t273 692.692
R246 avdd avdd.t472 688.231
R247 avdd avdd.t290 688.231
R248 avdd.n1856 avdd.n1855 682.918
R249 avdd.n1856 avdd.n1836 682.918
R250 avdd.n1196 avdd.t297 648.668
R251 avdd.n1211 avdd.t513 648.668
R252 avdd.n1226 avdd.t301 648.668
R253 avdd.n1241 avdd.t316 648.668
R254 avdd.n1256 avdd.t422 648.668
R255 avdd.n1271 avdd.t589 648.668
R256 avdd.n1286 avdd.t289 648.668
R257 avdd.n1301 avdd.t308 648.668
R258 avdd.n1316 avdd.t442 648.668
R259 avdd.n1533 avdd.t511 648.668
R260 avdd.n1548 avdd.t599 648.668
R261 avdd.n1563 avdd.t564 648.668
R262 avdd.n1578 avdd.t568 648.668
R263 avdd.n1593 avdd.t283 648.668
R264 avdd.n1608 avdd.t257 648.668
R265 avdd.n1623 avdd.t267 648.668
R266 avdd.n1638 avdd.t209 648.668
R267 avdd.n1653 avdd.t251 648.668
R268 avdd.n1191 avdd.t658 648.668
R269 avdd.n247 avdd.n31 624.808
R270 avdd.n245 avdd.n32 624.808
R271 avdd.n234 avdd.n233 624.808
R272 avdd.n222 avdd.n51 624.808
R273 avdd.n220 avdd.n52 624.808
R274 avdd.n209 avdd.n208 624.808
R275 avdd.n197 avdd.n71 624.808
R276 avdd.n195 avdd.n72 624.808
R277 avdd.n184 avdd.n183 624.808
R278 avdd.n172 avdd.n91 624.808
R279 avdd.n170 avdd.n92 624.808
R280 avdd.n159 avdd.n158 624.808
R281 avdd.n147 avdd.n111 624.808
R282 avdd.n145 avdd.n112 624.808
R283 avdd.n134 avdd.n133 624.808
R284 avdd.n456 avdd.n306 612.894
R285 avdd.n496 avdd.n281 612.894
R286 avdd.n880 avdd.n554 612.894
R287 avdd.n920 avdd.n529 612.894
R288 avdd.n1824 avdd.n1735 609.883
R289 avdd.n1828 avdd.n1827 555.672
R290 avdd.t378 avdd.t384 511.356
R291 avdd.t24 avdd.t380 511.356
R292 avdd.t550 avdd.t24 511.356
R293 avdd.t548 avdd.t550 511.356
R294 avdd.t115 avdd.t548 511.356
R295 avdd.t552 avdd.t115 511.356
R296 avdd.t554 avdd.t552 511.356
R297 avdd.t44 avdd.t554 511.356
R298 avdd.n455 avdd.n360 506.353
R299 avdd.n879 avdd.n608 506.353
R300 avdd.n6 avdd.t615 499.882
R301 avdd.t520 avdd.t524 484.288
R302 avdd.t574 avdd.t522 484.288
R303 avdd.t605 avdd.t609 484.288
R304 avdd.t460 avdd.t607 484.288
R305 avdd.n1818 avdd.n1816 481.507
R306 avdd.n1821 avdd.n1741 481.507
R307 avdd.n367 avdd.n366 479.625
R308 avdd.n366 avdd.n365 479.625
R309 avdd.n615 avdd.n614 479.625
R310 avdd.n614 avdd.n613 479.625
R311 avdd.t384 avdd.t386 475.098
R312 avdd.n493 avdd.n284 467.793
R313 avdd.n453 avdd.n305 467.793
R314 avdd.n917 avdd.n532 467.793
R315 avdd.n877 avdd.n553 467.793
R316 avdd.n1812 avdd.n1761 454.024
R317 avdd.n296 avdd.t574 437.699
R318 avdd.n544 avdd.t460 437.699
R319 avdd.n446 avdd.n364 437.082
R320 avdd.n446 avdd.n445 437.082
R321 avdd.n870 avdd.n612 437.082
R322 avdd.n870 avdd.n869 437.082
R323 avdd.n1815 avdd.n1761 423.818
R324 avdd.n299 avdd.n292 399.06
R325 avdd.n295 avdd.n292 399.06
R326 avdd.n547 avdd.n540 399.06
R327 avdd.n543 avdd.n540 399.06
R328 avdd.n1749 avdd.t175 397.264
R329 avdd.n1750 avdd.t119 397.135
R330 avdd.n1751 avdd.t107 397.135
R331 avdd.n15 avdd.t52 388.149
R332 avdd.n258 avdd.t98 388.149
R333 avdd.n259 avdd.t30 388.149
R334 avdd.n260 avdd.t117 388.149
R335 avdd.n261 avdd.t163 388.149
R336 avdd.n262 avdd.t66 388.149
R337 avdd.n263 avdd.t140 388.149
R338 avdd.n264 avdd.t37 388.149
R339 avdd.n266 avdd.t105 388.149
R340 avdd.n267 avdd.t156 388.149
R341 avdd.n268 avdd.t168 388.149
R342 avdd.n269 avdd.t72 388.149
R343 avdd.n270 avdd.t15 388.149
R344 avdd.n271 avdd.t39 388.149
R345 avdd.n272 avdd.t170 388.149
R346 avdd.n1155 avdd.t462 372.885
R347 avdd.n1134 avdd.t265 372.885
R348 avdd.n1113 avdd.t213 372.885
R349 avdd.n1092 avdd.t321 372.885
R350 avdd.n1071 avdd.t476 372.885
R351 avdd.n1050 avdd.t271 372.885
R352 avdd.n1029 avdd.t506 372.885
R353 avdd.n1008 avdd.t432 372.885
R354 avdd.n990 avdd.t656 372.885
R355 avdd.n1528 avdd.t428 372.885
R356 avdd.n1507 avdd.t305 372.885
R357 avdd.n1486 avdd.t438 372.885
R358 avdd.n1465 avdd.t652 372.885
R359 avdd.n1444 avdd.t457 372.885
R360 avdd.n1423 avdd.t263 372.885
R361 avdd.n1402 avdd.t516 372.885
R362 avdd.n1381 avdd.t495 372.885
R363 avdd.n1363 avdd.t498 372.885
R364 avdd.n1187 avdd.t217 372.885
R365 avdd.t619 avdd.n23 354.904
R366 avdd.n1827 avdd.n1736 352
R367 avdd.n1824 avdd.n1823 352
R368 avdd.n1773 avdd.t44 345.817
R369 avdd.n298 avdd.t520 343.495
R370 avdd.n546 avdd.t605 343.495
R371 avdd.n1817 avdd.n1736 325.647
R372 avdd.n1823 avdd.n1822 325.647
R373 avdd.n668 avdd.n667 325.039
R374 avdd.n362 avdd.t481 323.445
R375 avdd.n363 avdd.t499 323.445
R376 avdd.n610 avdd.t540 323.445
R377 avdd.n611 avdd.t544 323.445
R378 avdd.n132 avdd.n117 321.882
R379 avdd.n137 avdd.n136 321.882
R380 avdd.n136 avdd.n116 321.882
R381 avdd.n148 avdd.n108 321.882
R382 avdd.n144 avdd.n108 321.882
R383 avdd.n157 avdd.n97 321.882
R384 avdd.n110 avdd.n97 321.882
R385 avdd.n162 avdd.n161 321.882
R386 avdd.n161 avdd.n96 321.882
R387 avdd.n173 avdd.n88 321.882
R388 avdd.n169 avdd.n88 321.882
R389 avdd.n182 avdd.n77 321.882
R390 avdd.n90 avdd.n77 321.882
R391 avdd.n187 avdd.n186 321.882
R392 avdd.n186 avdd.n76 321.882
R393 avdd.n198 avdd.n68 321.882
R394 avdd.n194 avdd.n68 321.882
R395 avdd.n207 avdd.n57 321.882
R396 avdd.n70 avdd.n57 321.882
R397 avdd.n212 avdd.n211 321.882
R398 avdd.n211 avdd.n56 321.882
R399 avdd.n223 avdd.n48 321.882
R400 avdd.n219 avdd.n48 321.882
R401 avdd.n232 avdd.n37 321.882
R402 avdd.n50 avdd.n37 321.882
R403 avdd.n237 avdd.n236 321.882
R404 avdd.n236 avdd.n36 321.882
R405 avdd.n248 avdd.n29 321.882
R406 avdd.n244 avdd.n29 321.882
R407 avdd.n24 avdd.n23 321.882
R408 avdd.n25 avdd.n24 321.882
R409 avdd.n5 avdd.n4 321.882
R410 avdd.n1139 avdd.n1138 321.882
R411 avdd.n1149 avdd.n1148 321.882
R412 avdd.n1146 avdd.n1145 321.882
R413 avdd.n1118 avdd.n1117 321.882
R414 avdd.n1128 avdd.n1127 321.882
R415 avdd.n1125 avdd.n1124 321.882
R416 avdd.n1097 avdd.n1096 321.882
R417 avdd.n1107 avdd.n1106 321.882
R418 avdd.n1104 avdd.n1103 321.882
R419 avdd.n1076 avdd.n1075 321.882
R420 avdd.n1086 avdd.n1085 321.882
R421 avdd.n1083 avdd.n1082 321.882
R422 avdd.n1055 avdd.n1054 321.882
R423 avdd.n1065 avdd.n1064 321.882
R424 avdd.n1062 avdd.n1061 321.882
R425 avdd.n1034 avdd.n1033 321.882
R426 avdd.n1044 avdd.n1043 321.882
R427 avdd.n1041 avdd.n1040 321.882
R428 avdd.n1013 avdd.n1012 321.882
R429 avdd.n1023 avdd.n1022 321.882
R430 avdd.n1020 avdd.n1019 321.882
R431 avdd.n992 avdd.n991 321.882
R432 avdd.n1002 avdd.n1001 321.882
R433 avdd.n999 avdd.n998 321.882
R434 avdd.n980 avdd.n979 321.882
R435 avdd.n1321 avdd.n980 321.882
R436 avdd.n1321 avdd.n986 321.882
R437 avdd.n987 avdd.n986 321.882
R438 avdd.n1325 avdd.n987 321.882
R439 avdd.n1325 avdd.n1319 321.882
R440 avdd.n1329 avdd.n1319 321.882
R441 avdd.n1512 avdd.n1511 321.882
R442 avdd.n1522 avdd.n1521 321.882
R443 avdd.n1519 avdd.n1518 321.882
R444 avdd.n1491 avdd.n1490 321.882
R445 avdd.n1501 avdd.n1500 321.882
R446 avdd.n1498 avdd.n1497 321.882
R447 avdd.n1470 avdd.n1469 321.882
R448 avdd.n1480 avdd.n1479 321.882
R449 avdd.n1477 avdd.n1476 321.882
R450 avdd.n1449 avdd.n1448 321.882
R451 avdd.n1459 avdd.n1458 321.882
R452 avdd.n1456 avdd.n1455 321.882
R453 avdd.n1428 avdd.n1427 321.882
R454 avdd.n1438 avdd.n1437 321.882
R455 avdd.n1435 avdd.n1434 321.882
R456 avdd.n1407 avdd.n1406 321.882
R457 avdd.n1417 avdd.n1416 321.882
R458 avdd.n1414 avdd.n1413 321.882
R459 avdd.n1386 avdd.n1385 321.882
R460 avdd.n1396 avdd.n1395 321.882
R461 avdd.n1393 avdd.n1392 321.882
R462 avdd.n1365 avdd.n1364 321.882
R463 avdd.n1375 avdd.n1374 321.882
R464 avdd.n1372 avdd.n1371 321.882
R465 avdd.n1353 avdd.n1352 321.882
R466 avdd.n1658 avdd.n1359 321.882
R467 avdd.n1360 avdd.n1359 321.882
R468 avdd.n1662 avdd.n1360 321.882
R469 avdd.n1662 avdd.n1656 321.882
R470 avdd.n1666 avdd.n1656 321.882
R471 avdd.n1180 avdd.n1164 321.882
R472 avdd.n1170 avdd.n1169 321.882
R473 avdd.n1182 avdd.n1161 321.882
R474 avdd.n666 avdd.n663 321.882
R475 avdd.n672 avdd.n663 321.882
R476 avdd.n672 avdd.n661 321.882
R477 avdd.n677 avdd.n661 321.882
R478 avdd.n677 avdd.n657 321.882
R479 avdd.n683 avdd.n657 321.882
R480 avdd.n683 avdd.n656 321.882
R481 avdd.n687 avdd.n656 321.882
R482 avdd.n687 avdd.n652 321.882
R483 avdd.n693 avdd.n652 321.882
R484 avdd.n693 avdd.n650 321.882
R485 avdd.n698 avdd.n650 321.882
R486 avdd.n698 avdd.n646 321.882
R487 avdd.n704 avdd.n646 321.882
R488 avdd.n704 avdd.n645 321.882
R489 avdd.n708 avdd.n645 321.882
R490 avdd.n708 avdd.n641 321.882
R491 avdd.n714 avdd.n641 321.882
R492 avdd.n714 avdd.n639 321.882
R493 avdd.n719 avdd.n639 321.882
R494 avdd.n719 avdd.n635 321.882
R495 avdd.n725 avdd.n635 321.882
R496 avdd.n725 avdd.n634 321.882
R497 avdd.n730 avdd.n634 321.882
R498 avdd.n730 avdd.n630 321.882
R499 avdd.n736 avdd.n630 321.882
R500 avdd.n736 avdd.n629 321.882
R501 avdd.n741 avdd.n629 321.882
R502 avdd.n741 avdd.n624 321.882
R503 avdd.n768 avdd.n624 321.882
R504 avdd.n768 avdd.n622 321.882
R505 avdd.n772 avdd.n622 321.882
R506 avdd.n773 avdd.n772 321.882
R507 avdd.n773 avdd.n618 321.882
R508 avdd.n619 avdd.n618 321.882
R509 avdd.n621 avdd.n619 321.882
R510 avdd.n125 avdd.n124 318.757
R511 avdd.n778 avdd.n777 318.757
R512 avdd.n1658 avdd.n1353 318.529
R513 avdd.t13 avdd.t180 310.303
R514 avdd.t180 avdd.t182 310.303
R515 avdd.t195 avdd.t191 310.303
R516 avdd.t191 avdd.t3 310.303
R517 avdd.t33 avdd.t401 310.303
R518 avdd.t401 avdd.t403 310.303
R519 avdd.t392 avdd.t395 310.303
R520 avdd.t395 avdd.t27 310.303
R521 avdd.n450 avdd.n302 300.048
R522 avdd.n490 avdd.n489 300.048
R523 avdd.n300 avdd.n291 300.048
R524 avdd.n294 avdd.n291 300.048
R525 avdd.n874 avdd.n550 300.048
R526 avdd.n914 avdd.n913 300.048
R527 avdd.n548 avdd.n539 300.048
R528 avdd.n542 avdd.n539 300.048
R529 avdd.n359 avdd.n302 295.529
R530 avdd.n607 avdd.n550 295.529
R531 avdd.t524 avdd.n287 289.247
R532 avdd.t609 avdd.n535 289.247
R533 avdd.n495 avdd.n282 281.601
R534 avdd.n919 avdd.n530 281.601
R535 avdd.n759 avdd.t345 280.161
R536 avdd.n752 avdd.t353 279.486
R537 avdd.n8 avdd.n7 271.068
R538 avdd.n1153 avdd.n1152 271.068
R539 avdd.n1132 avdd.n1131 271.068
R540 avdd.n1111 avdd.n1110 271.068
R541 avdd.n1090 avdd.n1089 271.068
R542 avdd.n1069 avdd.n1068 271.068
R543 avdd.n1048 avdd.n1047 271.068
R544 avdd.n1027 avdd.n1026 271.068
R545 avdd.n1006 avdd.n1005 271.068
R546 avdd.n1526 avdd.n1525 271.068
R547 avdd.n1505 avdd.n1504 271.068
R548 avdd.n1484 avdd.n1483 271.068
R549 avdd.n1463 avdd.n1462 271.068
R550 avdd.n1442 avdd.n1441 271.068
R551 avdd.n1421 avdd.n1420 271.068
R552 avdd.n1400 avdd.n1399 271.068
R553 avdd.n1379 avdd.n1378 271.068
R554 avdd.n1823 avdd.n1740 257.882
R555 avdd.n1763 avdd.n1741 257.882
R556 avdd.n786 avdd.t444 257.603
R557 avdd.n760 avdd.t281 256.101
R558 avdd.n1772 avdd.t378 255.679
R559 avdd.t380 avdd.n1772 255.679
R560 avdd.n127 avdd.t508 252.983
R561 avdd.n121 avdd.t259 252.983
R562 avdd.n140 avdd.t1 252.983
R563 avdd.n152 avdd.t450 252.983
R564 avdd.n101 avdd.t601 252.983
R565 avdd.n165 avdd.t467 252.983
R566 avdd.n177 avdd.t593 252.983
R567 avdd.n81 avdd.t436 252.983
R568 avdd.n190 avdd.t424 252.983
R569 avdd.n202 avdd.t519 252.983
R570 avdd.n61 avdd.t474 252.983
R571 avdd.n215 avdd.t179 252.983
R572 avdd.n227 avdd.t573 252.983
R573 avdd.n41 avdd.t504 252.983
R574 avdd.n240 avdd.t391 252.983
R575 avdd.n251 avdd.t620 252.983
R576 avdd.n12 avdd.t616 252.983
R577 avdd.n788 avdd.t275 252.983
R578 avdd.n1876 avdd.n1875 241.459
R579 avdd.n1875 avdd.n17 240.66
R580 avdd.n1872 avdd.n1871 240.66
R581 avdd.n1872 avdd.n20 240.66
R582 avdd.t481 avdd.t491 233.565
R583 avdd.t491 avdd.t487 233.565
R584 avdd.t487 avdd.t485 233.565
R585 avdd.t485 avdd.t477 233.565
R586 avdd.t483 avdd.t489 233.565
R587 avdd.t479 avdd.t483 233.565
R588 avdd.t501 avdd.t479 233.565
R589 avdd.t499 avdd.t501 233.565
R590 avdd.t540 avdd.t532 233.565
R591 avdd.t532 avdd.t528 233.565
R592 avdd.t528 avdd.t538 233.565
R593 avdd.t538 avdd.t536 233.565
R594 avdd.t542 avdd.t530 233.565
R595 avdd.t534 avdd.t542 233.565
R596 avdd.t546 avdd.t534 233.565
R597 avdd.t544 avdd.t546 233.565
R598 avdd.n521 avdd.t523 232.686
R599 avdd.n945 avdd.t608 232.686
R600 avdd.n435 avdd.t482 231.989
R601 avdd.n444 avdd.t500 231.989
R602 avdd.n859 avdd.t541 231.989
R603 avdd.n868 avdd.t545 231.989
R604 avdd.n522 avdd.t521 231.974
R605 avdd.n521 avdd.t525 231.974
R606 avdd.n946 avdd.t606 231.974
R607 avdd.n945 avdd.t610 231.974
R608 avdd.n518 avdd.t58 227.478
R609 avdd.n516 avdd.t22 227.478
R610 avdd.n514 avdd.t19 227.478
R611 avdd.n512 avdd.t8 227.478
R612 avdd.n510 avdd.t11 227.478
R613 avdd.n508 avdd.t174 227.478
R614 avdd.n506 avdd.t5 227.478
R615 avdd.n504 avdd.t123 227.478
R616 avdd.n502 avdd.t167 227.478
R617 avdd.n500 avdd.t134 227.478
R618 avdd.n498 avdd.t126 227.478
R619 avdd.n431 avdd.t128 227.478
R620 avdd.t85 avdd.n426 227.478
R621 avdd.t78 avdd.n423 227.478
R622 avdd.n420 avdd.t60 227.478
R623 avdd.n417 avdd.t62 227.478
R624 avdd.t48 avdd.n412 227.478
R625 avdd.t55 avdd.n409 227.478
R626 avdd.n406 avdd.t14 227.478
R627 avdd.n403 avdd.t42 227.478
R628 avdd.t147 avdd.n398 227.478
R629 avdd.t145 avdd.n395 227.478
R630 avdd.n942 avdd.t155 227.478
R631 avdd.n940 avdd.t111 227.478
R632 avdd.n938 avdd.t150 227.478
R633 avdd.n936 avdd.t102 227.478
R634 avdd.n934 avdd.t139 227.478
R635 avdd.n932 avdd.t93 227.478
R636 avdd.n930 avdd.t90 227.478
R637 avdd.n928 avdd.t81 227.478
R638 avdd.n926 avdd.t76 227.478
R639 avdd.n924 avdd.t29 227.478
R640 avdd.n922 avdd.t65 227.478
R641 avdd.n854 avdd.t159 227.478
R642 avdd.t113 avdd.n849 227.478
R643 avdd.t152 avdd.n846 227.478
R644 avdd.n843 avdd.t104 227.478
R645 avdd.n840 avdd.t143 227.478
R646 avdd.t97 avdd.n835 227.478
R647 avdd.t95 avdd.n832 227.478
R648 avdd.n829 avdd.t87 227.478
R649 avdd.n826 avdd.t83 227.478
R650 avdd.t34 avdd.n821 227.478
R651 avdd.t71 avdd.n818 227.478
R652 avdd.n279 avdd.t51 227.345
R653 avdd.t69 avdd.n459 227.345
R654 avdd.n527 avdd.t131 227.345
R655 avdd.t136 avdd.n883 227.345
R656 avdd.n1181 avdd.t216 217.947
R657 avdd.n352 avdd.n282 211.953
R658 avdd.n600 avdd.n530 211.953
R659 avdd.n1815 avdd.t35 211.924
R660 avdd.n360 avdd.n359 210.825
R661 avdd.n608 avdd.n607 210.825
R662 avdd.n482 avdd.n481 204.31
R663 avdd.n461 avdd.n460 204.31
R664 avdd.n336 avdd.n335 204.31
R665 avdd.n906 avdd.n905 204.31
R666 avdd.n885 avdd.n884 204.31
R667 avdd.n584 avdd.n583 204.31
R668 avdd.n437 avdd.n436 204.294
R669 avdd.n439 avdd.n438 204.294
R670 avdd.n441 avdd.n440 204.294
R671 avdd.n443 avdd.n442 204.294
R672 avdd.n861 avdd.n860 204.294
R673 avdd.n863 avdd.n862 204.294
R674 avdd.n865 avdd.n864 204.294
R675 avdd.n867 avdd.n866 204.294
R676 avdd.n387 avdd.n386 204.284
R677 avdd.n385 avdd.n384 204.284
R678 avdd.n383 avdd.n382 204.284
R679 avdd.n381 avdd.n380 204.284
R680 avdd.n379 avdd.n378 204.284
R681 avdd.n377 avdd.n376 204.284
R682 avdd.n375 avdd.n374 204.284
R683 avdd.n373 avdd.n372 204.284
R684 avdd.n371 avdd.n370 204.284
R685 avdd.n369 avdd.n368 204.284
R686 avdd.n308 avdd.n307 204.284
R687 avdd.n430 avdd.n429 204.284
R688 avdd.n428 avdd.n427 204.284
R689 avdd.n425 avdd.n424 204.284
R690 avdd.n419 avdd.n391 204.284
R691 avdd.n416 avdd.n415 204.284
R692 avdd.n414 avdd.n413 204.284
R693 avdd.n411 avdd.n410 204.284
R694 avdd.n405 avdd.n393 204.284
R695 avdd.n402 avdd.n401 204.284
R696 avdd.n400 avdd.n399 204.284
R697 avdd.n397 avdd.n396 204.284
R698 avdd.n313 avdd.n312 204.284
R699 avdd.n315 avdd.n314 204.284
R700 avdd.n317 avdd.n316 204.284
R701 avdd.n319 avdd.n318 204.284
R702 avdd.n321 avdd.n320 204.284
R703 avdd.n323 avdd.n322 204.284
R704 avdd.n325 avdd.n324 204.284
R705 avdd.n327 avdd.n326 204.284
R706 avdd.n329 avdd.n328 204.284
R707 avdd.n331 avdd.n330 204.284
R708 avdd.n333 avdd.n332 204.284
R709 avdd.n810 avdd.n809 204.284
R710 avdd.n808 avdd.n807 204.284
R711 avdd.n806 avdd.n805 204.284
R712 avdd.n804 avdd.n803 204.284
R713 avdd.n802 avdd.n801 204.284
R714 avdd.n800 avdd.n799 204.284
R715 avdd.n798 avdd.n797 204.284
R716 avdd.n796 avdd.n795 204.284
R717 avdd.n794 avdd.n793 204.284
R718 avdd.n792 avdd.n791 204.284
R719 avdd.n556 avdd.n555 204.284
R720 avdd.n853 avdd.n852 204.284
R721 avdd.n851 avdd.n850 204.284
R722 avdd.n848 avdd.n847 204.284
R723 avdd.n842 avdd.n814 204.284
R724 avdd.n839 avdd.n838 204.284
R725 avdd.n837 avdd.n836 204.284
R726 avdd.n834 avdd.n833 204.284
R727 avdd.n828 avdd.n816 204.284
R728 avdd.n825 avdd.n824 204.284
R729 avdd.n823 avdd.n822 204.284
R730 avdd.n820 avdd.n819 204.284
R731 avdd.n561 avdd.n560 204.284
R732 avdd.n563 avdd.n562 204.284
R733 avdd.n565 avdd.n564 204.284
R734 avdd.n567 avdd.n566 204.284
R735 avdd.n569 avdd.n568 204.284
R736 avdd.n571 avdd.n570 204.284
R737 avdd.n573 avdd.n572 204.284
R738 avdd.n575 avdd.n574 204.284
R739 avdd.n577 avdd.n576 204.284
R740 avdd.n579 avdd.n578 204.284
R741 avdd.n581 avdd.n580 204.284
R742 avdd.n1752 avdd.n1736 203.672
R743 avdd.n1816 avdd.n1760 203.672
R744 avdd.n353 avdd.n352 201.788
R745 avdd.n601 avdd.n600 201.788
R746 avdd.n667 avdd.t352 201.107
R747 avdd.n1151 avdd.t461 197.562
R748 avdd.n1130 avdd.t264 197.562
R749 avdd.n1109 avdd.t212 197.562
R750 avdd.n1088 avdd.t320 197.562
R751 avdd.n1067 avdd.t475 197.562
R752 avdd.n1046 avdd.t270 197.562
R753 avdd.n1025 avdd.t505 197.562
R754 avdd.n1004 avdd.t431 197.562
R755 avdd.n1524 avdd.t427 197.562
R756 avdd.n1503 avdd.t304 197.562
R757 avdd.n1482 avdd.t437 197.562
R758 avdd.n1461 avdd.t651 197.562
R759 avdd.n1440 avdd.t456 197.562
R760 avdd.n1419 avdd.t262 197.562
R761 avdd.n1398 avdd.t515 197.562
R762 avdd.n1377 avdd.t494 197.562
R763 avdd.n1812 avdd.n1741 196.142
R764 avdd.t522 avdd.n287 195.042
R765 avdd.t607 avdd.n535 195.042
R766 avdd.t311 avdd.n979 193.774
R767 avdd.t272 avdd.n1352 193.774
R768 avdd.n353 avdd.n301 186.353
R769 avdd.n601 avdd.n549 186.353
R770 avdd.n249 avdd.n248 185
R771 avdd.n248 avdd.n247 185
R772 avdd.n29 avdd.n28 185
R773 avdd.n246 avdd.n29 185
R774 avdd.n244 avdd.n243 185
R775 avdd.n245 avdd.n244 185
R776 avdd.n238 avdd.n237 185
R777 avdd.n237 avdd.n32 185
R778 avdd.n236 avdd.n35 185
R779 avdd.n236 avdd.n235 185
R780 avdd.n38 avdd.n36 185
R781 avdd.n234 avdd.n36 185
R782 avdd.n232 avdd.n231 185
R783 avdd.n233 avdd.n232 185
R784 avdd.n230 avdd.n37 185
R785 avdd.n49 avdd.n37 185
R786 avdd.n50 avdd.n44 185
R787 avdd.n51 avdd.n50 185
R788 avdd.n224 avdd.n223 185
R789 avdd.n223 avdd.n222 185
R790 avdd.n48 avdd.n47 185
R791 avdd.n221 avdd.n48 185
R792 avdd.n219 avdd.n218 185
R793 avdd.n220 avdd.n219 185
R794 avdd.n213 avdd.n212 185
R795 avdd.n212 avdd.n52 185
R796 avdd.n211 avdd.n55 185
R797 avdd.n211 avdd.n210 185
R798 avdd.n58 avdd.n56 185
R799 avdd.n209 avdd.n56 185
R800 avdd.n207 avdd.n206 185
R801 avdd.n208 avdd.n207 185
R802 avdd.n205 avdd.n57 185
R803 avdd.n69 avdd.n57 185
R804 avdd.n70 avdd.n64 185
R805 avdd.n71 avdd.n70 185
R806 avdd.n199 avdd.n198 185
R807 avdd.n198 avdd.n197 185
R808 avdd.n68 avdd.n67 185
R809 avdd.n196 avdd.n68 185
R810 avdd.n194 avdd.n193 185
R811 avdd.n195 avdd.n194 185
R812 avdd.n188 avdd.n187 185
R813 avdd.n187 avdd.n72 185
R814 avdd.n186 avdd.n75 185
R815 avdd.n186 avdd.n185 185
R816 avdd.n78 avdd.n76 185
R817 avdd.n184 avdd.n76 185
R818 avdd.n182 avdd.n181 185
R819 avdd.n183 avdd.n182 185
R820 avdd.n180 avdd.n77 185
R821 avdd.n89 avdd.n77 185
R822 avdd.n90 avdd.n84 185
R823 avdd.n91 avdd.n90 185
R824 avdd.n174 avdd.n173 185
R825 avdd.n173 avdd.n172 185
R826 avdd.n88 avdd.n87 185
R827 avdd.n171 avdd.n88 185
R828 avdd.n169 avdd.n168 185
R829 avdd.n170 avdd.n169 185
R830 avdd.n163 avdd.n162 185
R831 avdd.n162 avdd.n92 185
R832 avdd.n161 avdd.n95 185
R833 avdd.n161 avdd.n160 185
R834 avdd.n98 avdd.n96 185
R835 avdd.n159 avdd.n96 185
R836 avdd.n157 avdd.n156 185
R837 avdd.n158 avdd.n157 185
R838 avdd.n155 avdd.n97 185
R839 avdd.n109 avdd.n97 185
R840 avdd.n110 avdd.n104 185
R841 avdd.n111 avdd.n110 185
R842 avdd.n149 avdd.n148 185
R843 avdd.n148 avdd.n147 185
R844 avdd.n108 avdd.n107 185
R845 avdd.n146 avdd.n108 185
R846 avdd.n144 avdd.n143 185
R847 avdd.n145 avdd.n144 185
R848 avdd.n138 avdd.n137 185
R849 avdd.n137 avdd.n112 185
R850 avdd.n136 avdd.n115 185
R851 avdd.n136 avdd.n135 185
R852 avdd.n118 avdd.n116 185
R853 avdd.n134 avdd.n116 185
R854 avdd.n132 avdd.n131 185
R855 avdd.n133 avdd.n132 185
R856 avdd.n130 avdd.n117 185
R857 avdd.n256 avdd.n23 185
R858 avdd.n255 avdd.n24 185
R859 avdd.n30 avdd.n24 185
R860 avdd.n254 avdd.n25 185
R861 avdd.n31 avdd.n25 185
R862 avdd.n5 avdd.n3 185
R863 avdd.n6 avdd.n5 185
R864 avdd.n9 avdd.n4 185
R865 avdd.n1208 avdd.n1138 185
R866 avdd.n1151 avdd.n1138 185
R867 avdd.n1207 avdd.n1139 185
R868 avdd.n1148 avdd.n1140 185
R869 avdd.n1149 avdd.n1144 185
R870 avdd.n1200 avdd.n1145 185
R871 avdd.n1199 avdd.n1146 185
R872 avdd.n1223 avdd.n1117 185
R873 avdd.n1130 avdd.n1117 185
R874 avdd.n1222 avdd.n1118 185
R875 avdd.n1127 avdd.n1119 185
R876 avdd.n1128 avdd.n1123 185
R877 avdd.n1215 avdd.n1124 185
R878 avdd.n1214 avdd.n1125 185
R879 avdd.n1238 avdd.n1096 185
R880 avdd.n1109 avdd.n1096 185
R881 avdd.n1237 avdd.n1097 185
R882 avdd.n1106 avdd.n1098 185
R883 avdd.n1107 avdd.n1102 185
R884 avdd.n1230 avdd.n1103 185
R885 avdd.n1229 avdd.n1104 185
R886 avdd.n1253 avdd.n1075 185
R887 avdd.n1088 avdd.n1075 185
R888 avdd.n1252 avdd.n1076 185
R889 avdd.n1085 avdd.n1077 185
R890 avdd.n1086 avdd.n1081 185
R891 avdd.n1245 avdd.n1082 185
R892 avdd.n1244 avdd.n1083 185
R893 avdd.n1268 avdd.n1054 185
R894 avdd.n1067 avdd.n1054 185
R895 avdd.n1267 avdd.n1055 185
R896 avdd.n1064 avdd.n1056 185
R897 avdd.n1065 avdd.n1060 185
R898 avdd.n1260 avdd.n1061 185
R899 avdd.n1259 avdd.n1062 185
R900 avdd.n1283 avdd.n1033 185
R901 avdd.n1046 avdd.n1033 185
R902 avdd.n1282 avdd.n1034 185
R903 avdd.n1043 avdd.n1035 185
R904 avdd.n1044 avdd.n1039 185
R905 avdd.n1275 avdd.n1040 185
R906 avdd.n1274 avdd.n1041 185
R907 avdd.n1298 avdd.n1012 185
R908 avdd.n1025 avdd.n1012 185
R909 avdd.n1297 avdd.n1013 185
R910 avdd.n1022 avdd.n1014 185
R911 avdd.n1023 avdd.n1018 185
R912 avdd.n1290 avdd.n1019 185
R913 avdd.n1289 avdd.n1020 185
R914 avdd.n1313 avdd.n991 185
R915 avdd.n1004 avdd.n991 185
R916 avdd.n1312 avdd.n992 185
R917 avdd.n1001 avdd.n993 185
R918 avdd.n1002 avdd.n997 185
R919 avdd.n1305 avdd.n998 185
R920 avdd.n1304 avdd.n999 185
R921 avdd.n1348 avdd.n979 185
R922 avdd.n1347 avdd.n980 185
R923 avdd.n1320 avdd.n980 185
R924 avdd.n1321 avdd.n981 185
R925 avdd.n1322 avdd.n1321 185
R926 avdd.n1343 avdd.n986 185
R927 avdd.n1323 avdd.n986 185
R928 avdd.n1342 avdd.n987 185
R929 avdd.n1324 avdd.n987 185
R930 avdd.n1325 avdd.n988 185
R931 avdd.n1326 avdd.n1325 185
R932 avdd.n1319 avdd.n1318 185
R933 avdd.n1327 avdd.n1319 185
R934 avdd.n1330 avdd.n1329 185
R935 avdd.n1329 avdd.n1328 185
R936 avdd.n1545 avdd.n1511 185
R937 avdd.n1524 avdd.n1511 185
R938 avdd.n1544 avdd.n1512 185
R939 avdd.n1521 avdd.n1513 185
R940 avdd.n1522 avdd.n1517 185
R941 avdd.n1537 avdd.n1518 185
R942 avdd.n1536 avdd.n1519 185
R943 avdd.n1560 avdd.n1490 185
R944 avdd.n1503 avdd.n1490 185
R945 avdd.n1559 avdd.n1491 185
R946 avdd.n1500 avdd.n1492 185
R947 avdd.n1501 avdd.n1496 185
R948 avdd.n1552 avdd.n1497 185
R949 avdd.n1551 avdd.n1498 185
R950 avdd.n1575 avdd.n1469 185
R951 avdd.n1482 avdd.n1469 185
R952 avdd.n1574 avdd.n1470 185
R953 avdd.n1479 avdd.n1471 185
R954 avdd.n1480 avdd.n1475 185
R955 avdd.n1567 avdd.n1476 185
R956 avdd.n1566 avdd.n1477 185
R957 avdd.n1590 avdd.n1448 185
R958 avdd.n1461 avdd.n1448 185
R959 avdd.n1589 avdd.n1449 185
R960 avdd.n1458 avdd.n1450 185
R961 avdd.n1459 avdd.n1454 185
R962 avdd.n1582 avdd.n1455 185
R963 avdd.n1581 avdd.n1456 185
R964 avdd.n1605 avdd.n1427 185
R965 avdd.n1440 avdd.n1427 185
R966 avdd.n1604 avdd.n1428 185
R967 avdd.n1437 avdd.n1429 185
R968 avdd.n1438 avdd.n1433 185
R969 avdd.n1597 avdd.n1434 185
R970 avdd.n1596 avdd.n1435 185
R971 avdd.n1620 avdd.n1406 185
R972 avdd.n1419 avdd.n1406 185
R973 avdd.n1619 avdd.n1407 185
R974 avdd.n1416 avdd.n1408 185
R975 avdd.n1417 avdd.n1412 185
R976 avdd.n1612 avdd.n1413 185
R977 avdd.n1611 avdd.n1414 185
R978 avdd.n1635 avdd.n1385 185
R979 avdd.n1398 avdd.n1385 185
R980 avdd.n1634 avdd.n1386 185
R981 avdd.n1395 avdd.n1387 185
R982 avdd.n1396 avdd.n1391 185
R983 avdd.n1627 avdd.n1392 185
R984 avdd.n1626 avdd.n1393 185
R985 avdd.n1650 avdd.n1364 185
R986 avdd.n1377 avdd.n1364 185
R987 avdd.n1649 avdd.n1365 185
R988 avdd.n1374 avdd.n1366 185
R989 avdd.n1375 avdd.n1370 185
R990 avdd.n1642 avdd.n1371 185
R991 avdd.n1641 avdd.n1372 185
R992 avdd.n1685 avdd.n1352 185
R993 avdd.n1684 avdd.n1353 185
R994 avdd.n1657 avdd.n1353 185
R995 avdd.n1658 avdd.n1354 185
R996 avdd.n1659 avdd.n1658 185
R997 avdd.n1680 avdd.n1359 185
R998 avdd.n1660 avdd.n1359 185
R999 avdd.n1679 avdd.n1360 185
R1000 avdd.n1661 avdd.n1360 185
R1001 avdd.n1662 avdd.n1361 185
R1002 avdd.n1663 avdd.n1662 185
R1003 avdd.n1656 avdd.n1655 185
R1004 avdd.n1664 avdd.n1656 185
R1005 avdd.n1667 avdd.n1666 185
R1006 avdd.n1666 avdd.n1665 185
R1007 avdd.n1180 avdd.n1179 185
R1008 avdd.n1181 avdd.n1180 185
R1009 avdd.n1165 avdd.n1164 185
R1010 avdd.n1171 avdd.n1170 185
R1011 avdd.n1169 avdd.n1160 185
R1012 avdd.n1184 avdd.n1161 185
R1013 avdd.n1183 avdd.n1182 185
R1014 avdd.n1182 avdd.n1181 185
R1015 avdd.n666 avdd.n665 185
R1016 avdd.n664 avdd.n663 185
R1017 avdd.n663 avdd.n662 185
R1018 avdd.n672 avdd.n671 185
R1019 avdd.n673 avdd.n672 185
R1020 avdd.n661 avdd.n660 185
R1021 avdd.n674 avdd.n661 185
R1022 avdd.n678 avdd.n677 185
R1023 avdd.n677 avdd.n676 185
R1024 avdd.n658 avdd.n657 185
R1025 avdd.n675 avdd.n657 185
R1026 avdd.n683 avdd.n682 185
R1027 avdd.n684 avdd.n683 185
R1028 avdd.n656 avdd.n655 185
R1029 avdd.n685 avdd.n656 185
R1030 avdd.n688 avdd.n687 185
R1031 avdd.n687 avdd.n686 185
R1032 avdd.n653 avdd.n652 185
R1033 avdd.n652 avdd.n651 185
R1034 avdd.n693 avdd.n692 185
R1035 avdd.n694 avdd.n693 185
R1036 avdd.n650 avdd.n649 185
R1037 avdd.n695 avdd.n650 185
R1038 avdd.n699 avdd.n698 185
R1039 avdd.n698 avdd.n697 185
R1040 avdd.n647 avdd.n646 185
R1041 avdd.n696 avdd.n646 185
R1042 avdd.n704 avdd.n703 185
R1043 avdd.n705 avdd.n704 185
R1044 avdd.n645 avdd.n644 185
R1045 avdd.n706 avdd.n645 185
R1046 avdd.n709 avdd.n708 185
R1047 avdd.n708 avdd.n707 185
R1048 avdd.n642 avdd.n641 185
R1049 avdd.n641 avdd.n640 185
R1050 avdd.n714 avdd.n713 185
R1051 avdd.n715 avdd.n714 185
R1052 avdd.n639 avdd.n638 185
R1053 avdd.n716 avdd.n639 185
R1054 avdd.n720 avdd.n719 185
R1055 avdd.n719 avdd.n718 185
R1056 avdd.n636 avdd.n635 185
R1057 avdd.n717 avdd.n635 185
R1058 avdd.n725 avdd.n724 185
R1059 avdd.n726 avdd.n725 185
R1060 avdd.n634 avdd.n633 185
R1061 avdd.n727 avdd.n634 185
R1062 avdd.n731 avdd.n730 185
R1063 avdd.n730 avdd.n729 185
R1064 avdd.n631 avdd.n630 185
R1065 avdd.n728 avdd.n630 185
R1066 avdd.n736 avdd.n735 185
R1067 avdd.n737 avdd.n736 185
R1068 avdd.n629 avdd.n628 185
R1069 avdd.n738 avdd.n629 185
R1070 avdd.n742 avdd.n741 185
R1071 avdd.n741 avdd.n740 185
R1072 avdd.n625 avdd.n624 185
R1073 avdd.n739 avdd.n624 185
R1074 avdd.n768 avdd.n767 185
R1075 avdd.n769 avdd.n768 185
R1076 avdd.n626 avdd.n622 185
R1077 avdd.n770 avdd.n622 185
R1078 avdd.n772 avdd.n623 185
R1079 avdd.n772 avdd.n771 185
R1080 avdd.n773 avdd.n617 185
R1081 avdd.n774 avdd.n773 185
R1082 avdd.n783 avdd.n618 185
R1083 avdd.n775 avdd.n618 185
R1084 avdd.n782 avdd.n619 185
R1085 avdd.n776 avdd.n619 185
R1086 avdd.n621 avdd.n620 185
R1087 avdd.n452 avdd.t13 180.231
R1088 avdd.n492 avdd.t3 180.231
R1089 avdd.n876 avdd.t33 180.231
R1090 avdd.n916 avdd.t27 180.231
R1091 avdd.n31 avdd.n30 175.386
R1092 avdd.n246 avdd.n245 175.386
R1093 avdd.n235 avdd.n234 175.386
R1094 avdd.n51 avdd.n49 175.386
R1095 avdd.n221 avdd.n220 175.386
R1096 avdd.n210 avdd.n209 175.386
R1097 avdd.n71 avdd.n69 175.386
R1098 avdd.n196 avdd.n195 175.386
R1099 avdd.n185 avdd.n184 175.386
R1100 avdd.n91 avdd.n89 175.386
R1101 avdd.n171 avdd.n170 175.386
R1102 avdd.n160 avdd.n159 175.386
R1103 avdd.n111 avdd.n109 175.386
R1104 avdd.n146 avdd.n145 175.386
R1105 avdd.n135 avdd.n134 175.386
R1106 avdd.n673 avdd.n662 175.386
R1107 avdd.n676 avdd.n675 175.386
R1108 avdd.n685 avdd.n684 175.386
R1109 avdd.n694 avdd.n651 175.386
R1110 avdd.n697 avdd.n695 175.386
R1111 avdd.n706 avdd.n705 175.386
R1112 avdd.n715 avdd.n640 175.386
R1113 avdd.n718 avdd.n716 175.386
R1114 avdd.n727 avdd.n726 175.386
R1115 avdd.n729 avdd.n728 175.386
R1116 avdd.n738 avdd.n737 175.386
R1117 avdd.n740 avdd.n739 175.386
R1118 avdd.n770 avdd.n769 175.386
R1119 avdd.n775 avdd.n774 175.386
R1120 avdd.n776 avdd.n775 175.386
R1121 avdd.n247 avdd.t390 169.905
R1122 avdd.t503 avdd.n32 169.905
R1123 avdd.n233 avdd.t572 169.905
R1124 avdd.n222 avdd.t178 169.905
R1125 avdd.t473 avdd.n52 169.905
R1126 avdd.n208 avdd.t518 169.905
R1127 avdd.n197 avdd.t423 169.905
R1128 avdd.t435 avdd.n72 169.905
R1129 avdd.n183 avdd.t592 169.905
R1130 avdd.n172 avdd.t466 169.905
R1131 avdd.t600 avdd.n92 169.905
R1132 avdd.n158 avdd.t449 169.905
R1133 avdd.n147 avdd.t0 169.905
R1134 avdd.t258 avdd.n112 169.905
R1135 avdd.n133 avdd.t507 169.905
R1136 avdd.t443 avdd.n776 169.905
R1137 avdd.t322 avdd.n674 168.077
R1138 avdd.n707 avdd.t326 168.077
R1139 avdd.t579 avdd.n1762 167.023
R1140 avdd.n1816 avdd.n1815 165.936
R1141 avdd.t280 avdd.n738 162.596
R1142 avdd.t338 avdd.n696 160.769
R1143 avdd.n737 avdd.t344 160.769
R1144 avdd.n1818 avdd.n1817 155.859
R1145 avdd.n1822 avdd.n1821 155.859
R1146 avdd.n486 avdd.t182 155.153
R1147 avdd.n486 avdd.t195 155.153
R1148 avdd.n910 avdd.t403 155.153
R1149 avdd.n910 avdd.t392 155.153
R1150 avdd.n758 avdd.n745 154.113
R1151 avdd.n757 avdd.n746 154.113
R1152 avdd.n756 avdd.n747 154.113
R1153 avdd.n755 avdd.n748 154.113
R1154 avdd.n754 avdd.n749 154.113
R1155 avdd.n753 avdd.n750 154.113
R1156 avdd.n752 avdd.n751 154.113
R1157 avdd.n762 avdd.n761 154.042
R1158 avdd.t36 avdd.t579 153.764
R1159 avdd.n1142 avdd.n1141 153.571
R1160 avdd.n1121 avdd.n1120 153.571
R1161 avdd.n1100 avdd.n1099 153.571
R1162 avdd.n1079 avdd.n1078 153.571
R1163 avdd.n1058 avdd.n1057 153.571
R1164 avdd.n1037 avdd.n1036 153.571
R1165 avdd.n1016 avdd.n1015 153.571
R1166 avdd.n995 avdd.n994 153.571
R1167 avdd.n1337 avdd.n1336 153.571
R1168 avdd.n1515 avdd.n1514 153.571
R1169 avdd.n1494 avdd.n1493 153.571
R1170 avdd.n1473 avdd.n1472 153.571
R1171 avdd.n1452 avdd.n1451 153.571
R1172 avdd.n1431 avdd.n1430 153.571
R1173 avdd.n1410 avdd.n1409 153.571
R1174 avdd.n1389 avdd.n1388 153.571
R1175 avdd.n1368 avdd.n1367 153.571
R1176 avdd.n1674 avdd.n1673 153.571
R1177 avdd.n1168 avdd.n1167 153.571
R1178 avdd.t218 avdd.n1858 149.893
R1179 avdd.n1860 avdd.t246 149.893
R1180 avdd.t434 avdd.n1873 149.893
R1181 avdd.n1874 avdd.t429 149.893
R1182 avdd.n686 avdd.t330 146.155
R1183 avdd.n717 avdd.t340 146.155
R1184 avdd.n771 avdd.t276 144.327
R1185 avdd.n771 avdd.t274 140.673
R1186 avdd.n686 avdd.t328 138.846
R1187 avdd.t334 avdd.n717 138.846
R1188 avdd.n1861 avdd.n1855 125.742
R1189 avdd.n1853 avdd.n1836 125.742
R1190 avdd.n696 avdd.t324 124.231
R1191 avdd.t611 avdd.t577 121.877
R1192 avdd.t613 avdd.t603 121.877
R1193 avdd.n1322 avdd.n1320 120.317
R1194 avdd.n1324 avdd.n1323 120.317
R1195 avdd.n1327 avdd.n1326 120.317
R1196 avdd.n1328 avdd.n1327 120.317
R1197 avdd.n1661 avdd.n1660 120.317
R1198 avdd.n1664 avdd.n1663 120.317
R1199 avdd.n1665 avdd.n1664 120.317
R1200 avdd.n1659 avdd.n1657 119.064
R1201 avdd.n1181 avdd.t657 117.838
R1202 avdd.n674 avdd.t348 116.924
R1203 avdd.n707 avdd.t346 116.924
R1204 avdd.n448 avdd.t477 116.782
R1205 avdd.n448 avdd.t489 116.782
R1206 avdd.n872 avdd.t536 116.782
R1207 avdd.n872 avdd.t530 116.782
R1208 avdd.t657 avdd.t445 112.624
R1209 avdd.t222 avdd.t218 110.959
R1210 avdd.t248 avdd.t222 110.959
R1211 avdd.t244 avdd.t248 110.959
R1212 avdd.t240 avdd.t244 110.959
R1213 avdd.t228 avdd.t240 110.959
R1214 avdd.t230 avdd.t228 110.959
R1215 avdd.t226 avdd.t230 110.959
R1216 avdd.t238 avdd.t224 110.959
R1217 avdd.t236 avdd.t238 110.959
R1218 avdd.t242 avdd.t236 110.959
R1219 avdd.t234 avdd.t242 110.959
R1220 avdd.t232 avdd.t234 110.959
R1221 avdd.t220 avdd.t232 110.959
R1222 avdd.t246 avdd.t220 110.959
R1223 avdd.t433 avdd.t434 110.959
R1224 avdd.t171 avdd.t433 110.959
R1225 avdd.t559 avdd.t171 110.959
R1226 avdd.t558 avdd.t559 110.959
R1227 avdd.t40 avdd.t558 110.959
R1228 avdd.t458 avdd.t40 110.959
R1229 avdd.t459 avdd.t458 110.959
R1230 avdd.t16 avdd.t459 110.959
R1231 avdd.t471 avdd.t16 110.959
R1232 avdd.t470 avdd.t471 110.959
R1233 avdd.t73 avdd.t470 110.959
R1234 avdd.t261 avdd.t73 110.959
R1235 avdd.t260 avdd.t261 110.959
R1236 avdd.t169 avdd.t260 110.959
R1237 avdd.t591 avdd.t169 110.959
R1238 avdd.t590 avdd.t591 110.959
R1239 avdd.t157 avdd.t590 110.959
R1240 avdd.t465 avdd.t157 110.959
R1241 avdd.t464 avdd.t465 110.959
R1242 avdd.t106 avdd.t464 110.959
R1243 avdd.t426 avdd.t106 110.959
R1244 avdd.t425 avdd.t426 110.959
R1245 avdd.t38 avdd.t425 110.959
R1246 avdd.t653 avdd.t38 110.959
R1247 avdd.t654 avdd.t653 110.959
R1248 avdd.t141 avdd.t654 110.959
R1249 avdd.t595 avdd.t141 110.959
R1250 avdd.t594 avdd.t595 110.959
R1251 avdd.t67 avdd.t594 110.959
R1252 avdd.t469 avdd.t67 110.959
R1253 avdd.t468 avdd.t469 110.959
R1254 avdd.t164 avdd.t468 110.959
R1255 avdd.t561 avdd.t164 110.959
R1256 avdd.t560 avdd.t561 110.959
R1257 avdd.t118 avdd.t560 110.959
R1258 avdd.t451 avdd.t118 110.959
R1259 avdd.t452 avdd.t451 110.959
R1260 avdd.t31 avdd.t452 110.959
R1261 avdd.t526 avdd.t31 110.959
R1262 avdd.t527 avdd.t526 110.959
R1263 avdd.t99 avdd.t527 110.959
R1264 avdd.t215 avdd.t99 110.959
R1265 avdd.t214 avdd.t215 110.959
R1266 avdd.t53 avdd.t214 110.959
R1267 avdd.t430 avdd.t53 110.959
R1268 avdd.t429 avdd.t430 110.959
R1269 avdd.n1151 avdd.t296 106.817
R1270 avdd.n1130 avdd.t512 106.817
R1271 avdd.n1109 avdd.t300 106.817
R1272 avdd.n1088 avdd.t315 106.817
R1273 avdd.n1067 avdd.t421 106.817
R1274 avdd.n1046 avdd.t588 106.817
R1275 avdd.n1025 avdd.t288 106.817
R1276 avdd.n1004 avdd.t307 106.817
R1277 avdd.n1524 avdd.t510 106.817
R1278 avdd.n1503 avdd.t598 106.817
R1279 avdd.n1482 avdd.t563 106.817
R1280 avdd.n1461 avdd.t567 106.817
R1281 avdd.n1440 avdd.t282 106.817
R1282 avdd.n1419 avdd.t256 106.817
R1283 avdd.n1398 avdd.t266 106.817
R1284 avdd.n1377 avdd.t208 106.817
R1285 avdd.t294 avdd.n1322 106.531
R1286 avdd.t447 avdd.n1659 106.531
R1287 avdd.n489 avdd.n301 105.412
R1288 avdd.n913 avdd.n549 105.412
R1289 avdd.n675 avdd.t350 102.308
R1290 avdd.t332 avdd.n715 102.308
R1291 avdd.t296 avdd.t298 102.091
R1292 avdd.t512 avdd.t453 102.091
R1293 avdd.t300 avdd.t302 102.091
R1294 avdd.t315 avdd.t317 102.091
R1295 avdd.t421 avdd.t419 102.091
R1296 avdd.t588 avdd.t556 102.091
R1297 avdd.t288 avdd.t286 102.091
R1298 avdd.t307 avdd.t292 102.091
R1299 avdd.t510 avdd.t309 102.091
R1300 avdd.t598 avdd.t596 102.091
R1301 avdd.t563 avdd.t313 102.091
R1302 avdd.t567 avdd.t565 102.091
R1303 avdd.t282 avdd.t284 102.091
R1304 avdd.t256 avdd.t254 102.091
R1305 avdd.t266 avdd.t268 102.091
R1306 avdd.t208 avdd.t210 102.091
R1307 avdd.n1320 avdd.t311 101.564
R1308 avdd.n1657 avdd.t272 101.564
R1309 avdd.n295 avdd.n294 99.0123
R1310 avdd.n300 avdd.n299 99.0123
R1311 avdd.n543 avdd.n542 99.0123
R1312 avdd.n548 avdd.n547 99.0123
R1313 avdd.n1328 avdd.t655 97.7578
R1314 avdd.n1665 avdd.t497 97.7578
R1315 avdd.n739 avdd.t278 96.8274
R1316 avdd.t584 avdd.n1744 96.5971
R1317 avdd.n695 avdd.t336 95.0005
R1318 avdd.n729 avdd.t342 95.0005
R1319 avdd.n495 avdd.n494 94.1181
R1320 avdd.n455 avdd.n454 94.1181
R1321 avdd.n919 avdd.n918 94.1181
R1322 avdd.n879 avdd.n878 94.1181
R1323 avdd.n344 avdd.n339 91.1064
R1324 avdd.n592 avdd.n587 91.1064
R1325 avdd.t388 avdd.t584 88.8801
R1326 avdd.n7 avdd.n4 86.068
R1327 avdd.n1147 avdd.n1139 86.068
R1328 avdd.n1150 avdd.n1149 86.068
R1329 avdd.n1152 avdd.n1146 86.068
R1330 avdd.n1148 avdd.n1147 86.068
R1331 avdd.n1150 avdd.n1145 86.068
R1332 avdd.n1126 avdd.n1118 86.068
R1333 avdd.n1129 avdd.n1128 86.068
R1334 avdd.n1131 avdd.n1125 86.068
R1335 avdd.n1127 avdd.n1126 86.068
R1336 avdd.n1129 avdd.n1124 86.068
R1337 avdd.n1105 avdd.n1097 86.068
R1338 avdd.n1108 avdd.n1107 86.068
R1339 avdd.n1110 avdd.n1104 86.068
R1340 avdd.n1106 avdd.n1105 86.068
R1341 avdd.n1108 avdd.n1103 86.068
R1342 avdd.n1084 avdd.n1076 86.068
R1343 avdd.n1087 avdd.n1086 86.068
R1344 avdd.n1089 avdd.n1083 86.068
R1345 avdd.n1085 avdd.n1084 86.068
R1346 avdd.n1087 avdd.n1082 86.068
R1347 avdd.n1063 avdd.n1055 86.068
R1348 avdd.n1066 avdd.n1065 86.068
R1349 avdd.n1068 avdd.n1062 86.068
R1350 avdd.n1064 avdd.n1063 86.068
R1351 avdd.n1066 avdd.n1061 86.068
R1352 avdd.n1042 avdd.n1034 86.068
R1353 avdd.n1045 avdd.n1044 86.068
R1354 avdd.n1047 avdd.n1041 86.068
R1355 avdd.n1043 avdd.n1042 86.068
R1356 avdd.n1045 avdd.n1040 86.068
R1357 avdd.n1021 avdd.n1013 86.068
R1358 avdd.n1024 avdd.n1023 86.068
R1359 avdd.n1026 avdd.n1020 86.068
R1360 avdd.n1022 avdd.n1021 86.068
R1361 avdd.n1024 avdd.n1019 86.068
R1362 avdd.n1000 avdd.n992 86.068
R1363 avdd.n1003 avdd.n1002 86.068
R1364 avdd.n1005 avdd.n999 86.068
R1365 avdd.n1001 avdd.n1000 86.068
R1366 avdd.n1003 avdd.n998 86.068
R1367 avdd.n1520 avdd.n1512 86.068
R1368 avdd.n1523 avdd.n1522 86.068
R1369 avdd.n1525 avdd.n1519 86.068
R1370 avdd.n1521 avdd.n1520 86.068
R1371 avdd.n1523 avdd.n1518 86.068
R1372 avdd.n1499 avdd.n1491 86.068
R1373 avdd.n1502 avdd.n1501 86.068
R1374 avdd.n1504 avdd.n1498 86.068
R1375 avdd.n1500 avdd.n1499 86.068
R1376 avdd.n1502 avdd.n1497 86.068
R1377 avdd.n1478 avdd.n1470 86.068
R1378 avdd.n1481 avdd.n1480 86.068
R1379 avdd.n1483 avdd.n1477 86.068
R1380 avdd.n1479 avdd.n1478 86.068
R1381 avdd.n1481 avdd.n1476 86.068
R1382 avdd.n1457 avdd.n1449 86.068
R1383 avdd.n1460 avdd.n1459 86.068
R1384 avdd.n1462 avdd.n1456 86.068
R1385 avdd.n1458 avdd.n1457 86.068
R1386 avdd.n1460 avdd.n1455 86.068
R1387 avdd.n1436 avdd.n1428 86.068
R1388 avdd.n1439 avdd.n1438 86.068
R1389 avdd.n1441 avdd.n1435 86.068
R1390 avdd.n1437 avdd.n1436 86.068
R1391 avdd.n1439 avdd.n1434 86.068
R1392 avdd.n1415 avdd.n1407 86.068
R1393 avdd.n1418 avdd.n1417 86.068
R1394 avdd.n1420 avdd.n1414 86.068
R1395 avdd.n1416 avdd.n1415 86.068
R1396 avdd.n1418 avdd.n1413 86.068
R1397 avdd.n1394 avdd.n1386 86.068
R1398 avdd.n1397 avdd.n1396 86.068
R1399 avdd.n1399 avdd.n1393 86.068
R1400 avdd.n1395 avdd.n1394 86.068
R1401 avdd.n1397 avdd.n1392 86.068
R1402 avdd.n1373 avdd.n1365 86.068
R1403 avdd.n1376 avdd.n1375 86.068
R1404 avdd.n1378 avdd.n1372 86.068
R1405 avdd.n1374 avdd.n1373 86.068
R1406 avdd.n1376 avdd.n1371 86.068
R1407 avdd.n1164 avdd.n1162 86.068
R1408 avdd.n1169 avdd.n1163 86.068
R1409 avdd.n1170 avdd.n1162 86.068
R1410 avdd.n1163 avdd.n1161 86.068
R1411 avdd.n124 avdd.t507 82.3568
R1412 avdd.n777 avdd.t443 82.3568
R1413 avdd.t336 avdd.n694 80.3851
R1414 avdd.t342 avdd.n727 80.3851
R1415 avdd.n769 avdd.t278 78.5582
R1416 avdd.t613 avdd.t382 73.4459
R1417 avdd.n684 avdd.t350 73.0774
R1418 avdd.n716 avdd.t332 73.0774
R1419 avdd.t439 avdd.n1324 72.6918
R1420 avdd.t252 avdd.n1661 72.6918
R1421 avdd.n294 avdd.n282 71.5299
R1422 avdd.n301 avdd.n300 71.5299
R1423 avdd.n542 avdd.n530 71.5299
R1424 avdd.n549 avdd.n548 71.5299
R1425 avdd.t617 avdd.n1765 69.9865
R1426 avdd.n124 avdd.n117 68.6629
R1427 avdd.n667 avdd.n666 68.6629
R1428 avdd.n777 avdd.n621 68.6629
R1429 avdd.n1771 avdd.t570 59.3422
R1430 avdd.t348 avdd.n673 58.462
R1431 avdd.t346 avdd.n706 58.462
R1432 avdd.t161 avdd.t611 58.0117
R1433 avdd.n1859 avdd.t226 55.4795
R1434 avdd.t224 avdd.n1859 55.4795
R1435 avdd.n1851 avdd.t247 54.6604
R1436 avdd.n1834 avdd.t219 54.6604
R1437 avdd.n1754 avdd.t585 53.8832
R1438 avdd.n1748 avdd.t618 53.8832
R1439 avdd.n1747 avdd.t580 53.8832
R1440 avdd.t352 avdd.n662 51.1543
R1441 avdd.n705 avdd.t324 51.1543
R1442 avdd.n1732 avdd.n1731 50.4475
R1443 avdd.n1794 avdd.t23 49.5908
R1444 avdd.n1778 avdd.t23 49.5908
R1445 avdd.n7 avdd.n6 49.4675
R1446 avdd.n1151 avdd.n1147 49.4675
R1447 avdd.n1151 avdd.n1150 49.4675
R1448 avdd.n1152 avdd.n1151 49.4675
R1449 avdd.n1130 avdd.n1126 49.4675
R1450 avdd.n1130 avdd.n1129 49.4675
R1451 avdd.n1131 avdd.n1130 49.4675
R1452 avdd.n1109 avdd.n1105 49.4675
R1453 avdd.n1109 avdd.n1108 49.4675
R1454 avdd.n1110 avdd.n1109 49.4675
R1455 avdd.n1088 avdd.n1084 49.4675
R1456 avdd.n1088 avdd.n1087 49.4675
R1457 avdd.n1089 avdd.n1088 49.4675
R1458 avdd.n1067 avdd.n1063 49.4675
R1459 avdd.n1067 avdd.n1066 49.4675
R1460 avdd.n1068 avdd.n1067 49.4675
R1461 avdd.n1046 avdd.n1042 49.4675
R1462 avdd.n1046 avdd.n1045 49.4675
R1463 avdd.n1047 avdd.n1046 49.4675
R1464 avdd.n1025 avdd.n1021 49.4675
R1465 avdd.n1025 avdd.n1024 49.4675
R1466 avdd.n1026 avdd.n1025 49.4675
R1467 avdd.n1004 avdd.n1000 49.4675
R1468 avdd.n1004 avdd.n1003 49.4675
R1469 avdd.n1005 avdd.n1004 49.4675
R1470 avdd.n1524 avdd.n1520 49.4675
R1471 avdd.n1524 avdd.n1523 49.4675
R1472 avdd.n1525 avdd.n1524 49.4675
R1473 avdd.n1503 avdd.n1499 49.4675
R1474 avdd.n1503 avdd.n1502 49.4675
R1475 avdd.n1504 avdd.n1503 49.4675
R1476 avdd.n1482 avdd.n1478 49.4675
R1477 avdd.n1482 avdd.n1481 49.4675
R1478 avdd.n1483 avdd.n1482 49.4675
R1479 avdd.n1461 avdd.n1457 49.4675
R1480 avdd.n1461 avdd.n1460 49.4675
R1481 avdd.n1462 avdd.n1461 49.4675
R1482 avdd.n1440 avdd.n1436 49.4675
R1483 avdd.n1440 avdd.n1439 49.4675
R1484 avdd.n1441 avdd.n1440 49.4675
R1485 avdd.n1419 avdd.n1415 49.4675
R1486 avdd.n1419 avdd.n1418 49.4675
R1487 avdd.n1420 avdd.n1419 49.4675
R1488 avdd.n1398 avdd.n1394 49.4675
R1489 avdd.n1398 avdd.n1397 49.4675
R1490 avdd.n1399 avdd.n1398 49.4675
R1491 avdd.n1377 avdd.n1373 49.4675
R1492 avdd.n1377 avdd.n1376 49.4675
R1493 avdd.n1378 avdd.n1377 49.4675
R1494 avdd.n1181 avdd.n1162 49.4675
R1495 avdd.n1181 avdd.n1163 49.4675
R1496 avdd.n1850 avdd.n1849 49.1214
R1497 avdd.n1848 avdd.n1847 49.1214
R1498 avdd.n1846 avdd.n1845 49.1214
R1499 avdd.n1844 avdd.n1843 49.1214
R1500 avdd.n1842 avdd.n1841 49.1214
R1501 avdd.n1840 avdd.n1839 49.1214
R1502 avdd.n1838 avdd.n1837 49.1214
R1503 avdd.t577 avdd.t382 48.4319
R1504 avdd.n1756 avdd.n1755 48.3442
R1505 avdd.n1758 avdd.n1757 48.3442
R1506 avdd.n1783 avdd.n1782 48.2034
R1507 avdd.n1785 avdd.n1784 48.2034
R1508 avdd.n1791 avdd.n1790 48.2034
R1509 avdd.n1798 avdd.n1797 48.2034
R1510 avdd.n1800 avdd.n1799 48.2034
R1511 avdd.n1802 avdd.n1801 48.2034
R1512 avdd.n1804 avdd.n1803 48.2034
R1513 avdd.n1780 avdd.t46 48.0365
R1514 avdd.n1805 avdd.t162 48.0365
R1515 avdd.n1326 avdd.t439 47.6258
R1516 avdd.n1663 avdd.t252 47.6258
R1517 avdd.t571 avdd.t575 47.3674
R1518 avdd.t575 avdd.t108 47.3674
R1519 avdd.t108 avdd.t576 47.3674
R1520 avdd.t120 avdd.t576 47.3674
R1521 avdd.t176 avdd.t583 47.3674
R1522 avdd.t581 avdd.t176 47.3674
R1523 avdd.t570 avdd.t581 47.3674
R1524 avdd.n496 avdd.n495 44.8005
R1525 avdd.n456 avdd.n455 44.8005
R1526 avdd.n920 avdd.n919 44.8005
R1527 avdd.n880 avdd.n879 44.8005
R1528 avdd.n1687 avdd 43.959
R1529 avdd.n345 avdd.n340 43.2946
R1530 avdd.n593 avdd.n588 43.2946
R1531 avdd.n1744 avdd.t623 42.8436
R1532 avdd.n1787 avdd.n1786 42.4975
R1533 avdd.n1789 avdd.n1779 42.4505
R1534 avdd.n1811 avdd.t617 41.247
R1535 avdd.n1765 avdd.t161 38.5859
R1536 avdd.n299 avdd.n298 37.0005
R1537 avdd.n296 avdd.n295 37.0005
R1538 avdd.n547 avdd.n546 37.0005
R1539 avdd.n544 avdd.n543 37.0005
R1540 avdd.t328 avdd.n685 36.539
R1541 avdd.n718 avdd.t334 36.539
R1542 avdd.n1709 avdd.n1708 36.4934
R1543 avdd.n131 avdd.n130 36.1417
R1544 avdd.n130 avdd.n125 36.1417
R1545 avdd.n138 avdd.n115 36.1417
R1546 avdd.n118 avdd.n115 36.1417
R1547 avdd.n149 avdd.n107 36.1417
R1548 avdd.n143 avdd.n107 36.1417
R1549 avdd.n156 avdd.n155 36.1417
R1550 avdd.n155 avdd.n104 36.1417
R1551 avdd.n163 avdd.n95 36.1417
R1552 avdd.n98 avdd.n95 36.1417
R1553 avdd.n174 avdd.n87 36.1417
R1554 avdd.n168 avdd.n87 36.1417
R1555 avdd.n181 avdd.n180 36.1417
R1556 avdd.n180 avdd.n84 36.1417
R1557 avdd.n188 avdd.n75 36.1417
R1558 avdd.n78 avdd.n75 36.1417
R1559 avdd.n199 avdd.n67 36.1417
R1560 avdd.n193 avdd.n67 36.1417
R1561 avdd.n206 avdd.n205 36.1417
R1562 avdd.n205 avdd.n64 36.1417
R1563 avdd.n213 avdd.n55 36.1417
R1564 avdd.n58 avdd.n55 36.1417
R1565 avdd.n224 avdd.n47 36.1417
R1566 avdd.n218 avdd.n47 36.1417
R1567 avdd.n231 avdd.n230 36.1417
R1568 avdd.n230 avdd.n44 36.1417
R1569 avdd.n238 avdd.n35 36.1417
R1570 avdd.n38 avdd.n35 36.1417
R1571 avdd.n249 avdd.n28 36.1417
R1572 avdd.n243 avdd.n28 36.1417
R1573 avdd.n256 avdd.n255 36.1417
R1574 avdd.n255 avdd.n254 36.1417
R1575 avdd.n9 avdd.n3 36.1417
R1576 avdd.n9 avdd.n8 36.1417
R1577 avdd.n1208 avdd.n1207 36.1417
R1578 avdd.n1207 avdd.n1140 36.1417
R1579 avdd.n1144 avdd.n1140 36.1417
R1580 avdd.n1200 avdd.n1144 36.1417
R1581 avdd.n1200 avdd.n1199 36.1417
R1582 avdd.n1199 avdd.n1153 36.1417
R1583 avdd.n1223 avdd.n1222 36.1417
R1584 avdd.n1222 avdd.n1119 36.1417
R1585 avdd.n1123 avdd.n1119 36.1417
R1586 avdd.n1215 avdd.n1123 36.1417
R1587 avdd.n1215 avdd.n1214 36.1417
R1588 avdd.n1214 avdd.n1132 36.1417
R1589 avdd.n1238 avdd.n1237 36.1417
R1590 avdd.n1237 avdd.n1098 36.1417
R1591 avdd.n1102 avdd.n1098 36.1417
R1592 avdd.n1230 avdd.n1102 36.1417
R1593 avdd.n1230 avdd.n1229 36.1417
R1594 avdd.n1229 avdd.n1111 36.1417
R1595 avdd.n1253 avdd.n1252 36.1417
R1596 avdd.n1252 avdd.n1077 36.1417
R1597 avdd.n1081 avdd.n1077 36.1417
R1598 avdd.n1245 avdd.n1081 36.1417
R1599 avdd.n1245 avdd.n1244 36.1417
R1600 avdd.n1244 avdd.n1090 36.1417
R1601 avdd.n1268 avdd.n1267 36.1417
R1602 avdd.n1267 avdd.n1056 36.1417
R1603 avdd.n1060 avdd.n1056 36.1417
R1604 avdd.n1260 avdd.n1060 36.1417
R1605 avdd.n1260 avdd.n1259 36.1417
R1606 avdd.n1259 avdd.n1069 36.1417
R1607 avdd.n1283 avdd.n1282 36.1417
R1608 avdd.n1282 avdd.n1035 36.1417
R1609 avdd.n1039 avdd.n1035 36.1417
R1610 avdd.n1275 avdd.n1039 36.1417
R1611 avdd.n1275 avdd.n1274 36.1417
R1612 avdd.n1274 avdd.n1048 36.1417
R1613 avdd.n1298 avdd.n1297 36.1417
R1614 avdd.n1297 avdd.n1014 36.1417
R1615 avdd.n1018 avdd.n1014 36.1417
R1616 avdd.n1290 avdd.n1018 36.1417
R1617 avdd.n1290 avdd.n1289 36.1417
R1618 avdd.n1289 avdd.n1027 36.1417
R1619 avdd.n1313 avdd.n1312 36.1417
R1620 avdd.n1312 avdd.n993 36.1417
R1621 avdd.n997 avdd.n993 36.1417
R1622 avdd.n1305 avdd.n997 36.1417
R1623 avdd.n1305 avdd.n1304 36.1417
R1624 avdd.n1304 avdd.n1006 36.1417
R1625 avdd.n1348 avdd.n1347 36.1417
R1626 avdd.n1347 avdd.n981 36.1417
R1627 avdd.n1343 avdd.n981 36.1417
R1628 avdd.n1343 avdd.n1342 36.1417
R1629 avdd.n1342 avdd.n988 36.1417
R1630 avdd.n1318 avdd.n988 36.1417
R1631 avdd.n1330 avdd.n1318 36.1417
R1632 avdd.n1545 avdd.n1544 36.1417
R1633 avdd.n1544 avdd.n1513 36.1417
R1634 avdd.n1517 avdd.n1513 36.1417
R1635 avdd.n1537 avdd.n1517 36.1417
R1636 avdd.n1537 avdd.n1536 36.1417
R1637 avdd.n1536 avdd.n1526 36.1417
R1638 avdd.n1560 avdd.n1559 36.1417
R1639 avdd.n1559 avdd.n1492 36.1417
R1640 avdd.n1496 avdd.n1492 36.1417
R1641 avdd.n1552 avdd.n1496 36.1417
R1642 avdd.n1552 avdd.n1551 36.1417
R1643 avdd.n1551 avdd.n1505 36.1417
R1644 avdd.n1575 avdd.n1574 36.1417
R1645 avdd.n1574 avdd.n1471 36.1417
R1646 avdd.n1475 avdd.n1471 36.1417
R1647 avdd.n1567 avdd.n1475 36.1417
R1648 avdd.n1567 avdd.n1566 36.1417
R1649 avdd.n1566 avdd.n1484 36.1417
R1650 avdd.n1590 avdd.n1589 36.1417
R1651 avdd.n1589 avdd.n1450 36.1417
R1652 avdd.n1454 avdd.n1450 36.1417
R1653 avdd.n1582 avdd.n1454 36.1417
R1654 avdd.n1582 avdd.n1581 36.1417
R1655 avdd.n1581 avdd.n1463 36.1417
R1656 avdd.n1605 avdd.n1604 36.1417
R1657 avdd.n1604 avdd.n1429 36.1417
R1658 avdd.n1433 avdd.n1429 36.1417
R1659 avdd.n1597 avdd.n1433 36.1417
R1660 avdd.n1597 avdd.n1596 36.1417
R1661 avdd.n1596 avdd.n1442 36.1417
R1662 avdd.n1620 avdd.n1619 36.1417
R1663 avdd.n1619 avdd.n1408 36.1417
R1664 avdd.n1412 avdd.n1408 36.1417
R1665 avdd.n1612 avdd.n1412 36.1417
R1666 avdd.n1612 avdd.n1611 36.1417
R1667 avdd.n1611 avdd.n1421 36.1417
R1668 avdd.n1635 avdd.n1634 36.1417
R1669 avdd.n1634 avdd.n1387 36.1417
R1670 avdd.n1391 avdd.n1387 36.1417
R1671 avdd.n1627 avdd.n1391 36.1417
R1672 avdd.n1627 avdd.n1626 36.1417
R1673 avdd.n1626 avdd.n1400 36.1417
R1674 avdd.n1650 avdd.n1649 36.1417
R1675 avdd.n1649 avdd.n1366 36.1417
R1676 avdd.n1370 avdd.n1366 36.1417
R1677 avdd.n1642 avdd.n1370 36.1417
R1678 avdd.n1642 avdd.n1641 36.1417
R1679 avdd.n1641 avdd.n1379 36.1417
R1680 avdd.n1685 avdd.n1684 36.1417
R1681 avdd.n1680 avdd.n1354 36.1417
R1682 avdd.n1680 avdd.n1679 36.1417
R1683 avdd.n1679 avdd.n1361 36.1417
R1684 avdd.n1655 avdd.n1361 36.1417
R1685 avdd.n1667 avdd.n1655 36.1417
R1686 avdd.n1179 avdd.n1165 36.1417
R1687 avdd.n1171 avdd.n1165 36.1417
R1688 avdd.n1171 avdd.n1160 36.1417
R1689 avdd.n1184 avdd.n1160 36.1417
R1690 avdd.n1184 avdd.n1183 36.1417
R1691 avdd.n665 avdd.n664 36.1417
R1692 avdd.n671 avdd.n664 36.1417
R1693 avdd.n671 avdd.n660 36.1417
R1694 avdd.n678 avdd.n660 36.1417
R1695 avdd.n678 avdd.n658 36.1417
R1696 avdd.n682 avdd.n658 36.1417
R1697 avdd.n682 avdd.n655 36.1417
R1698 avdd.n688 avdd.n655 36.1417
R1699 avdd.n688 avdd.n653 36.1417
R1700 avdd.n692 avdd.n653 36.1417
R1701 avdd.n692 avdd.n649 36.1417
R1702 avdd.n699 avdd.n649 36.1417
R1703 avdd.n699 avdd.n647 36.1417
R1704 avdd.n703 avdd.n647 36.1417
R1705 avdd.n703 avdd.n644 36.1417
R1706 avdd.n709 avdd.n644 36.1417
R1707 avdd.n709 avdd.n642 36.1417
R1708 avdd.n713 avdd.n642 36.1417
R1709 avdd.n713 avdd.n638 36.1417
R1710 avdd.n720 avdd.n638 36.1417
R1711 avdd.n720 avdd.n636 36.1417
R1712 avdd.n724 avdd.n636 36.1417
R1713 avdd.n724 avdd.n633 36.1417
R1714 avdd.n731 avdd.n633 36.1417
R1715 avdd.n731 avdd.n631 36.1417
R1716 avdd.n735 avdd.n631 36.1417
R1717 avdd.n735 avdd.n628 36.1417
R1718 avdd.n742 avdd.n628 36.1417
R1719 avdd.n742 avdd.n625 36.1417
R1720 avdd.n767 avdd.n625 36.1417
R1721 avdd.n767 avdd.n626 36.1417
R1722 avdd.n626 avdd.n623 36.1417
R1723 avdd.n623 avdd.n617 36.1417
R1724 avdd.n783 avdd.n617 36.1417
R1725 avdd.n783 avdd.n782 36.1417
R1726 avdd.n782 avdd.n620 36.1417
R1727 avdd.n778 avdd.n620 36.1417
R1728 avdd.n1684 avdd.n1354 35.7652
R1729 avdd.n774 avdd.t274 34.712
R1730 avdd.t603 avdd.t388 32.9977
R1731 avdd.n1752 avdd.n1740 31.624
R1732 avdd.n1763 avdd.n1760 31.624
R1733 avdd.n1828 avdd.n1735 31.624
R1734 avdd.n445 avdd.n367 31.2476
R1735 avdd.n365 avdd.n364 31.2476
R1736 avdd.n869 avdd.n615 31.2476
R1737 avdd.n613 avdd.n612 31.2476
R1738 avdd.n1708 avdd.n959 31.2285
R1739 avdd.t276 avdd.n770 31.0582
R1740 avdd.n454 avdd.n453 30.8338
R1741 avdd.n453 avdd.n452 30.8338
R1742 avdd.n494 avdd.n493 30.8338
R1743 avdd.n493 avdd.n492 30.8338
R1744 avdd.n367 avdd.n363 30.8338
R1745 avdd.n365 avdd.n362 30.8338
R1746 avdd.n878 avdd.n877 30.8338
R1747 avdd.n877 avdd.n876 30.8338
R1748 avdd.n918 avdd.n917 30.8338
R1749 avdd.n917 avdd.n916 30.8338
R1750 avdd.n615 avdd.n611 30.8338
R1751 avdd.n613 avdd.n610 30.8338
R1752 avdd.n968 avdd.n966 30.3029
R1753 avdd.t330 avdd.n651 29.2313
R1754 avdd.n726 avdd.t340 29.2313
R1755 avdd.n1714 avdd.n1709 27.9872
R1756 avdd.n386 avdd.t361 27.6955
R1757 avdd.n386 avdd.t207 27.6955
R1758 avdd.n384 avdd.t359 27.6955
R1759 avdd.n384 avdd.t201 27.6955
R1760 avdd.n382 avdd.t358 27.6955
R1761 avdd.n382 avdd.t198 27.6955
R1762 avdd.n380 avdd.t355 27.6955
R1763 avdd.n380 avdd.t196 27.6955
R1764 avdd.n378 avdd.t186 27.6955
R1765 avdd.n378 avdd.t363 27.6955
R1766 avdd.n376 avdd.t183 27.6955
R1767 avdd.n376 avdd.t365 27.6955
R1768 avdd.n374 avdd.t185 27.6955
R1769 avdd.n374 avdd.t364 27.6955
R1770 avdd.n372 avdd.t202 27.6955
R1771 avdd.n372 avdd.t373 27.6955
R1772 avdd.n370 avdd.t206 27.6955
R1773 avdd.n370 avdd.t368 27.6955
R1774 avdd.n368 avdd.t189 27.6955
R1775 avdd.n368 avdd.t374 27.6955
R1776 avdd.n307 avdd.t187 27.6955
R1777 avdd.n307 avdd.t375 27.6955
R1778 avdd.n481 avdd.t199 27.6955
R1779 avdd.n481 avdd.t362 27.6955
R1780 avdd.t128 avdd.n430 27.6955
R1781 avdd.n430 avdd.t360 27.6955
R1782 avdd.n427 avdd.t85 27.6955
R1783 avdd.n427 avdd.t357 27.6955
R1784 avdd.n424 avdd.t78 27.6955
R1785 avdd.n424 avdd.t356 27.6955
R1786 avdd.t60 avdd.n419 27.6955
R1787 avdd.n419 avdd.t354 27.6955
R1788 avdd.t62 avdd.n416 27.6955
R1789 avdd.n416 avdd.t184 27.6955
R1790 avdd.n413 avdd.t48 27.6955
R1791 avdd.n413 avdd.t205 27.6955
R1792 avdd.n410 avdd.t55 27.6955
R1793 avdd.n410 avdd.t181 27.6955
R1794 avdd.t14 avdd.n405 27.6955
R1795 avdd.n405 avdd.t197 27.6955
R1796 avdd.t42 avdd.n402 27.6955
R1797 avdd.n402 avdd.t204 27.6955
R1798 avdd.n399 avdd.t147 27.6955
R1799 avdd.n399 avdd.t190 27.6955
R1800 avdd.n396 avdd.t145 27.6955
R1801 avdd.n396 avdd.t188 27.6955
R1802 avdd.n460 avdd.t69 27.6955
R1803 avdd.n460 avdd.t200 27.6955
R1804 avdd.n312 avdd.t203 27.6955
R1805 avdd.n312 avdd.t57 27.6955
R1806 avdd.n314 avdd.t194 27.6955
R1807 avdd.n314 avdd.t21 27.6955
R1808 avdd.n316 avdd.t193 27.6955
R1809 avdd.n316 avdd.t18 27.6955
R1810 avdd.n318 avdd.t192 27.6955
R1811 avdd.n318 avdd.t7 27.6955
R1812 avdd.n320 avdd.t369 27.6955
R1813 avdd.n320 avdd.t10 27.6955
R1814 avdd.n322 avdd.t371 27.6955
R1815 avdd.n322 avdd.t173 27.6955
R1816 avdd.n324 avdd.t370 27.6955
R1817 avdd.n324 avdd.t4 27.6955
R1818 avdd.n326 avdd.t377 27.6955
R1819 avdd.n326 avdd.t122 27.6955
R1820 avdd.n328 avdd.t372 27.6955
R1821 avdd.n328 avdd.t166 27.6955
R1822 avdd.n330 avdd.t366 27.6955
R1823 avdd.n330 avdd.t133 27.6955
R1824 avdd.n332 avdd.t367 27.6955
R1825 avdd.n332 avdd.t125 27.6955
R1826 avdd.n335 avdd.t376 27.6955
R1827 avdd.n335 avdd.t50 27.6955
R1828 avdd.n436 avdd.t492 27.6955
R1829 avdd.n436 avdd.t488 27.6955
R1830 avdd.n438 avdd.t486 27.6955
R1831 avdd.n438 avdd.t478 27.6955
R1832 avdd.n440 avdd.t490 27.6955
R1833 avdd.n440 avdd.t484 27.6955
R1834 avdd.n442 avdd.t480 27.6955
R1835 avdd.n442 avdd.t502 27.6955
R1836 avdd.n809 avdd.t632 27.6955
R1837 avdd.n809 avdd.t399 27.6955
R1838 avdd.n807 avdd.t628 27.6955
R1839 avdd.n807 avdd.t394 27.6955
R1840 avdd.n805 avdd.t631 27.6955
R1841 avdd.n805 avdd.t398 27.6955
R1842 avdd.n803 avdd.t627 27.6955
R1843 avdd.n803 avdd.t393 27.6955
R1844 avdd.n801 avdd.t404 27.6955
R1845 avdd.n801 avdd.t640 27.6955
R1846 avdd.n799 avdd.t411 27.6955
R1847 avdd.n799 avdd.t644 27.6955
R1848 avdd.n797 avdd.t412 27.6955
R1849 avdd.n797 avdd.t645 27.6955
R1850 avdd.n795 avdd.t413 27.6955
R1851 avdd.n795 avdd.t646 27.6955
R1852 avdd.n793 avdd.t414 27.6955
R1853 avdd.n793 avdd.t647 27.6955
R1854 avdd.n791 avdd.t417 27.6955
R1855 avdd.n791 avdd.t638 27.6955
R1856 avdd.n555 avdd.t415 27.6955
R1857 avdd.n555 avdd.t648 27.6955
R1858 avdd.n905 avdd.t405 27.6955
R1859 avdd.n905 avdd.t641 27.6955
R1860 avdd.t159 avdd.n853 27.6955
R1861 avdd.n853 avdd.t626 27.6955
R1862 avdd.n850 avdd.t113 27.6955
R1863 avdd.n850 avdd.t630 27.6955
R1864 avdd.n847 avdd.t152 27.6955
R1865 avdd.n847 avdd.t625 27.6955
R1866 avdd.t104 avdd.n842 27.6955
R1867 avdd.n842 avdd.t629 27.6955
R1868 avdd.t143 avdd.n839 27.6955
R1869 avdd.n839 avdd.t418 27.6955
R1870 avdd.n836 avdd.t97 27.6955
R1871 avdd.n836 avdd.t406 27.6955
R1872 avdd.n833 avdd.t95 27.6955
R1873 avdd.n833 avdd.t407 27.6955
R1874 avdd.t87 avdd.n828 27.6955
R1875 avdd.n828 avdd.t408 27.6955
R1876 avdd.t83 avdd.n825 27.6955
R1877 avdd.n825 avdd.t409 27.6955
R1878 avdd.n822 avdd.t34 27.6955
R1879 avdd.n822 avdd.t416 27.6955
R1880 avdd.n819 avdd.t71 27.6955
R1881 avdd.n819 avdd.t410 27.6955
R1882 avdd.n884 avdd.t136 27.6955
R1883 avdd.n884 avdd.t402 27.6955
R1884 avdd.n560 avdd.t397 27.6955
R1885 avdd.n560 avdd.t154 27.6955
R1886 avdd.n562 avdd.t455 27.6955
R1887 avdd.n562 avdd.t110 27.6955
R1888 avdd.n564 avdd.t396 27.6955
R1889 avdd.n564 avdd.t149 27.6955
R1890 avdd.n566 avdd.t400 27.6955
R1891 avdd.n566 avdd.t101 27.6955
R1892 avdd.n568 avdd.t642 27.6955
R1893 avdd.n568 avdd.t138 27.6955
R1894 avdd.n570 avdd.t633 27.6955
R1895 avdd.n570 avdd.t92 27.6955
R1896 avdd.n572 avdd.t634 27.6955
R1897 avdd.n572 avdd.t89 27.6955
R1898 avdd.n574 avdd.t635 27.6955
R1899 avdd.n574 avdd.t80 27.6955
R1900 avdd.n576 avdd.t636 27.6955
R1901 avdd.n576 avdd.t75 27.6955
R1902 avdd.n578 avdd.t639 27.6955
R1903 avdd.n578 avdd.t28 27.6955
R1904 avdd.n580 avdd.t637 27.6955
R1905 avdd.n580 avdd.t64 27.6955
R1906 avdd.n583 avdd.t643 27.6955
R1907 avdd.n583 avdd.t130 27.6955
R1908 avdd.n860 avdd.t533 27.6955
R1909 avdd.n860 avdd.t529 27.6955
R1910 avdd.n862 avdd.t539 27.6955
R1911 avdd.n862 avdd.t537 27.6955
R1912 avdd.n864 avdd.t531 27.6955
R1913 avdd.n864 avdd.t543 27.6955
R1914 avdd.n866 avdd.t535 27.6955
R1915 avdd.n866 avdd.t547 27.6955
R1916 avdd.t36 avdd.n1811 26.7523
R1917 avdd.n1780 avdd.t43 25.5567
R1918 avdd.n1805 avdd.t160 25.5567
R1919 avdd.n1787 avdd.t114 25.4942
R1920 avdd.t583 avdd.t621 25.0145
R1921 avdd.n1695 avdd.n1694 24.9671
R1922 avdd.n1141 avdd.t299 23.5572
R1923 avdd.n1120 avdd.t514 23.5572
R1924 avdd.n1099 avdd.t303 23.5572
R1925 avdd.n1078 avdd.t318 23.5572
R1926 avdd.n1057 avdd.t420 23.5572
R1927 avdd.n1036 avdd.t587 23.5572
R1928 avdd.n1015 avdd.t287 23.5572
R1929 avdd.n994 avdd.t306 23.5572
R1930 avdd.n1336 avdd.t440 23.5572
R1931 avdd.n1514 avdd.t509 23.5572
R1932 avdd.n1493 avdd.t597 23.5572
R1933 avdd.n1472 avdd.t562 23.5572
R1934 avdd.n1451 avdd.t566 23.5572
R1935 avdd.n1430 avdd.t285 23.5572
R1936 avdd.n1409 avdd.t255 23.5572
R1937 avdd.n1388 avdd.t269 23.5572
R1938 avdd.n1367 avdd.t211 23.5572
R1939 avdd.n1673 avdd.t253 23.5572
R1940 avdd.n1167 avdd.t659 23.5572
R1941 avdd.t120 avdd.t621 22.3534
R1942 avdd.n1713 avdd.n1710 21.9177
R1943 avdd.n1725 avdd.n1724 20.3986
R1944 avdd.n1724 avdd.n949 20.2792
R1945 avdd.n978 avdd 20.0949
R1946 avdd.n968 avdd.n948 19.4414
R1947 avdd.n1700 avdd.n1699 18.824
R1948 avdd.n984 avdd 18.3657
R1949 avdd.n1357 avdd 18.3657
R1950 avdd.n1141 avdd.t493 17.8272
R1951 avdd.n1120 avdd.t454 17.8272
R1952 avdd.n1099 avdd.t496 17.8272
R1953 avdd.n1078 avdd.t319 17.8272
R1954 avdd.n1057 avdd.t517 17.8272
R1955 avdd.n1036 avdd.t557 17.8272
R1956 avdd.n1015 avdd.t291 17.8272
R1957 avdd.n994 avdd.t293 17.8272
R1958 avdd.n1336 avdd.t295 17.8272
R1959 avdd.n1514 avdd.t310 17.8272
R1960 avdd.n1493 avdd.t650 17.8272
R1961 avdd.n1472 avdd.t314 17.8272
R1962 avdd.n1451 avdd.t569 17.8272
R1963 avdd.n1430 avdd.t649 17.8272
R1964 avdd.n1409 avdd.t463 17.8272
R1965 avdd.n1388 avdd.t586 17.8272
R1966 avdd.n1367 avdd.t602 17.8272
R1967 avdd.n1673 avdd.t448 17.8272
R1968 avdd.n1167 avdd.t446 17.8272
R1969 avdd.n745 avdd.t341 17.8272
R1970 avdd.n745 avdd.t343 17.8272
R1971 avdd.n746 avdd.t333 17.8272
R1972 avdd.n746 avdd.t335 17.8272
R1973 avdd.n747 avdd.t347 17.8272
R1974 avdd.n747 avdd.t327 17.8272
R1975 avdd.n748 avdd.t339 17.8272
R1976 avdd.n748 avdd.t325 17.8272
R1977 avdd.n749 avdd.t331 17.8272
R1978 avdd.n749 avdd.t337 17.8272
R1979 avdd.n750 avdd.t351 17.8272
R1980 avdd.n750 avdd.t329 17.8272
R1981 avdd.n751 avdd.t349 17.8272
R1982 avdd.n751 avdd.t323 17.8272
R1983 avdd.n761 avdd.t279 17.8272
R1984 avdd.n761 avdd.t277 17.8272
R1985 avdd.n452 avdd.n448 17.7802
R1986 avdd.n492 avdd.n287 17.7802
R1987 avdd.n876 avdd.n872 17.7802
R1988 avdd.n916 avdd.n535 17.7802
R1989 avdd.n1196 avdd.n1195 17.7258
R1990 avdd.n1211 avdd.n1210 17.7258
R1991 avdd.n1226 avdd.n1225 17.7258
R1992 avdd.n1241 avdd.n1240 17.7258
R1993 avdd.n1256 avdd.n1255 17.7258
R1994 avdd.n1271 avdd.n1270 17.7258
R1995 avdd.n1286 avdd.n1285 17.7258
R1996 avdd.n1301 avdd.n1300 17.7258
R1997 avdd.n1317 avdd.n1316 17.7258
R1998 avdd.n1533 avdd.n1532 17.7258
R1999 avdd.n1548 avdd.n1547 17.7258
R2000 avdd.n1563 avdd.n1562 17.7258
R2001 avdd.n1578 avdd.n1577 17.7258
R2002 avdd.n1593 avdd.n1592 17.7258
R2003 avdd.n1608 avdd.n1607 17.7258
R2004 avdd.n1623 avdd.n1622 17.7258
R2005 avdd.n1638 avdd.n1637 17.7258
R2006 avdd.n1654 avdd.n1653 17.7258
R2007 avdd.n1192 avdd.n1191 17.7258
R2008 avdd.n984 avdd.n983 17.3701
R2009 avdd.n983 avdd.n982 17.3701
R2010 avdd.n1357 avdd.n1356 17.3701
R2011 avdd.n1356 avdd.n1355 17.3701
R2012 avdd.n1807 avdd.n1770 16.6169
R2013 avdd.t623 avdd.t571 16.4991
R2014 avdd.n1807 avdd.n1796 16.3798
R2015 avdd.n1753 avdd.n1752 14.9605
R2016 avdd.n1760 avdd.n1759 14.9605
R2017 avdd.n1194 avdd.n1193 14.7017
R2018 avdd.n965 avdd.n960 14.6829
R2019 avdd.n1777 avdd.n1776 14.6449
R2020 avdd.n697 avdd.t338 14.6159
R2021 avdd.n728 avdd.t344 14.6159
R2022 avdd.n279 avdd.t49 14.6083
R2023 avdd.n459 avdd.t68 14.6083
R2024 avdd.n527 avdd.t129 14.6083
R2025 avdd.n883 avdd.t135 14.6083
R2026 avdd.n1714 avdd.n1713 14.4431
R2027 avdd.n510 avdd.t9 14.4262
R2028 avdd.n508 avdd.t172 14.4262
R2029 avdd.n506 avdd.t2 14.4262
R2030 avdd.n504 avdd.t121 14.4262
R2031 avdd.n502 avdd.t165 14.4262
R2032 avdd.n500 avdd.t132 14.4262
R2033 avdd.n498 avdd.t124 14.4262
R2034 avdd.n417 avdd.t61 14.4262
R2035 avdd.n412 avdd.t47 14.4262
R2036 avdd.n409 avdd.t54 14.4262
R2037 avdd.n406 avdd.t12 14.4262
R2038 avdd.n403 avdd.t41 14.4262
R2039 avdd.n398 avdd.t146 14.4262
R2040 avdd.n395 avdd.t144 14.4262
R2041 avdd.n934 avdd.t137 14.4262
R2042 avdd.n932 avdd.t91 14.4262
R2043 avdd.n930 avdd.t88 14.4262
R2044 avdd.n928 avdd.t79 14.4262
R2045 avdd.n926 avdd.t74 14.4262
R2046 avdd.n924 avdd.t26 14.4262
R2047 avdd.n922 avdd.t63 14.4262
R2048 avdd.n840 avdd.t142 14.4262
R2049 avdd.n835 avdd.t96 14.4262
R2050 avdd.n832 avdd.t94 14.4262
R2051 avdd.n829 avdd.t86 14.4262
R2052 avdd.n826 avdd.t82 14.4262
R2053 avdd.n821 avdd.t32 14.4262
R2054 avdd.n818 avdd.t70 14.4262
R2055 avdd.n518 avdd.t56 14.4191
R2056 avdd.n516 avdd.t20 14.4191
R2057 avdd.n514 avdd.t17 14.4191
R2058 avdd.n512 avdd.t6 14.4191
R2059 avdd.n431 avdd.t127 14.4191
R2060 avdd.n426 avdd.t84 14.4191
R2061 avdd.n423 avdd.t77 14.4191
R2062 avdd.n420 avdd.t59 14.4191
R2063 avdd.n942 avdd.t153 14.4191
R2064 avdd.n940 avdd.t109 14.4191
R2065 avdd.n938 avdd.t148 14.4191
R2066 avdd.n936 avdd.t100 14.4191
R2067 avdd.n854 avdd.t158 14.4191
R2068 avdd.n849 avdd.t112 14.4191
R2069 avdd.n846 avdd.t151 14.4191
R2070 avdd.n843 avdd.t103 14.4191
R2071 avdd.n1795 avdd.n1776 14.4078
R2072 avdd.n1813 avdd.n1812 14.2313
R2073 avdd.t36 avdd.n1813 14.2313
R2074 avdd.n1815 avdd.n1814 14.2313
R2075 avdd.n1814 avdd.t36 14.2313
R2076 avdd.n975 avdd.n966 14.1829
R2077 avdd.n445 avdd.n444 14.0622
R2078 avdd.n869 avdd.n868 14.0622
R2079 avdd.n1698 avdd.n1697 13.9971
R2080 avdd.n1878 avdd.n1877 13.8347
R2081 avdd.n1868 avdd.n1867 13.8322
R2082 avdd.n274 avdd.n273 13.822
R2083 avdd.n1870 avdd.n275 13.822
R2084 avdd.n497 avdd.n496 13.8005
R2085 avdd.n484 avdd.n483 13.8005
R2086 avdd.n350 avdd.n306 13.8005
R2087 avdd.n334 avdd.n281 13.8005
R2088 avdd.n457 avdd.n456 13.8005
R2089 avdd.n434 avdd.n364 13.8005
R2090 avdd.n921 avdd.n920 13.8005
R2091 avdd.n908 avdd.n907 13.8005
R2092 avdd.n598 avdd.n554 13.8005
R2093 avdd.n582 avdd.n529 13.8005
R2094 avdd.n881 avdd.n880 13.8005
R2095 avdd.n858 avdd.n612 13.8005
R2096 avdd.n1323 avdd.t294 13.7868
R2097 avdd.n1660 avdd.t447 13.7868
R2098 avdd.n349 avdd.n309 13.436
R2099 avdd.n476 avdd.n337 13.436
R2100 avdd.n463 avdd.n462 13.436
R2101 avdd.n597 avdd.n557 13.436
R2102 avdd.n900 avdd.n585 13.436
R2103 avdd.n887 avdd.n886 13.436
R2104 avdd.n466 avdd.n465 13.177
R2105 avdd.n890 avdd.n889 13.177
R2106 avdd.n357 avdd.n356 13.0943
R2107 avdd.n356 avdd.n355 13.0943
R2108 avdd.n605 avdd.n604 13.0943
R2109 avdd.n604 avdd.n603 13.0943
R2110 avdd.n740 avdd.t280 12.789
R2111 avdd.n1197 avdd.n1196 12.541
R2112 avdd.n1212 avdd.n1211 12.541
R2113 avdd.n1227 avdd.n1226 12.541
R2114 avdd.n1242 avdd.n1241 12.541
R2115 avdd.n1257 avdd.n1256 12.541
R2116 avdd.n1272 avdd.n1271 12.541
R2117 avdd.n1287 avdd.n1286 12.541
R2118 avdd.n1302 avdd.n1301 12.541
R2119 avdd.n1316 avdd.n1315 12.541
R2120 avdd.n1534 avdd.n1533 12.541
R2121 avdd.n1549 avdd.n1548 12.541
R2122 avdd.n1564 avdd.n1563 12.541
R2123 avdd.n1579 avdd.n1578 12.541
R2124 avdd.n1594 avdd.n1593 12.541
R2125 avdd.n1609 avdd.n1608 12.541
R2126 avdd.n1624 avdd.n1623 12.541
R2127 avdd.n1639 avdd.n1638 12.541
R2128 avdd.n1653 avdd.n1652 12.541
R2129 avdd.n1191 avdd.n1190 12.541
R2130 avdd.n1153 avdd 12.424
R2131 avdd.n1132 avdd 12.424
R2132 avdd.n1111 avdd 12.424
R2133 avdd.n1090 avdd 12.424
R2134 avdd.n1069 avdd 12.424
R2135 avdd.n1048 avdd 12.424
R2136 avdd.n1027 avdd 12.424
R2137 avdd.n1006 avdd 12.424
R2138 avdd.n1330 avdd 12.424
R2139 avdd.n1526 avdd 12.424
R2140 avdd.n1505 avdd 12.424
R2141 avdd.n1484 avdd 12.424
R2142 avdd.n1463 avdd 12.424
R2143 avdd.n1442 avdd 12.424
R2144 avdd.n1421 avdd 12.424
R2145 avdd.n1400 avdd 12.424
R2146 avdd.n1379 avdd 12.424
R2147 avdd.n1667 avdd 12.424
R2148 avdd.n1687 avdd 12.424
R2149 avdd.n1183 avdd 12.424
R2150 avdd.n1691 avdd 12.2439
R2151 avdd.n974 avdd.n964 11.2946
R2152 avdd.n1710 avdd.n949 11.1593
R2153 avdd.n1775 avdd.n1774 11.0005
R2154 avdd.n1809 avdd.n1808 11.0005
R2155 avdd.n357 avdd.n303 10.9402
R2156 avdd.n355 avdd.n303 10.9402
R2157 avdd.n605 avdd.n551 10.9402
R2158 avdd.n603 avdd.n551 10.9402
R2159 avdd.n1861 avdd.n1860 10.8829
R2160 avdd.n1858 avdd.n1853 10.8829
R2161 avdd.n1875 avdd.n1874 10.8829
R2162 avdd.n1873 avdd.n1872 10.8829
R2163 avdd.n1762 avdd.n1761 10.2783
R2164 avdd.n1764 avdd.n1763 10.2783
R2165 avdd.n1765 avdd.n1764 10.2783
R2166 avdd.n1743 avdd.n1740 10.2783
R2167 avdd.n1744 avdd.n1743 10.2783
R2168 avdd.n1738 avdd.n1735 10.2783
R2169 avdd.n1771 avdd.n1738 10.2783
R2170 avdd.n1774 avdd.n1773 10.2783
R2171 avdd.n1810 avdd.n1809 10.2783
R2172 avdd.n1811 avdd.n1810 10.2783
R2173 avdd.n1193 avdd.n977 10.0697
R2174 avdd.t655 avdd.t441 10.0269
R2175 avdd.t497 avdd.t250 10.0269
R2176 avdd.n479 avdd.n310 9.71534
R2177 avdd.n903 avdd.n558 9.71534
R2178 avdd.n1156 avdd.n1155 9.5406
R2179 avdd.n1135 avdd.n1134 9.5406
R2180 avdd.n1114 avdd.n1113 9.5406
R2181 avdd.n1093 avdd.n1092 9.5406
R2182 avdd.n1072 avdd.n1071 9.5406
R2183 avdd.n1051 avdd.n1050 9.5406
R2184 avdd.n1030 avdd.n1029 9.5406
R2185 avdd.n1009 avdd.n1008 9.5406
R2186 avdd.n1333 avdd.n990 9.5406
R2187 avdd.n1529 avdd.n1528 9.5406
R2188 avdd.n1508 avdd.n1507 9.5406
R2189 avdd.n1487 avdd.n1486 9.5406
R2190 avdd.n1466 avdd.n1465 9.5406
R2191 avdd.n1445 avdd.n1444 9.5406
R2192 avdd.n1424 avdd.n1423 9.5406
R2193 avdd.n1403 avdd.n1402 9.5406
R2194 avdd.n1382 avdd.n1381 9.5406
R2195 avdd.n1670 avdd.n1363 9.5406
R2196 avdd.n1188 avdd.n1187 9.5406
R2197 avdd.n1697 avdd.n959 9.42955
R2198 avdd.n1707 avdd.n1706 9.41227
R2199 avdd.n1855 avdd.n1852 9.3005
R2200 avdd.n1864 avdd.n1836 9.3005
R2201 avdd.n1868 avdd.n17 9.3005
R2202 avdd.n1871 avdd.n1870 9.3005
R2203 avdd.n273 avdd.n20 9.3005
R2204 avdd.n1877 avdd.n1876 9.3005
R2205 avdd.n12 avdd.n11 9.3005
R2206 avdd.n13 avdd.n12 9.3005
R2207 avdd.n3 avdd.n1 9.3005
R2208 avdd.n10 avdd.n9 9.3005
R2209 avdd.n8 avdd.n2 9.3005
R2210 avdd.n985 avdd.n982 9.3005
R2211 avdd.n1333 avdd.n1332 9.3005
R2212 avdd.n1334 avdd.n1333 9.3005
R2213 avdd.n1010 avdd.n1009 9.3005
R2214 avdd.n1009 avdd.n1007 9.3005
R2215 avdd.n1031 avdd.n1030 9.3005
R2216 avdd.n1030 avdd.n1028 9.3005
R2217 avdd.n1052 avdd.n1051 9.3005
R2218 avdd.n1051 avdd.n1049 9.3005
R2219 avdd.n1073 avdd.n1072 9.3005
R2220 avdd.n1072 avdd.n1070 9.3005
R2221 avdd.n1094 avdd.n1093 9.3005
R2222 avdd.n1093 avdd.n1091 9.3005
R2223 avdd.n1115 avdd.n1114 9.3005
R2224 avdd.n1114 avdd.n1112 9.3005
R2225 avdd.n1136 avdd.n1135 9.3005
R2226 avdd.n1135 avdd.n1133 9.3005
R2227 avdd.n1157 avdd.n1156 9.3005
R2228 avdd.n1156 avdd.n1154 9.3005
R2229 avdd.n985 avdd.n984 9.3005
R2230 avdd.n1340 avdd.n1339 9.3005
R2231 avdd.n1339 avdd.n1338 9.3005
R2232 avdd.n1308 avdd.n1307 9.3005
R2233 avdd.n1309 avdd.n1308 9.3005
R2234 avdd.n1293 avdd.n1292 9.3005
R2235 avdd.n1294 avdd.n1293 9.3005
R2236 avdd.n1278 avdd.n1277 9.3005
R2237 avdd.n1279 avdd.n1278 9.3005
R2238 avdd.n1263 avdd.n1262 9.3005
R2239 avdd.n1264 avdd.n1263 9.3005
R2240 avdd.n1248 avdd.n1247 9.3005
R2241 avdd.n1249 avdd.n1248 9.3005
R2242 avdd.n1233 avdd.n1232 9.3005
R2243 avdd.n1234 avdd.n1233 9.3005
R2244 avdd.n1218 avdd.n1217 9.3005
R2245 avdd.n1219 avdd.n1218 9.3005
R2246 avdd.n1203 avdd.n1202 9.3005
R2247 avdd.n1204 avdd.n1203 9.3005
R2248 avdd.n1349 avdd.n1348 9.3005
R2249 avdd.n1347 avdd.n1346 9.3005
R2250 avdd.n1345 avdd.n981 9.3005
R2251 avdd.n1344 avdd.n1343 9.3005
R2252 avdd.n1342 avdd.n1341 9.3005
R2253 avdd.n1335 avdd.n988 9.3005
R2254 avdd.n1318 avdd.n989 9.3005
R2255 avdd.n1331 avdd.n1330 9.3005
R2256 avdd.n1314 avdd.n1313 9.3005
R2257 avdd.n1312 avdd.n1311 9.3005
R2258 avdd.n1310 avdd.n993 9.3005
R2259 avdd.n997 avdd.n996 9.3005
R2260 avdd.n1306 avdd.n1305 9.3005
R2261 avdd.n1304 avdd.n1303 9.3005
R2262 avdd.n1011 avdd.n1006 9.3005
R2263 avdd.n1299 avdd.n1298 9.3005
R2264 avdd.n1297 avdd.n1296 9.3005
R2265 avdd.n1295 avdd.n1014 9.3005
R2266 avdd.n1018 avdd.n1017 9.3005
R2267 avdd.n1291 avdd.n1290 9.3005
R2268 avdd.n1289 avdd.n1288 9.3005
R2269 avdd.n1032 avdd.n1027 9.3005
R2270 avdd.n1284 avdd.n1283 9.3005
R2271 avdd.n1282 avdd.n1281 9.3005
R2272 avdd.n1280 avdd.n1035 9.3005
R2273 avdd.n1039 avdd.n1038 9.3005
R2274 avdd.n1276 avdd.n1275 9.3005
R2275 avdd.n1274 avdd.n1273 9.3005
R2276 avdd.n1053 avdd.n1048 9.3005
R2277 avdd.n1269 avdd.n1268 9.3005
R2278 avdd.n1267 avdd.n1266 9.3005
R2279 avdd.n1265 avdd.n1056 9.3005
R2280 avdd.n1060 avdd.n1059 9.3005
R2281 avdd.n1261 avdd.n1260 9.3005
R2282 avdd.n1259 avdd.n1258 9.3005
R2283 avdd.n1074 avdd.n1069 9.3005
R2284 avdd.n1254 avdd.n1253 9.3005
R2285 avdd.n1252 avdd.n1251 9.3005
R2286 avdd.n1250 avdd.n1077 9.3005
R2287 avdd.n1081 avdd.n1080 9.3005
R2288 avdd.n1246 avdd.n1245 9.3005
R2289 avdd.n1244 avdd.n1243 9.3005
R2290 avdd.n1095 avdd.n1090 9.3005
R2291 avdd.n1239 avdd.n1238 9.3005
R2292 avdd.n1237 avdd.n1236 9.3005
R2293 avdd.n1235 avdd.n1098 9.3005
R2294 avdd.n1102 avdd.n1101 9.3005
R2295 avdd.n1231 avdd.n1230 9.3005
R2296 avdd.n1229 avdd.n1228 9.3005
R2297 avdd.n1116 avdd.n1111 9.3005
R2298 avdd.n1224 avdd.n1223 9.3005
R2299 avdd.n1222 avdd.n1221 9.3005
R2300 avdd.n1220 avdd.n1119 9.3005
R2301 avdd.n1123 avdd.n1122 9.3005
R2302 avdd.n1216 avdd.n1215 9.3005
R2303 avdd.n1214 avdd.n1213 9.3005
R2304 avdd.n1137 avdd.n1132 9.3005
R2305 avdd.n1209 avdd.n1208 9.3005
R2306 avdd.n1207 avdd.n1206 9.3005
R2307 avdd.n1205 avdd.n1140 9.3005
R2308 avdd.n1144 avdd.n1143 9.3005
R2309 avdd.n1201 avdd.n1200 9.3005
R2310 avdd.n1199 avdd.n1198 9.3005
R2311 avdd.n1158 avdd.n1153 9.3005
R2312 avdd.n1358 avdd.n1355 9.3005
R2313 avdd.n1670 avdd.n1669 9.3005
R2314 avdd.n1671 avdd.n1670 9.3005
R2315 avdd.n1383 avdd.n1382 9.3005
R2316 avdd.n1382 avdd.n1380 9.3005
R2317 avdd.n1404 avdd.n1403 9.3005
R2318 avdd.n1403 avdd.n1401 9.3005
R2319 avdd.n1425 avdd.n1424 9.3005
R2320 avdd.n1424 avdd.n1422 9.3005
R2321 avdd.n1446 avdd.n1445 9.3005
R2322 avdd.n1445 avdd.n1443 9.3005
R2323 avdd.n1467 avdd.n1466 9.3005
R2324 avdd.n1466 avdd.n1464 9.3005
R2325 avdd.n1488 avdd.n1487 9.3005
R2326 avdd.n1487 avdd.n1485 9.3005
R2327 avdd.n1509 avdd.n1508 9.3005
R2328 avdd.n1508 avdd.n1506 9.3005
R2329 avdd.n1530 avdd.n1529 9.3005
R2330 avdd.n1529 avdd.n1527 9.3005
R2331 avdd.n1358 avdd.n1357 9.3005
R2332 avdd.n1677 avdd.n1676 9.3005
R2333 avdd.n1676 avdd.n1675 9.3005
R2334 avdd.n1645 avdd.n1644 9.3005
R2335 avdd.n1646 avdd.n1645 9.3005
R2336 avdd.n1630 avdd.n1629 9.3005
R2337 avdd.n1631 avdd.n1630 9.3005
R2338 avdd.n1615 avdd.n1614 9.3005
R2339 avdd.n1616 avdd.n1615 9.3005
R2340 avdd.n1600 avdd.n1599 9.3005
R2341 avdd.n1601 avdd.n1600 9.3005
R2342 avdd.n1585 avdd.n1584 9.3005
R2343 avdd.n1586 avdd.n1585 9.3005
R2344 avdd.n1570 avdd.n1569 9.3005
R2345 avdd.n1571 avdd.n1570 9.3005
R2346 avdd.n1555 avdd.n1554 9.3005
R2347 avdd.n1556 avdd.n1555 9.3005
R2348 avdd.n1540 avdd.n1539 9.3005
R2349 avdd.n1541 avdd.n1540 9.3005
R2350 avdd.n1688 avdd.n1687 9.3005
R2351 avdd.n1686 avdd.n1685 9.3005
R2352 avdd.n1684 avdd.n1683 9.3005
R2353 avdd.n1682 avdd.n1354 9.3005
R2354 avdd.n1681 avdd.n1680 9.3005
R2355 avdd.n1679 avdd.n1678 9.3005
R2356 avdd.n1672 avdd.n1361 9.3005
R2357 avdd.n1655 avdd.n1362 9.3005
R2358 avdd.n1668 avdd.n1667 9.3005
R2359 avdd.n1651 avdd.n1650 9.3005
R2360 avdd.n1649 avdd.n1648 9.3005
R2361 avdd.n1647 avdd.n1366 9.3005
R2362 avdd.n1370 avdd.n1369 9.3005
R2363 avdd.n1643 avdd.n1642 9.3005
R2364 avdd.n1641 avdd.n1640 9.3005
R2365 avdd.n1384 avdd.n1379 9.3005
R2366 avdd.n1636 avdd.n1635 9.3005
R2367 avdd.n1634 avdd.n1633 9.3005
R2368 avdd.n1632 avdd.n1387 9.3005
R2369 avdd.n1391 avdd.n1390 9.3005
R2370 avdd.n1628 avdd.n1627 9.3005
R2371 avdd.n1626 avdd.n1625 9.3005
R2372 avdd.n1405 avdd.n1400 9.3005
R2373 avdd.n1621 avdd.n1620 9.3005
R2374 avdd.n1619 avdd.n1618 9.3005
R2375 avdd.n1617 avdd.n1408 9.3005
R2376 avdd.n1412 avdd.n1411 9.3005
R2377 avdd.n1613 avdd.n1612 9.3005
R2378 avdd.n1611 avdd.n1610 9.3005
R2379 avdd.n1426 avdd.n1421 9.3005
R2380 avdd.n1606 avdd.n1605 9.3005
R2381 avdd.n1604 avdd.n1603 9.3005
R2382 avdd.n1602 avdd.n1429 9.3005
R2383 avdd.n1433 avdd.n1432 9.3005
R2384 avdd.n1598 avdd.n1597 9.3005
R2385 avdd.n1596 avdd.n1595 9.3005
R2386 avdd.n1447 avdd.n1442 9.3005
R2387 avdd.n1591 avdd.n1590 9.3005
R2388 avdd.n1589 avdd.n1588 9.3005
R2389 avdd.n1587 avdd.n1450 9.3005
R2390 avdd.n1454 avdd.n1453 9.3005
R2391 avdd.n1583 avdd.n1582 9.3005
R2392 avdd.n1581 avdd.n1580 9.3005
R2393 avdd.n1468 avdd.n1463 9.3005
R2394 avdd.n1576 avdd.n1575 9.3005
R2395 avdd.n1574 avdd.n1573 9.3005
R2396 avdd.n1572 avdd.n1471 9.3005
R2397 avdd.n1475 avdd.n1474 9.3005
R2398 avdd.n1568 avdd.n1567 9.3005
R2399 avdd.n1566 avdd.n1565 9.3005
R2400 avdd.n1489 avdd.n1484 9.3005
R2401 avdd.n1561 avdd.n1560 9.3005
R2402 avdd.n1559 avdd.n1558 9.3005
R2403 avdd.n1557 avdd.n1492 9.3005
R2404 avdd.n1496 avdd.n1495 9.3005
R2405 avdd.n1553 avdd.n1552 9.3005
R2406 avdd.n1551 avdd.n1550 9.3005
R2407 avdd.n1510 avdd.n1505 9.3005
R2408 avdd.n1546 avdd.n1545 9.3005
R2409 avdd.n1544 avdd.n1543 9.3005
R2410 avdd.n1542 avdd.n1513 9.3005
R2411 avdd.n1517 avdd.n1516 9.3005
R2412 avdd.n1538 avdd.n1537 9.3005
R2413 avdd.n1536 avdd.n1535 9.3005
R2414 avdd.n1531 avdd.n1526 9.3005
R2415 avdd.n1189 avdd.n1188 9.3005
R2416 avdd.n1188 avdd.n1186 9.3005
R2417 avdd.n1175 avdd.n1174 9.3005
R2418 avdd.n1176 avdd.n1175 9.3005
R2419 avdd.n1179 avdd.n1178 9.3005
R2420 avdd.n1177 avdd.n1165 9.3005
R2421 avdd.n1172 avdd.n1171 9.3005
R2422 avdd.n1173 avdd.n1160 9.3005
R2423 avdd.n1185 avdd.n1184 9.3005
R2424 avdd.n1183 avdd.n1159 9.3005
R2425 avdd.n1829 avdd.n1828 9.3005
R2426 avdd.n1808 avdd.n1807 9.3005
R2427 avdd.n1776 avdd.n1775 9.3005
R2428 avdd.n788 avdd.n787 9.3005
R2429 avdd.n784 avdd.n783 9.3005
R2430 avdd.n782 avdd.n781 9.3005
R2431 avdd.n780 avdd.n620 9.3005
R2432 avdd.n779 avdd.n778 9.3005
R2433 avdd.n669 avdd.n664 9.3005
R2434 avdd.n671 avdd.n670 9.3005
R2435 avdd.n660 avdd.n659 9.3005
R2436 avdd.n679 avdd.n678 9.3005
R2437 avdd.n680 avdd.n658 9.3005
R2438 avdd.n682 avdd.n681 9.3005
R2439 avdd.n655 avdd.n654 9.3005
R2440 avdd.n689 avdd.n688 9.3005
R2441 avdd.n690 avdd.n653 9.3005
R2442 avdd.n692 avdd.n691 9.3005
R2443 avdd.n649 avdd.n648 9.3005
R2444 avdd.n700 avdd.n699 9.3005
R2445 avdd.n701 avdd.n647 9.3005
R2446 avdd.n703 avdd.n702 9.3005
R2447 avdd.n644 avdd.n643 9.3005
R2448 avdd.n710 avdd.n709 9.3005
R2449 avdd.n711 avdd.n642 9.3005
R2450 avdd.n713 avdd.n712 9.3005
R2451 avdd.n638 avdd.n637 9.3005
R2452 avdd.n721 avdd.n720 9.3005
R2453 avdd.n722 avdd.n636 9.3005
R2454 avdd.n724 avdd.n723 9.3005
R2455 avdd.n633 avdd.n632 9.3005
R2456 avdd.n732 avdd.n731 9.3005
R2457 avdd.n733 avdd.n631 9.3005
R2458 avdd.n735 avdd.n734 9.3005
R2459 avdd.n628 avdd.n627 9.3005
R2460 avdd.n743 avdd.n742 9.3005
R2461 avdd.n744 avdd.n625 9.3005
R2462 avdd.n767 avdd.n766 9.3005
R2463 avdd.n765 avdd.n626 9.3005
R2464 avdd.n764 avdd.n623 9.3005
R2465 avdd.n789 avdd.n788 9.3005
R2466 avdd.n617 avdd.n616 9.3005
R2467 avdd.n251 avdd.n26 9.3005
R2468 avdd.n252 avdd.n251 9.3005
R2469 avdd.n240 avdd.n33 9.3005
R2470 avdd.n241 avdd.n240 9.3005
R2471 avdd.n41 avdd.n40 9.3005
R2472 avdd.n42 avdd.n41 9.3005
R2473 avdd.n228 avdd.n227 9.3005
R2474 avdd.n227 avdd.n226 9.3005
R2475 avdd.n215 avdd.n53 9.3005
R2476 avdd.n216 avdd.n215 9.3005
R2477 avdd.n61 avdd.n60 9.3005
R2478 avdd.n62 avdd.n61 9.3005
R2479 avdd.n203 avdd.n202 9.3005
R2480 avdd.n202 avdd.n201 9.3005
R2481 avdd.n190 avdd.n73 9.3005
R2482 avdd.n191 avdd.n190 9.3005
R2483 avdd.n81 avdd.n80 9.3005
R2484 avdd.n82 avdd.n81 9.3005
R2485 avdd.n178 avdd.n177 9.3005
R2486 avdd.n177 avdd.n176 9.3005
R2487 avdd.n165 avdd.n93 9.3005
R2488 avdd.n166 avdd.n165 9.3005
R2489 avdd.n101 avdd.n100 9.3005
R2490 avdd.n102 avdd.n101 9.3005
R2491 avdd.n153 avdd.n152 9.3005
R2492 avdd.n152 avdd.n151 9.3005
R2493 avdd.n140 avdd.n113 9.3005
R2494 avdd.n141 avdd.n140 9.3005
R2495 avdd.n121 avdd.n120 9.3005
R2496 avdd.n122 avdd.n121 9.3005
R2497 avdd.n128 avdd.n127 9.3005
R2498 avdd.n127 avdd.n0 9.3005
R2499 avdd.n257 avdd.n256 9.3005
R2500 avdd.n255 avdd.n22 9.3005
R2501 avdd.n254 avdd.n253 9.3005
R2502 avdd.n250 avdd.n249 9.3005
R2503 avdd.n28 avdd.n27 9.3005
R2504 avdd.n243 avdd.n242 9.3005
R2505 avdd.n239 avdd.n238 9.3005
R2506 avdd.n35 avdd.n34 9.3005
R2507 avdd.n39 avdd.n38 9.3005
R2508 avdd.n231 avdd.n43 9.3005
R2509 avdd.n230 avdd.n229 9.3005
R2510 avdd.n45 avdd.n44 9.3005
R2511 avdd.n225 avdd.n224 9.3005
R2512 avdd.n47 avdd.n46 9.3005
R2513 avdd.n218 avdd.n217 9.3005
R2514 avdd.n214 avdd.n213 9.3005
R2515 avdd.n55 avdd.n54 9.3005
R2516 avdd.n59 avdd.n58 9.3005
R2517 avdd.n206 avdd.n63 9.3005
R2518 avdd.n205 avdd.n204 9.3005
R2519 avdd.n65 avdd.n64 9.3005
R2520 avdd.n200 avdd.n199 9.3005
R2521 avdd.n67 avdd.n66 9.3005
R2522 avdd.n193 avdd.n192 9.3005
R2523 avdd.n189 avdd.n188 9.3005
R2524 avdd.n75 avdd.n74 9.3005
R2525 avdd.n79 avdd.n78 9.3005
R2526 avdd.n181 avdd.n83 9.3005
R2527 avdd.n180 avdd.n179 9.3005
R2528 avdd.n85 avdd.n84 9.3005
R2529 avdd.n175 avdd.n174 9.3005
R2530 avdd.n87 avdd.n86 9.3005
R2531 avdd.n168 avdd.n167 9.3005
R2532 avdd.n164 avdd.n163 9.3005
R2533 avdd.n95 avdd.n94 9.3005
R2534 avdd.n99 avdd.n98 9.3005
R2535 avdd.n156 avdd.n103 9.3005
R2536 avdd.n155 avdd.n154 9.3005
R2537 avdd.n105 avdd.n104 9.3005
R2538 avdd.n150 avdd.n149 9.3005
R2539 avdd.n107 avdd.n106 9.3005
R2540 avdd.n143 avdd.n142 9.3005
R2541 avdd.n139 avdd.n138 9.3005
R2542 avdd.n115 avdd.n114 9.3005
R2543 avdd.n119 avdd.n118 9.3005
R2544 avdd.n131 avdd.n123 9.3005
R2545 avdd.n130 avdd.n129 9.3005
R2546 avdd.n126 avdd.n125 9.3005
R2547 avdd.n1870 avdd.n1869 9.2699
R2548 avdd.n1869 avdd.n1868 9.2699
R2549 avdd.n1698 avdd.n975 8.94982
R2550 avdd.n293 avdd.n291 8.40959
R2551 avdd.n293 avdd.n287 8.40959
R2552 avdd.n297 avdd.n292 8.40959
R2553 avdd.n297 avdd.n287 8.40959
R2554 avdd.n451 avdd.n450 8.40959
R2555 avdd.n452 avdd.n451 8.40959
R2556 avdd.n491 avdd.n490 8.40959
R2557 avdd.n492 avdd.n491 8.40959
R2558 avdd.n541 avdd.n539 8.40959
R2559 avdd.n541 avdd.n535 8.40959
R2560 avdd.n545 avdd.n540 8.40959
R2561 avdd.n545 avdd.n535 8.40959
R2562 avdd.n875 avdd.n874 8.40959
R2563 avdd.n876 avdd.n875 8.40959
R2564 avdd.n915 avdd.n914 8.40959
R2565 avdd.n916 avdd.n915 8.40959
R2566 avdd.n464 avdd.n347 8.24855
R2567 avdd.n888 avdd.n595 8.24855
R2568 avdd.n523 avdd.n522 8.24253
R2569 avdd.n947 avdd.n946 8.24253
R2570 avdd.n474 avdd.n337 8.18605
R2571 avdd.n898 avdd.n585 8.18605
R2572 avdd.n475 avdd.n474 8.17238
R2573 avdd.n899 avdd.n898 8.17238
R2574 avdd.n464 avdd.n463 8.10988
R2575 avdd.n888 avdd.n887 8.10988
R2576 avdd.n1833 avdd.n1832 7.90948
R2577 avdd.n434 avdd.n433 7.90079
R2578 avdd.n858 avdd.n857 7.68198
R2579 avdd.n1728 avdd.n1727 7.56644
R2580 avdd.n1829 avdd.n1733 7.55653
R2581 avdd.n1746 avdd.n1733 7.55653
R2582 avdd.n1825 avdd.n1824 7.4005
R2583 avdd.t120 avdd.n1825 7.4005
R2584 avdd.n1827 avdd.n1826 7.4005
R2585 avdd.n1826 avdd.t120 7.4005
R2586 avdd.n676 avdd.t322 7.30819
R2587 avdd.t326 avdd.n640 7.30819
R2588 avdd.n348 avdd.n337 7.29542
R2589 avdd.n596 avdd.n585 7.29542
R2590 avdd.n1746 avdd.n1734 7.06516
R2591 avdd.n1829 avdd.n1734 7.06516
R2592 avdd.n1155 avdd 7.01471
R2593 avdd.n1134 avdd 7.01471
R2594 avdd.n1113 avdd 7.01471
R2595 avdd.n1092 avdd 7.01471
R2596 avdd.n1071 avdd 7.01471
R2597 avdd.n1050 avdd 7.01471
R2598 avdd.n1029 avdd 7.01471
R2599 avdd.n1008 avdd 7.01471
R2600 avdd.n990 avdd 7.01471
R2601 avdd.n1528 avdd 7.01471
R2602 avdd.n1507 avdd 7.01471
R2603 avdd.n1486 avdd 7.01471
R2604 avdd.n1465 avdd 7.01471
R2605 avdd.n1444 avdd 7.01471
R2606 avdd.n1423 avdd 7.01471
R2607 avdd.n1402 avdd 7.01471
R2608 avdd.n1381 avdd 7.01471
R2609 avdd.n1363 avdd 7.01471
R2610 avdd.n1187 avdd 7.01471
R2611 avdd.n463 avdd.n349 6.77003
R2612 avdd.n347 avdd.n346 6.77003
R2613 avdd.n887 avdd.n597 6.77003
R2614 avdd.n595 avdd.n594 6.77003
R2615 avdd.n366 avdd.n361 6.60764
R2616 avdd.n448 avdd.n361 6.60764
R2617 avdd.n447 avdd.n446 6.60764
R2618 avdd.n448 avdd.n447 6.60764
R2619 avdd.n614 avdd.n609 6.60764
R2620 avdd.n872 avdd.n609 6.60764
R2621 avdd.n871 avdd.n870 6.60764
R2622 avdd.n872 avdd.n871 6.60764
R2623 avdd.n475 avdd.n338 6.59816
R2624 avdd.n899 avdd.n586 6.59816
R2625 avdd.n479 avdd.n478 6.47706
R2626 avdd.n903 avdd.n902 6.47706
R2627 avdd.n668 avdd.n665 6.11192
R2628 avdd.n1833 avdd.n276 5.9555
R2629 avdd.n1166 avdd 5.7342
R2630 avdd.n1866 avdd.n1865 5.7183
R2631 avdd.n1781 avdd.n1780 5.70732
R2632 avdd.n1806 avdd.n1805 5.70732
R2633 avdd.n1788 avdd.n1787 5.70732
R2634 avdd.n1781 avdd.n1776 5.70369
R2635 avdd.n1852 avdd.n1851 5.70305
R2636 avdd.n1807 avdd.n1806 5.70274
R2637 avdd.n1747 avdd.n1746 5.70242
R2638 avdd.n1865 avdd.n1864 5.6605
R2639 avdd.n1830 avdd.n1829 5.6605
R2640 avdd.n1793 avdd.n1792 5.6605
R2641 avdd.n1849 avdd.t233 5.5395
R2642 avdd.n1849 avdd.t221 5.5395
R2643 avdd.n1847 avdd.t243 5.5395
R2644 avdd.n1847 avdd.t235 5.5395
R2645 avdd.n1845 avdd.t239 5.5395
R2646 avdd.n1845 avdd.t237 5.5395
R2647 avdd.n1843 avdd.t227 5.5395
R2648 avdd.n1843 avdd.t225 5.5395
R2649 avdd.n1841 avdd.t229 5.5395
R2650 avdd.n1841 avdd.t231 5.5395
R2651 avdd.n1839 avdd.t245 5.5395
R2652 avdd.n1839 avdd.t241 5.5395
R2653 avdd.n1837 avdd.t223 5.5395
R2654 avdd.n1837 avdd.t249 5.5395
R2655 avdd.n1789 avdd.t381 5.5395
R2656 avdd.t25 avdd.n1789 5.5395
R2657 avdd.n1731 avdd.t177 5.5395
R2658 avdd.n1731 avdd.t582 5.5395
R2659 avdd.n1755 avdd.t614 5.5395
R2660 avdd.n1755 avdd.t604 5.5395
R2661 avdd.n1757 avdd.t612 5.5395
R2662 avdd.n1757 avdd.t578 5.5395
R2663 avdd.n1786 avdd.t549 5.5395
R2664 avdd.n1786 avdd.t116 5.5395
R2665 avdd.n1782 avdd.t555 5.5395
R2666 avdd.n1782 avdd.t45 5.5395
R2667 avdd.t116 avdd.n1785 5.5395
R2668 avdd.n1785 avdd.t553 5.5395
R2669 avdd.n1790 avdd.t25 5.5395
R2670 avdd.n1790 avdd.t551 5.5395
R2671 avdd.n1797 avdd.t385 5.5395
R2672 avdd.n1797 avdd.t379 5.5395
R2673 avdd.n1799 avdd.t622 5.5395
R2674 avdd.n1799 avdd.t387 5.5395
R2675 avdd.n1801 avdd.t389 5.5395
R2676 avdd.n1801 avdd.t624 5.5395
R2677 avdd.t162 avdd.n1804 5.5395
R2678 avdd.n1804 avdd.t383 5.5395
R2679 avdd.n1863 avdd.n1852 5.48326
R2680 avdd.n1864 avdd.n1863 5.48326
R2681 avdd.n30 avdd.t619 5.48127
R2682 avdd.t390 avdd.n246 5.48127
R2683 avdd.n235 avdd.t503 5.48127
R2684 avdd.n49 avdd.t572 5.48127
R2685 avdd.t178 avdd.n221 5.48127
R2686 avdd.n210 avdd.t473 5.48127
R2687 avdd.n69 avdd.t518 5.48127
R2688 avdd.t423 avdd.n196 5.48127
R2689 avdd.n185 avdd.t435 5.48127
R2690 avdd.n89 avdd.t592 5.48127
R2691 avdd.t466 avdd.n171 5.48127
R2692 avdd.n160 avdd.t600 5.48127
R2693 avdd.n109 avdd.t449 5.48127
R2694 avdd.t0 avdd.n146 5.48127
R2695 avdd.n135 avdd.t258 5.48127
R2696 avdd.n1693 avdd.n525 5.3849
R2697 avdd.n1821 avdd.n1820 5.28621
R2698 avdd.n1820 avdd.t613 5.28621
R2699 avdd.n1819 avdd.n1818 5.28621
R2700 avdd.t613 avdd.n1819 5.28621
R2701 avdd.n311 avdd.n280 5.22511
R2702 avdd.n458 avdd.n310 5.22511
R2703 avdd.n559 avdd.n528 5.22511
R2704 avdd.n882 avdd.n558 5.22511
R2705 avdd.n462 avdd.n461 5.11573
R2706 avdd.n886 avdd.n885 5.11573
R2707 avdd.n358 avdd.n310 4.98102
R2708 avdd.n606 avdd.n558 4.98102
R2709 avdd.n354 avdd.n311 4.94972
R2710 avdd.n602 avdd.n559 4.94972
R2711 avdd.n973 avdd.n970 4.89462
R2712 avdd.n969 avdd.n967 4.89462
R2713 avdd.n449 avdd.n360 4.86892
R2714 avdd.n452 avdd.n449 4.86892
R2715 avdd.n352 avdd.n286 4.86892
R2716 avdd.n492 avdd.n286 4.86892
R2717 avdd.n873 avdd.n608 4.86892
R2718 avdd.n876 avdd.n873 4.86892
R2719 avdd.n600 avdd.n534 4.86892
R2720 avdd.n916 avdd.n534 4.86892
R2721 avdd.n1693 avdd.n524 4.85844
R2722 avdd.n857 avdd.n790 4.76569
R2723 avdd.n280 avdd.n279 4.66083
R2724 avdd.n459 avdd.n458 4.66083
R2725 avdd.n528 avdd.n527 4.66083
R2726 avdd.n883 avdd.n882 4.66083
R2727 avdd.n1694 avdd.n1692 4.55185
R2728 avdd.n499 avdd.n498 4.5005
R2729 avdd.n501 avdd.n500 4.5005
R2730 avdd.n503 avdd.n502 4.5005
R2731 avdd.n505 avdd.n504 4.5005
R2732 avdd.n507 avdd.n506 4.5005
R2733 avdd.n509 avdd.n508 4.5005
R2734 avdd.n511 avdd.n510 4.5005
R2735 avdd.n513 avdd.n512 4.5005
R2736 avdd.n515 avdd.n514 4.5005
R2737 avdd.n517 avdd.n516 4.5005
R2738 avdd.n519 avdd.n518 4.5005
R2739 avdd.n476 avdd.n475 4.5005
R2740 avdd.n346 avdd.n309 4.5005
R2741 avdd.n462 avdd.n347 4.5005
R2742 avdd.n395 avdd.n351 4.5005
R2743 avdd.n398 avdd.n394 4.5005
R2744 avdd.n404 avdd.n403 4.5005
R2745 avdd.n407 avdd.n406 4.5005
R2746 avdd.n409 avdd.n408 4.5005
R2747 avdd.n412 avdd.n392 4.5005
R2748 avdd.n418 avdd.n417 4.5005
R2749 avdd.n421 avdd.n420 4.5005
R2750 avdd.n423 avdd.n422 4.5005
R2751 avdd.n426 avdd.n390 4.5005
R2752 avdd.n432 avdd.n431 4.5005
R2753 avdd.n480 avdd.n479 4.5005
R2754 avdd.n478 avdd.n477 4.5005
R2755 avdd.n923 avdd.n922 4.5005
R2756 avdd.n925 avdd.n924 4.5005
R2757 avdd.n927 avdd.n926 4.5005
R2758 avdd.n929 avdd.n928 4.5005
R2759 avdd.n931 avdd.n930 4.5005
R2760 avdd.n933 avdd.n932 4.5005
R2761 avdd.n935 avdd.n934 4.5005
R2762 avdd.n937 avdd.n936 4.5005
R2763 avdd.n939 avdd.n938 4.5005
R2764 avdd.n941 avdd.n940 4.5005
R2765 avdd.n943 avdd.n942 4.5005
R2766 avdd.n900 avdd.n899 4.5005
R2767 avdd.n594 avdd.n557 4.5005
R2768 avdd.n886 avdd.n595 4.5005
R2769 avdd.n818 avdd.n599 4.5005
R2770 avdd.n821 avdd.n817 4.5005
R2771 avdd.n827 avdd.n826 4.5005
R2772 avdd.n830 avdd.n829 4.5005
R2773 avdd.n832 avdd.n831 4.5005
R2774 avdd.n835 avdd.n815 4.5005
R2775 avdd.n841 avdd.n840 4.5005
R2776 avdd.n844 avdd.n843 4.5005
R2777 avdd.n846 avdd.n845 4.5005
R2778 avdd.n849 avdd.n813 4.5005
R2779 avdd.n855 avdd.n854 4.5005
R2780 avdd.n904 avdd.n903 4.5005
R2781 avdd.n902 avdd.n901 4.5005
R2782 avdd.n1832 avdd.n1729 4.4965
R2783 avdd.n984 avdd 4.46111
R2784 avdd.n984 avdd 4.46111
R2785 avdd.n1357 avdd 4.46111
R2786 avdd.n1357 avdd 4.46111
R2787 avdd.n520 avdd.n519 4.45347
R2788 avdd.n388 avdd.n387 4.45347
R2789 avdd.n429 avdd.n389 4.45347
R2790 avdd.n313 avdd.n278 4.45347
R2791 avdd.n433 avdd.n432 4.45347
R2792 avdd.n944 avdd.n943 4.45347
R2793 avdd.n811 avdd.n810 4.45347
R2794 avdd.n852 avdd.n812 4.45347
R2795 avdd.n561 avdd.n526 4.45347
R2796 avdd.n856 avdd.n855 4.45347
R2797 avdd.n477 avdd.n476 4.39112
R2798 avdd.n901 avdd.n900 4.39112
R2799 avdd.n1692 avdd.n276 4.28658
R2800 avdd.n1862 avdd.n1854 4.20505
R2801 avdd.n1859 avdd.n1854 4.20505
R2802 avdd.n1857 avdd.n1856 4.20505
R2803 avdd.n1859 avdd.n1857 4.20505
R2804 avdd.n480 avdd.n309 4.16066
R2805 avdd.n904 avdd.n557 4.16066
R2806 avdd.n1832 avdd.n1831 4.15861
R2807 avdd.n1716 avdd.n1715 4.14168
R2808 avdd.n1351 avdd.n977 4.12179
R2809 avdd.n1831 avdd.n1830 4.01324
R2810 avdd.n1864 avdd.n1835 3.91429
R2811 avdd.n1852 avdd.n1835 3.91429
R2812 avdd.n1142 avdd 3.7406
R2813 avdd.n1121 avdd 3.7406
R2814 avdd.n1100 avdd 3.7406
R2815 avdd.n1079 avdd 3.7406
R2816 avdd.n1058 avdd 3.7406
R2817 avdd.n1037 avdd 3.7406
R2818 avdd.n1016 avdd 3.7406
R2819 avdd.n995 avdd 3.7406
R2820 avdd.n1337 avdd 3.7406
R2821 avdd.n1515 avdd 3.7406
R2822 avdd.n1494 avdd 3.7406
R2823 avdd.n1473 avdd 3.7406
R2824 avdd.n1452 avdd 3.7406
R2825 avdd.n1431 avdd 3.7406
R2826 avdd.n1410 avdd 3.7406
R2827 avdd.n1389 avdd 3.7406
R2828 avdd.n1368 avdd 3.7406
R2829 avdd.n1674 avdd 3.7406
R2830 avdd.n1168 avdd 3.7406
R2831 avdd.n1166 avdd 3.56469
R2832 avdd.n1166 avdd 3.56469
R2833 avdd.n964 avdd.n963 3.55819
R2834 avdd.n963 avdd.n962 3.55819
R2835 avdd.n1696 avdd.n1695 3.40737
R2836 avdd.n478 avdd.n311 3.23878
R2837 avdd.n902 avdd.n559 3.23878
R2838 avdd.n1717 avdd.n1716 2.93701
R2839 avdd.n1718 avdd.n1717 2.93701
R2840 avdd.n467 avdd.n466 2.80353
R2841 avdd.n468 avdd.n467 2.80353
R2842 avdd.n472 avdd.n471 2.80353
R2843 avdd.n471 avdd.n470 2.80353
R2844 avdd.n891 avdd.n890 2.80353
R2845 avdd.n892 avdd.n891 2.80353
R2846 avdd.n896 avdd.n895 2.80353
R2847 avdd.n895 avdd.n894 2.80353
R2848 avdd.n977 avdd.n525 2.68185
R2849 avdd.n1701 avdd.n1700 2.28445
R2850 avdd.n1702 avdd.n1701 2.28445
R2851 avdd.n1726 avdd.n1725 2.27397
R2852 avdd.n1694 avdd 2.19329
R2853 avdd.n1193 avdd 2.07277
R2854 avdd.n1831 avdd.n1730 1.97988
R2855 avdd.n1777 avdd.n1770 1.97248
R2856 avdd.n1796 avdd.n1795 1.97248
R2857 avdd.n669 avdd.n668 1.87847
R2858 avdd.t386 avdd.n1771 1.86325
R2859 avdd.n1727 avdd.n1726 1.7055
R2860 avdd.n1194 avdd.n976 1.69386
R2861 avdd.n355 avdd.n354 1.61378
R2862 avdd.n603 avdd.n602 1.61378
R2863 avdd.n358 avdd.n357 1.55875
R2864 avdd.n606 avdd.n605 1.55875
R2865 avdd.n950 avdd.n948 1.5505
R2866 avdd.n1779 avdd.n1778 1.52433
R2867 avdd.n473 avdd.n472 1.50638
R2868 avdd.n897 avdd.n896 1.50638
R2869 avdd.n18 avdd.n16 1.4805
R2870 avdd.t38 avdd.n18 1.4805
R2871 avdd.n21 avdd.n19 1.4805
R2872 avdd.t38 avdd.n19 1.4805
R2873 avdd.n1695 avdd.n976 1.37843
R2874 avdd.n1794 avdd.n1793 1.31832
R2875 avdd.n273 avdd.n272 1.28283
R2876 avdd.n290 avdd.n288 1.2505
R2877 avdd.n486 avdd.n288 1.2505
R2878 avdd.n488 avdd.n487 1.2505
R2879 avdd.n487 avdd.n486 1.2505
R2880 avdd.n485 avdd.n484 1.2505
R2881 avdd.n486 avdd.n485 1.2505
R2882 avdd.n285 avdd.n283 1.2505
R2883 avdd.n486 avdd.n285 1.2505
R2884 avdd.n538 avdd.n536 1.2505
R2885 avdd.n910 avdd.n536 1.2505
R2886 avdd.n912 avdd.n911 1.2505
R2887 avdd.n911 avdd.n910 1.2505
R2888 avdd.n909 avdd.n908 1.2505
R2889 avdd.n910 avdd.n909 1.2505
R2890 avdd.n533 avdd.n531 1.2505
R2891 avdd.n910 avdd.n533 1.2505
R2892 avdd.n1351 avdd.n1350 1.20459
R2893 avdd.n1690 avdd.n1689 1.1873
R2894 avdd.n274 avdd.n257 1.16964
R2895 avdd.n272 avdd.n271 1.15136
R2896 avdd.n271 avdd.n270 1.15136
R2897 avdd.n270 avdd.n269 1.15136
R2898 avdd.n269 avdd.n268 1.15136
R2899 avdd.n268 avdd.n267 1.15136
R2900 avdd.n267 avdd.n266 1.15136
R2901 avdd.n264 avdd.n263 1.15136
R2902 avdd.n263 avdd.n262 1.15136
R2903 avdd.n262 avdd.n261 1.15136
R2904 avdd.n261 avdd.n260 1.15136
R2905 avdd.n260 avdd.n259 1.15136
R2906 avdd.n259 avdd.n258 1.15136
R2907 avdd.n258 avdd.n15 1.15136
R2908 avdd.n344 avdd.n341 1.14248
R2909 avdd.n343 avdd.n341 1.14248
R2910 avdd.n342 avdd.n340 1.14248
R2911 avdd.n469 avdd.n342 1.14248
R2912 avdd.n592 avdd.n589 1.14248
R2913 avdd.n591 avdd.n589 1.14248
R2914 avdd.n590 avdd.n588 1.14248
R2915 avdd.n893 avdd.n590 1.14248
R2916 avdd.n524 avdd 1.13913
R2917 avdd.n1877 avdd.n15 1.13628
R2918 avdd.n1712 avdd.n958 1.12991
R2919 avdd.n266 avdd.n265 1.0824
R2920 avdd.n389 avdd.n388 1.05355
R2921 avdd.n388 avdd.n278 1.05355
R2922 avdd.n812 avdd.n811 1.05355
R2923 avdd.n811 avdd.n526 1.05355
R2924 avdd.n513 avdd.n511 1.04347
R2925 avdd.n381 avdd.n379 1.04347
R2926 avdd.n321 avdd.n319 1.04347
R2927 avdd.n415 avdd.n391 1.04347
R2928 avdd.n421 avdd.n418 1.04347
R2929 avdd.n937 avdd.n935 1.04347
R2930 avdd.n804 avdd.n802 1.04347
R2931 avdd.n569 avdd.n567 1.04347
R2932 avdd.n838 avdd.n814 1.04347
R2933 avdd.n844 avdd.n841 1.04347
R2934 avdd.n951 avdd.n277 1.03383
R2935 avdd.n958 avdd.n953 0.989805
R2936 avdd.n1719 avdd.n953 0.989805
R2937 avdd.n276 avdd.n275 0.986125
R2938 avdd avdd.n1194 0.983
R2939 avdd avdd.n976 0.983
R2940 avdd.n973 avdd.n972 0.954108
R2941 avdd.n972 avdd.n971 0.954108
R2942 avdd.n1768 avdd.n1766 0.907363
R2943 avdd.n1772 avdd.n1766 0.907363
R2944 avdd.n1769 avdd.n1767 0.907363
R2945 avdd.n1772 avdd.n1767 0.907363
R2946 avdd.n1866 avdd.n1833 0.90425
R2947 avdd.n1706 avdd.n1705 0.877277
R2948 avdd.n1705 avdd.n1704 0.877277
R2949 avdd.n1697 avdd 0.876125
R2950 avdd.n275 avdd.n274 0.83425
R2951 avdd.n346 avdd.n338 0.773938
R2952 avdd.n594 avdd.n586 0.773938
R2953 avdd avdd.n1314 0.755
R2954 avdd avdd.n1299 0.755
R2955 avdd avdd.n1284 0.755
R2956 avdd avdd.n1269 0.755
R2957 avdd avdd.n1254 0.755
R2958 avdd avdd.n1239 0.755
R2959 avdd avdd.n1224 0.755
R2960 avdd avdd.n1209 0.755
R2961 avdd avdd.n1651 0.755
R2962 avdd avdd.n1636 0.755
R2963 avdd avdd.n1621 0.755
R2964 avdd avdd.n1606 0.755
R2965 avdd avdd.n1591 0.755
R2966 avdd avdd.n1576 0.755
R2967 avdd avdd.n1561 0.755
R2968 avdd avdd.n1546 0.755
R2969 avdd.n477 avdd.n336 0.725109
R2970 avdd.n901 avdd.n584 0.725109
R2971 avdd.n522 avdd.n521 0.713391
R2972 avdd.n519 avdd.n517 0.713391
R2973 avdd.n517 avdd.n515 0.713391
R2974 avdd.n515 avdd.n513 0.713391
R2975 avdd.n511 avdd.n509 0.713391
R2976 avdd.n509 avdd.n507 0.713391
R2977 avdd.n507 avdd.n505 0.713391
R2978 avdd.n505 avdd.n503 0.713391
R2979 avdd.n503 avdd.n501 0.713391
R2980 avdd.n501 avdd.n499 0.713391
R2981 avdd.n387 avdd.n385 0.713391
R2982 avdd.n385 avdd.n383 0.713391
R2983 avdd.n383 avdd.n381 0.713391
R2984 avdd.n379 avdd.n377 0.713391
R2985 avdd.n377 avdd.n375 0.713391
R2986 avdd.n375 avdd.n373 0.713391
R2987 avdd.n373 avdd.n371 0.713391
R2988 avdd.n371 avdd.n369 0.713391
R2989 avdd.n369 avdd.n308 0.713391
R2990 avdd.n315 avdd.n313 0.713391
R2991 avdd.n317 avdd.n315 0.713391
R2992 avdd.n319 avdd.n317 0.713391
R2993 avdd.n323 avdd.n321 0.713391
R2994 avdd.n325 avdd.n323 0.713391
R2995 avdd.n327 avdd.n325 0.713391
R2996 avdd.n329 avdd.n327 0.713391
R2997 avdd.n331 avdd.n329 0.713391
R2998 avdd.n333 avdd.n331 0.713391
R2999 avdd.n429 avdd.n428 0.713391
R3000 avdd.n428 avdd.n425 0.713391
R3001 avdd.n425 avdd.n391 0.713391
R3002 avdd.n415 avdd.n414 0.713391
R3003 avdd.n414 avdd.n411 0.713391
R3004 avdd.n411 avdd.n393 0.713391
R3005 avdd.n401 avdd.n393 0.713391
R3006 avdd.n401 avdd.n400 0.713391
R3007 avdd.n400 avdd.n397 0.713391
R3008 avdd.n432 avdd.n390 0.713391
R3009 avdd.n422 avdd.n390 0.713391
R3010 avdd.n422 avdd.n421 0.713391
R3011 avdd.n418 avdd.n392 0.713391
R3012 avdd.n408 avdd.n392 0.713391
R3013 avdd.n408 avdd.n407 0.713391
R3014 avdd.n407 avdd.n404 0.713391
R3015 avdd.n404 avdd.n394 0.713391
R3016 avdd.n394 avdd.n351 0.713391
R3017 avdd.n946 avdd.n945 0.713391
R3018 avdd.n943 avdd.n941 0.713391
R3019 avdd.n941 avdd.n939 0.713391
R3020 avdd.n939 avdd.n937 0.713391
R3021 avdd.n935 avdd.n933 0.713391
R3022 avdd.n933 avdd.n931 0.713391
R3023 avdd.n931 avdd.n929 0.713391
R3024 avdd.n929 avdd.n927 0.713391
R3025 avdd.n927 avdd.n925 0.713391
R3026 avdd.n925 avdd.n923 0.713391
R3027 avdd.n810 avdd.n808 0.713391
R3028 avdd.n808 avdd.n806 0.713391
R3029 avdd.n806 avdd.n804 0.713391
R3030 avdd.n802 avdd.n800 0.713391
R3031 avdd.n800 avdd.n798 0.713391
R3032 avdd.n798 avdd.n796 0.713391
R3033 avdd.n796 avdd.n794 0.713391
R3034 avdd.n794 avdd.n792 0.713391
R3035 avdd.n792 avdd.n556 0.713391
R3036 avdd.n563 avdd.n561 0.713391
R3037 avdd.n565 avdd.n563 0.713391
R3038 avdd.n567 avdd.n565 0.713391
R3039 avdd.n571 avdd.n569 0.713391
R3040 avdd.n573 avdd.n571 0.713391
R3041 avdd.n575 avdd.n573 0.713391
R3042 avdd.n577 avdd.n575 0.713391
R3043 avdd.n579 avdd.n577 0.713391
R3044 avdd.n581 avdd.n579 0.713391
R3045 avdd.n852 avdd.n851 0.713391
R3046 avdd.n851 avdd.n848 0.713391
R3047 avdd.n848 avdd.n814 0.713391
R3048 avdd.n838 avdd.n837 0.713391
R3049 avdd.n837 avdd.n834 0.713391
R3050 avdd.n834 avdd.n816 0.713391
R3051 avdd.n824 avdd.n816 0.713391
R3052 avdd.n824 avdd.n823 0.713391
R3053 avdd.n823 avdd.n820 0.713391
R3054 avdd.n855 avdd.n813 0.713391
R3055 avdd.n845 avdd.n813 0.713391
R3056 avdd.n845 avdd.n844 0.713391
R3057 avdd.n841 avdd.n815 0.713391
R3058 avdd.n831 avdd.n815 0.713391
R3059 avdd.n831 avdd.n830 0.713391
R3060 avdd.n830 avdd.n827 0.713391
R3061 avdd.n827 avdd.n817 0.713391
R3062 avdd.n817 avdd.n599 0.713391
R3063 avdd.n1692 avdd.n1691 0.70362
R3064 avdd.n437 avdd.n435 0.695812
R3065 avdd.n439 avdd.n437 0.695812
R3066 avdd.n441 avdd.n439 0.695812
R3067 avdd.n443 avdd.n441 0.695812
R3068 avdd.n444 avdd.n443 0.695812
R3069 avdd.n861 avdd.n859 0.695812
R3070 avdd.n863 avdd.n861 0.695812
R3071 avdd.n865 avdd.n863 0.695812
R3072 avdd.n867 avdd.n865 0.695812
R3073 avdd.n868 avdd.n867 0.695812
R3074 avdd avdd.n1686 0.664
R3075 avdd.n482 avdd.n480 0.662609
R3076 avdd.n906 avdd.n904 0.662609
R3077 avdd.n1350 avdd.n1349 0.649
R3078 avdd.n1879 avdd.n1878 0.624875
R3079 avdd.n1727 avdd.n525 0.597647
R3080 avdd.n763 avdd 0.576587
R3081 avdd.n1696 avdd 0.563625
R3082 avdd.n961 avdd.n960 0.56281
R3083 avdd.n1703 avdd.n961 0.56281
R3084 avdd.n967 avdd.n952 0.559412
R3085 avdd.n954 avdd.n952 0.559412
R3086 avdd.n1867 avdd.n14 0.55425
R3087 avdd.n1803 avdd.n1802 0.545446
R3088 avdd.n1802 avdd.n1800 0.545446
R3089 avdd.n1800 avdd.n1798 0.545446
R3090 avdd.n1791 avdd.n1788 0.545446
R3091 avdd.n1784 avdd.n1783 0.545446
R3092 avdd.n1728 avdd.n524 0.541125
R3093 avdd.n433 avdd.n389 0.527027
R3094 avdd.n520 avdd.n278 0.527027
R3095 avdd.n856 avdd.n812 0.527027
R3096 avdd.n944 avdd.n526 0.527027
R3097 avdd.n753 avdd.n752 0.526374
R3098 avdd.n754 avdd.n753 0.526374
R3099 avdd.n755 avdd.n754 0.526374
R3100 avdd.n756 avdd.n755 0.526374
R3101 avdd.n757 avdd.n756 0.526374
R3102 avdd.n758 avdd.n757 0.526374
R3103 avdd.n759 avdd.n758 0.49141
R3104 avdd.n499 avdd.n497 0.477062
R3105 avdd.n483 avdd.n308 0.477062
R3106 avdd.n334 avdd.n333 0.477062
R3107 avdd.n397 avdd.n350 0.477062
R3108 avdd.n457 avdd.n351 0.477062
R3109 avdd.n923 avdd.n921 0.477062
R3110 avdd.n907 avdd.n556 0.477062
R3111 avdd.n582 avdd.n581 0.477062
R3112 avdd.n820 avdd.n598 0.477062
R3113 avdd.n881 avdd.n599 0.477062
R3114 avdd.n762 avdd.n760 0.469796
R3115 avdd.n957 avdd.n956 0.444145
R3116 avdd.n956 avdd.n955 0.444145
R3117 avdd.n1725 avdd.n948 0.418878
R3118 avdd.n1729 avdd.n277 0.4145
R3119 avdd.n1697 avdd.n1696 0.407375
R3120 avdd.n763 avdd 0.358608
R3121 avdd avdd.n786 0.357024
R3122 avdd.n1722 avdd.n1721 0.330857
R3123 avdd.n1721 avdd.n1720 0.330857
R3124 avdd.n763 avdd.n762 0.325765
R3125 avdd avdd.n1879 0.32398
R3126 avdd.n497 avdd.n280 0.318859
R3127 avdd.n483 avdd.n482 0.318859
R3128 avdd.n336 avdd.n334 0.318859
R3129 avdd.n461 avdd.n350 0.318859
R3130 avdd.n458 avdd.n457 0.318859
R3131 avdd.n921 avdd.n528 0.318859
R3132 avdd.n907 avdd.n906 0.318859
R3133 avdd.n584 avdd.n582 0.318859
R3134 avdd.n885 avdd.n598 0.318859
R3135 avdd.n882 avdd.n881 0.318859
R3136 avdd.n1792 avdd.n1730 0.316162
R3137 avdd.n1758 avdd.n1756 0.291392
R3138 avdd.n1756 avdd.n1754 0.291392
R3139 avdd.n1778 avdd.n1777 0.284354
R3140 avdd.n1795 avdd.n1794 0.284354
R3141 avdd.n1878 avdd.n14 0.2805
R3142 avdd.n1792 avdd.n1791 0.273291
R3143 avdd.n1806 avdd.n1803 0.272973
R3144 avdd.n1788 avdd.n1784 0.272973
R3145 avdd.n1783 avdd.n1781 0.272973
R3146 avdd.n435 avdd.n434 0.262219
R3147 avdd.n859 avdd.n858 0.262219
R3148 avdd.n781 avdd.n780 0.26137
R3149 avdd.n780 avdd.n779 0.26137
R3150 avdd.n670 avdd.n669 0.26137
R3151 avdd.n670 avdd.n659 0.26137
R3152 avdd.n679 avdd.n659 0.26137
R3153 avdd.n680 avdd.n679 0.26137
R3154 avdd.n681 avdd.n680 0.26137
R3155 avdd.n681 avdd.n654 0.26137
R3156 avdd.n689 avdd.n654 0.26137
R3157 avdd.n690 avdd.n689 0.26137
R3158 avdd.n691 avdd.n690 0.26137
R3159 avdd.n691 avdd.n648 0.26137
R3160 avdd.n700 avdd.n648 0.26137
R3161 avdd.n702 avdd.n701 0.26137
R3162 avdd.n702 avdd.n643 0.26137
R3163 avdd.n710 avdd.n643 0.26137
R3164 avdd.n711 avdd.n710 0.26137
R3165 avdd.n712 avdd.n711 0.26137
R3166 avdd.n712 avdd.n637 0.26137
R3167 avdd.n721 avdd.n637 0.26137
R3168 avdd.n722 avdd.n721 0.26137
R3169 avdd.n723 avdd.n722 0.26137
R3170 avdd.n723 avdd.n632 0.26137
R3171 avdd.n732 avdd.n632 0.26137
R3172 avdd.n733 avdd.n732 0.26137
R3173 avdd.n734 avdd.n733 0.26137
R3174 avdd.n743 avdd.n627 0.26137
R3175 avdd.n744 avdd.n743 0.26137
R3176 avdd.n766 avdd.n744 0.26137
R3177 avdd.n766 avdd.n765 0.26137
R3178 avdd.n765 avdd.n764 0.26137
R3179 avdd.n1729 avdd.n1728 0.2505
R3180 avdd avdd.n250 0.248811
R3181 avdd avdd.n239 0.248811
R3182 avdd.n43 avdd 0.248811
R3183 avdd avdd.n225 0.248811
R3184 avdd avdd.n214 0.248811
R3185 avdd.n63 avdd 0.248811
R3186 avdd avdd.n200 0.248811
R3187 avdd avdd.n189 0.248811
R3188 avdd.n83 avdd 0.248811
R3189 avdd avdd.n175 0.248811
R3190 avdd avdd.n164 0.248811
R3191 avdd.n103 avdd 0.248811
R3192 avdd avdd.n150 0.248811
R3193 avdd avdd.n139 0.248811
R3194 avdd.n123 avdd 0.248811
R3195 avdd.n1748 avdd.n1747 0.246297
R3196 avdd.n1726 avdd 0.242804
R3197 avdd.n1867 avdd.n1866 0.238625
R3198 avdd.n1798 avdd.n1730 0.229784
R3199 avdd.n523 avdd.n520 0.227878
R3200 avdd.n947 avdd.n944 0.227878
R3201 avdd.n1856 avdd.n1835 0.227329
R3202 avdd.n1863 avdd.n1862 0.227329
R3203 avdd.n857 avdd.n856 0.219304
R3204 avdd.n1690 avdd.n1351 0.204245
R3205 avdd.n1691 avdd.n1690 0.195903
R3206 avdd.n1759 avdd.n1758 0.1885
R3207 avdd.n975 avdd.n974 0.1865
R3208 avdd.n1753 avdd.n1751 0.183736
R3209 avdd avdd.n1693 0.178865
R3210 avdd.n14 avdd.n13 0.175331
R3211 avdd.n1830 avdd.n1732 0.156108
R3212 avdd.n474 avdd.n473 0.152959
R3213 avdd.n465 avdd.n464 0.152959
R3214 avdd.n898 avdd.n897 0.152959
R3215 avdd.n889 avdd.n888 0.152959
R3216 avdd.n1715 avdd.n1714 0.152959
R3217 avdd.n760 avdd 0.144186
R3218 avdd.n359 avdd.n358 0.143577
R3219 avdd.n607 avdd.n606 0.143577
R3220 avdd.n354 avdd.n353 0.141409
R3221 avdd.n602 avdd.n601 0.141409
R3222 avdd avdd.n759 0.132362
R3223 avdd.n784 avdd 0.130935
R3224 avdd.n781 avdd 0.130935
R3225 avdd.n779 avdd 0.130935
R3226 avdd avdd.n700 0.130935
R3227 avdd.n701 avdd 0.130935
R3228 avdd.n734 avdd 0.130935
R3229 avdd avdd.n627 0.130935
R3230 avdd.n786 avdd 0.130673
R3231 avdd.n1817 avdd.n1734 0.126176
R3232 avdd.n1822 avdd.n1733 0.126176
R3233 avdd.n1699 avdd.n1698 0.119731
R3234 avdd.n1838 avdd.n1834 0.113554
R3235 avdd.n1840 avdd.n1838 0.113554
R3236 avdd.n1842 avdd.n1840 0.113554
R3237 avdd.n1844 avdd.n1842 0.113554
R3238 avdd.n1846 avdd.n1844 0.113554
R3239 avdd.n1848 avdd.n1846 0.113554
R3240 avdd.n1850 avdd.n1848 0.113554
R3241 avdd.n1851 avdd.n1850 0.113554
R3242 avdd.n1751 avdd.n1750 0.113554
R3243 avdd.n1750 avdd.n1749 0.113554
R3244 avdd.n1793 avdd.n1779 0.0934054
R3245 avdd.n10 avdd.n2 0.0815811
R3246 avdd.n257 avdd.n22 0.0815811
R3247 avdd.n250 avdd.n27 0.0815811
R3248 avdd.n239 avdd.n34 0.0815811
R3249 avdd.n229 avdd.n43 0.0815811
R3250 avdd.n225 avdd.n46 0.0815811
R3251 avdd.n214 avdd.n54 0.0815811
R3252 avdd.n204 avdd.n63 0.0815811
R3253 avdd.n200 avdd.n66 0.0815811
R3254 avdd.n189 avdd.n74 0.0815811
R3255 avdd.n179 avdd.n83 0.0815811
R3256 avdd.n175 avdd.n86 0.0815811
R3257 avdd.n164 avdd.n94 0.0815811
R3258 avdd.n154 avdd.n103 0.0815811
R3259 avdd.n150 avdd.n106 0.0815811
R3260 avdd.n139 avdd.n114 0.0815811
R3261 avdd.n129 avdd.n123 0.0815811
R3262 avdd.n1869 avdd.n21 0.0793136
R3263 avdd.n265 avdd.n16 0.0793136
R3264 avdd.n349 avdd.n348 0.0766719
R3265 avdd.n597 avdd.n596 0.0766719
R3266 avdd.n764 avdd.n763 0.076587
R3267 avdd.n787 avdd 0.0697568
R3268 avdd.n265 avdd.n264 0.0694655
R3269 avdd.n479 avdd.n283 0.0674065
R3270 avdd.n903 avdd.n531 0.0674065
R3271 avdd.n488 avdd.n303 0.0669286
R3272 avdd.n356 avdd.n290 0.0669286
R3273 avdd.n912 avdd.n551 0.0669286
R3274 avdd.n604 avdd.n538 0.0669286
R3275 avdd.n348 avdd.n345 0.0650833
R3276 avdd.n339 avdd.n338 0.0650833
R3277 avdd.n596 avdd.n593 0.0650833
R3278 avdd.n587 avdd.n586 0.0650833
R3279 avdd.n1203 avdd.n1142 0.0579519
R3280 avdd.n1218 avdd.n1121 0.0579519
R3281 avdd.n1233 avdd.n1100 0.0579519
R3282 avdd.n1248 avdd.n1079 0.0579519
R3283 avdd.n1263 avdd.n1058 0.0579519
R3284 avdd.n1278 avdd.n1037 0.0579519
R3285 avdd.n1293 avdd.n1016 0.0579519
R3286 avdd.n1308 avdd.n995 0.0579519
R3287 avdd.n1339 avdd.n1337 0.0579519
R3288 avdd.n1540 avdd.n1515 0.0579519
R3289 avdd.n1555 avdd.n1494 0.0579519
R3290 avdd.n1570 avdd.n1473 0.0579519
R3291 avdd.n1585 avdd.n1452 0.0579519
R3292 avdd.n1600 avdd.n1431 0.0579519
R3293 avdd.n1615 avdd.n1410 0.0579519
R3294 avdd.n1630 avdd.n1389 0.0579519
R3295 avdd.n1645 avdd.n1368 0.0579519
R3296 avdd.n1676 avdd.n1674 0.0579519
R3297 avdd.n1175 avdd.n1168 0.0579519
R3298 avdd.n763 avdd.n616 0.057547
R3299 avdd.n11 avdd.n1 0.0553986
R3300 avdd.n253 avdd.n26 0.0553986
R3301 avdd.n242 avdd.n33 0.0553986
R3302 avdd.n40 avdd.n39 0.0553986
R3303 avdd.n228 avdd.n45 0.0553986
R3304 avdd.n217 avdd.n53 0.0553986
R3305 avdd.n60 avdd.n59 0.0553986
R3306 avdd.n203 avdd.n65 0.0553986
R3307 avdd.n192 avdd.n73 0.0553986
R3308 avdd.n80 avdd.n79 0.0553986
R3309 avdd.n178 avdd.n85 0.0553986
R3310 avdd.n167 avdd.n93 0.0553986
R3311 avdd.n100 avdd.n99 0.0553986
R3312 avdd.n153 avdd.n105 0.0553986
R3313 avdd.n142 avdd.n113 0.0553986
R3314 avdd.n120 avdd.n119 0.0553986
R3315 avdd.n128 avdd.n126 0.0553986
R3316 avdd.n1713 avdd.n1712 0.0527472
R3317 avdd.n789 avdd.n785 0.0516745
R3318 avdd.n1711 avdd.n1710 0.0510435
R3319 avdd.n970 avdd.n966 0.0507703
R3320 avdd.n1770 avdd.n1768 0.0489375
R3321 avdd.n1796 avdd.n1769 0.0489375
R3322 avdd.n1708 avdd.n1707 0.0467687
R3323 avdd.n1879 avdd 0.04675
R3324 avdd.n785 avdd 0.0441242
R3325 avdd.n1754 avdd.n1753 0.0436892
R3326 avdd.n1865 avdd.n1834 0.0430541
R3327 avdd.n1759 avdd.n1748 0.0430541
R3328 avdd.n2 avdd 0.0410405
R3329 avdd avdd.n1344 0.04
R3330 avdd avdd.n1310 0.04
R3331 avdd avdd.n1295 0.04
R3332 avdd avdd.n1280 0.04
R3333 avdd avdd.n1265 0.04
R3334 avdd avdd.n1250 0.04
R3335 avdd avdd.n1235 0.04
R3336 avdd avdd.n1220 0.04
R3337 avdd avdd.n1205 0.04
R3338 avdd avdd.n1681 0.04
R3339 avdd avdd.n1647 0.04
R3340 avdd avdd.n1632 0.04
R3341 avdd avdd.n1617 0.04
R3342 avdd avdd.n1602 0.04
R3343 avdd avdd.n1587 0.04
R3344 avdd avdd.n1572 0.04
R3345 avdd avdd.n1557 0.04
R3346 avdd avdd.n1542 0.04
R3347 avdd avdd.n1177 0.04
R3348 avdd.n1689 avdd 0.038
R3349 avdd.n949 avdd.n277 0.0375
R3350 avdd avdd.n1335 0.0365
R3351 avdd avdd.n1306 0.0365
R3352 avdd avdd.n1291 0.0365
R3353 avdd avdd.n1276 0.0365
R3354 avdd avdd.n1261 0.0365
R3355 avdd avdd.n1246 0.0365
R3356 avdd avdd.n1231 0.0365
R3357 avdd avdd.n1216 0.0365
R3358 avdd avdd.n1201 0.0365
R3359 avdd avdd.n1672 0.0365
R3360 avdd avdd.n1643 0.0365
R3361 avdd avdd.n1628 0.0365
R3362 avdd avdd.n1613 0.0365
R3363 avdd avdd.n1598 0.0365
R3364 avdd avdd.n1583 0.0365
R3365 avdd avdd.n1568 0.0365
R3366 avdd avdd.n1553 0.0365
R3367 avdd avdd.n1538 0.0365
R3368 avdd avdd.n1173 0.0365
R3369 avdd.n252 avdd 0.0351284
R3370 avdd.n241 avdd 0.0351284
R3371 avdd avdd.n42 0.0351284
R3372 avdd.n226 avdd 0.0351284
R3373 avdd.n216 avdd 0.0351284
R3374 avdd avdd.n62 0.0351284
R3375 avdd.n201 avdd 0.0351284
R3376 avdd.n191 avdd 0.0351284
R3377 avdd avdd.n82 0.0351284
R3378 avdd.n176 avdd 0.0351284
R3379 avdd.n166 avdd 0.0351284
R3380 avdd avdd.n102 0.0351284
R3381 avdd.n151 avdd 0.0351284
R3382 avdd.n141 avdd 0.0351284
R3383 avdd avdd.n122 0.0351284
R3384 avdd avdd.n0 0.0351284
R3385 avdd.n978 avdd 0.0335784
R3386 avdd avdd.n1334 0.032
R3387 avdd.n1007 avdd 0.032
R3388 avdd.n1028 avdd 0.032
R3389 avdd.n1049 avdd 0.032
R3390 avdd.n1070 avdd 0.032
R3391 avdd.n1091 avdd 0.032
R3392 avdd.n1112 avdd 0.032
R3393 avdd.n1133 avdd 0.032
R3394 avdd.n1154 avdd 0.032
R3395 avdd avdd.n1671 0.032
R3396 avdd.n1380 avdd 0.032
R3397 avdd.n1401 avdd 0.032
R3398 avdd.n1422 avdd 0.032
R3399 avdd.n1443 avdd 0.032
R3400 avdd.n1464 avdd 0.032
R3401 avdd.n1485 avdd 0.032
R3402 avdd.n1506 avdd 0.032
R3403 avdd.n1527 avdd 0.032
R3404 avdd.n1186 avdd 0.032
R3405 avdd.n965 avdd.n959 0.0301178
R3406 avdd.n969 avdd.n968 0.0300238
R3407 avdd.n1749 avdd.n1732 0.0287635
R3408 avdd.n1724 avdd.n1723 0.0283443
R3409 avdd.n985 avdd 0.028
R3410 avdd.n1358 avdd 0.028
R3411 avdd.n11 avdd.n10 0.0266824
R3412 avdd.n26 avdd.n22 0.0266824
R3413 avdd.n33 avdd.n27 0.0266824
R3414 avdd.n40 avdd.n34 0.0266824
R3415 avdd.n229 avdd.n228 0.0266824
R3416 avdd.n53 avdd.n46 0.0266824
R3417 avdd.n60 avdd.n54 0.0266824
R3418 avdd.n204 avdd.n203 0.0266824
R3419 avdd.n73 avdd.n66 0.0266824
R3420 avdd.n80 avdd.n74 0.0266824
R3421 avdd.n179 avdd.n178 0.0266824
R3422 avdd.n93 avdd.n86 0.0266824
R3423 avdd.n100 avdd.n94 0.0266824
R3424 avdd.n154 avdd.n153 0.0266824
R3425 avdd.n113 avdd.n106 0.0266824
R3426 avdd.n120 avdd.n114 0.0266824
R3427 avdd.n129 avdd.n128 0.0266824
R3428 avdd avdd.n1345 0.0245
R3429 avdd.n1341 avdd 0.0245
R3430 avdd.n1311 avdd 0.0245
R3431 avdd.n996 avdd 0.0245
R3432 avdd.n1296 avdd 0.0245
R3433 avdd.n1017 avdd 0.0245
R3434 avdd.n1281 avdd 0.0245
R3435 avdd.n1038 avdd 0.0245
R3436 avdd.n1266 avdd 0.0245
R3437 avdd.n1059 avdd 0.0245
R3438 avdd.n1251 avdd 0.0245
R3439 avdd.n1080 avdd 0.0245
R3440 avdd.n1236 avdd 0.0245
R3441 avdd.n1101 avdd 0.0245
R3442 avdd.n1221 avdd 0.0245
R3443 avdd.n1122 avdd 0.0245
R3444 avdd.n1206 avdd 0.0245
R3445 avdd.n1143 avdd 0.0245
R3446 avdd.n1678 avdd 0.0245
R3447 avdd.n1648 avdd 0.0245
R3448 avdd.n1369 avdd 0.0245
R3449 avdd.n1633 avdd 0.0245
R3450 avdd.n1390 avdd 0.0245
R3451 avdd.n1618 avdd 0.0245
R3452 avdd.n1411 avdd 0.0245
R3453 avdd.n1603 avdd 0.0245
R3454 avdd.n1432 avdd 0.0245
R3455 avdd.n1588 avdd 0.0245
R3456 avdd.n1453 avdd 0.0245
R3457 avdd.n1573 avdd 0.0245
R3458 avdd.n1474 avdd 0.0245
R3459 avdd.n1558 avdd 0.0245
R3460 avdd.n1495 avdd 0.0245
R3461 avdd.n1543 avdd 0.0245
R3462 avdd.n1516 avdd 0.0245
R3463 avdd.n1172 avdd 0.0245
R3464 avdd.n1709 avdd.n957 0.0240443
R3465 avdd avdd.n1682 0.024
R3466 avdd.n1178 avdd.n1166 0.0235
R3467 avdd.n787 avdd.n785 0.0190811
R3468 avdd.n790 avdd.n789 0.0164396
R3469 avdd avdd.n978 0.0163924
R3470 avdd.n1350 avdd 0.0155
R3471 avdd avdd.n523 0.01225
R3472 avdd avdd.n947 0.01225
R3473 avdd avdd.n1331 0.012
R3474 avdd.n1011 avdd 0.012
R3475 avdd.n1032 avdd 0.012
R3476 avdd.n1053 avdd 0.012
R3477 avdd.n1074 avdd 0.012
R3478 avdd.n1095 avdd 0.012
R3479 avdd.n1116 avdd 0.012
R3480 avdd.n1137 avdd 0.012
R3481 avdd.n1158 avdd 0.012
R3482 avdd avdd.n1668 0.012
R3483 avdd.n1384 avdd 0.012
R3484 avdd.n1405 avdd 0.012
R3485 avdd.n1426 avdd 0.012
R3486 avdd.n1447 avdd 0.012
R3487 avdd.n1468 avdd 0.012
R3488 avdd.n1489 avdd 0.012
R3489 avdd.n1510 avdd 0.012
R3490 avdd.n1531 avdd 0.012
R3491 avdd avdd.n1159 0.012
R3492 avdd.n785 avdd.n784 0.0113696
R3493 avdd.n790 avdd.n616 0.0105671
R3494 avdd.n1349 avdd 0.009
R3495 avdd.n983 avdd 0.009
R3496 avdd.n1345 avdd 0.009
R3497 avdd.n1344 avdd 0.009
R3498 avdd.n1338 avdd 0.009
R3499 avdd.n1335 avdd 0.009
R3500 avdd.n1315 avdd 0.009
R3501 avdd.n1315 avdd 0.009
R3502 avdd.n1332 avdd 0.009
R3503 avdd.n1314 avdd 0.009
R3504 avdd.n1311 avdd 0.009
R3505 avdd.n1310 avdd 0.009
R3506 avdd.n1309 avdd 0.009
R3507 avdd.n1306 avdd 0.009
R3508 avdd avdd.n1302 0.009
R3509 avdd.n1302 avdd 0.009
R3510 avdd avdd.n1010 0.009
R3511 avdd.n1299 avdd 0.009
R3512 avdd.n1296 avdd 0.009
R3513 avdd.n1295 avdd 0.009
R3514 avdd.n1294 avdd 0.009
R3515 avdd.n1291 avdd 0.009
R3516 avdd avdd.n1287 0.009
R3517 avdd.n1287 avdd 0.009
R3518 avdd avdd.n1031 0.009
R3519 avdd.n1284 avdd 0.009
R3520 avdd.n1281 avdd 0.009
R3521 avdd.n1280 avdd 0.009
R3522 avdd.n1279 avdd 0.009
R3523 avdd.n1276 avdd 0.009
R3524 avdd avdd.n1272 0.009
R3525 avdd.n1272 avdd 0.009
R3526 avdd avdd.n1052 0.009
R3527 avdd.n1269 avdd 0.009
R3528 avdd.n1266 avdd 0.009
R3529 avdd.n1265 avdd 0.009
R3530 avdd.n1264 avdd 0.009
R3531 avdd.n1261 avdd 0.009
R3532 avdd avdd.n1257 0.009
R3533 avdd.n1257 avdd 0.009
R3534 avdd avdd.n1073 0.009
R3535 avdd.n1254 avdd 0.009
R3536 avdd.n1251 avdd 0.009
R3537 avdd.n1250 avdd 0.009
R3538 avdd.n1249 avdd 0.009
R3539 avdd.n1246 avdd 0.009
R3540 avdd avdd.n1242 0.009
R3541 avdd.n1242 avdd 0.009
R3542 avdd avdd.n1094 0.009
R3543 avdd.n1239 avdd 0.009
R3544 avdd.n1236 avdd 0.009
R3545 avdd.n1235 avdd 0.009
R3546 avdd.n1234 avdd 0.009
R3547 avdd.n1231 avdd 0.009
R3548 avdd avdd.n1227 0.009
R3549 avdd.n1227 avdd 0.009
R3550 avdd avdd.n1115 0.009
R3551 avdd.n1224 avdd 0.009
R3552 avdd.n1221 avdd 0.009
R3553 avdd.n1220 avdd 0.009
R3554 avdd.n1219 avdd 0.009
R3555 avdd.n1216 avdd 0.009
R3556 avdd avdd.n1212 0.009
R3557 avdd.n1212 avdd 0.009
R3558 avdd avdd.n1136 0.009
R3559 avdd.n1209 avdd 0.009
R3560 avdd.n1206 avdd 0.009
R3561 avdd.n1205 avdd 0.009
R3562 avdd.n1204 avdd 0.009
R3563 avdd.n1201 avdd 0.009
R3564 avdd avdd.n1197 0.009
R3565 avdd.n1197 avdd 0.009
R3566 avdd avdd.n1157 0.009
R3567 avdd.n1688 avdd 0.009
R3568 avdd.n1686 avdd 0.009
R3569 avdd.n1356 avdd 0.009
R3570 avdd.n1682 avdd 0.009
R3571 avdd.n1681 avdd 0.009
R3572 avdd.n1675 avdd 0.009
R3573 avdd.n1672 avdd 0.009
R3574 avdd.n1652 avdd 0.009
R3575 avdd.n1652 avdd 0.009
R3576 avdd.n1669 avdd 0.009
R3577 avdd.n1651 avdd 0.009
R3578 avdd.n1648 avdd 0.009
R3579 avdd.n1647 avdd 0.009
R3580 avdd.n1646 avdd 0.009
R3581 avdd.n1643 avdd 0.009
R3582 avdd avdd.n1639 0.009
R3583 avdd.n1639 avdd 0.009
R3584 avdd avdd.n1383 0.009
R3585 avdd.n1636 avdd 0.009
R3586 avdd.n1633 avdd 0.009
R3587 avdd.n1632 avdd 0.009
R3588 avdd.n1631 avdd 0.009
R3589 avdd.n1628 avdd 0.009
R3590 avdd avdd.n1624 0.009
R3591 avdd.n1624 avdd 0.009
R3592 avdd avdd.n1404 0.009
R3593 avdd.n1621 avdd 0.009
R3594 avdd.n1618 avdd 0.009
R3595 avdd.n1617 avdd 0.009
R3596 avdd.n1616 avdd 0.009
R3597 avdd.n1613 avdd 0.009
R3598 avdd avdd.n1609 0.009
R3599 avdd.n1609 avdd 0.009
R3600 avdd avdd.n1425 0.009
R3601 avdd.n1606 avdd 0.009
R3602 avdd.n1603 avdd 0.009
R3603 avdd.n1602 avdd 0.009
R3604 avdd.n1601 avdd 0.009
R3605 avdd.n1598 avdd 0.009
R3606 avdd avdd.n1594 0.009
R3607 avdd.n1594 avdd 0.009
R3608 avdd avdd.n1446 0.009
R3609 avdd.n1591 avdd 0.009
R3610 avdd.n1588 avdd 0.009
R3611 avdd.n1587 avdd 0.009
R3612 avdd.n1586 avdd 0.009
R3613 avdd.n1583 avdd 0.009
R3614 avdd avdd.n1579 0.009
R3615 avdd.n1579 avdd 0.009
R3616 avdd avdd.n1467 0.009
R3617 avdd.n1576 avdd 0.009
R3618 avdd.n1573 avdd 0.009
R3619 avdd.n1572 avdd 0.009
R3620 avdd.n1571 avdd 0.009
R3621 avdd.n1568 avdd 0.009
R3622 avdd avdd.n1564 0.009
R3623 avdd.n1564 avdd 0.009
R3624 avdd avdd.n1488 0.009
R3625 avdd.n1561 avdd 0.009
R3626 avdd.n1558 avdd 0.009
R3627 avdd.n1557 avdd 0.009
R3628 avdd.n1556 avdd 0.009
R3629 avdd.n1553 avdd 0.009
R3630 avdd avdd.n1549 0.009
R3631 avdd.n1549 avdd 0.009
R3632 avdd avdd.n1509 0.009
R3633 avdd.n1546 avdd 0.009
R3634 avdd.n1543 avdd 0.009
R3635 avdd.n1542 avdd 0.009
R3636 avdd.n1541 avdd 0.009
R3637 avdd.n1538 avdd 0.009
R3638 avdd avdd.n1534 0.009
R3639 avdd.n1534 avdd 0.009
R3640 avdd avdd.n1530 0.009
R3641 avdd.n1178 avdd 0.009
R3642 avdd.n1177 avdd 0.009
R3643 avdd.n1176 avdd 0.009
R3644 avdd.n1173 avdd 0.009
R3645 avdd.n1190 avdd 0.009
R3646 avdd.n1190 avdd 0.009
R3647 avdd.n1189 avdd 0.009
R3648 avdd.n1346 avdd 0.0085
R3649 avdd.n1334 avdd.n989 0.0085
R3650 avdd.n1303 avdd.n1007 0.0085
R3651 avdd.n1288 avdd.n1028 0.0085
R3652 avdd.n1273 avdd.n1049 0.0085
R3653 avdd.n1258 avdd.n1070 0.0085
R3654 avdd.n1243 avdd.n1091 0.0085
R3655 avdd.n1228 avdd.n1112 0.0085
R3656 avdd.n1213 avdd.n1133 0.0085
R3657 avdd.n1198 avdd.n1154 0.0085
R3658 avdd.n1683 avdd 0.0085
R3659 avdd.n1671 avdd.n1362 0.0085
R3660 avdd.n1640 avdd.n1380 0.0085
R3661 avdd.n1625 avdd.n1401 0.0085
R3662 avdd.n1610 avdd.n1422 0.0085
R3663 avdd.n1595 avdd.n1443 0.0085
R3664 avdd.n1580 avdd.n1464 0.0085
R3665 avdd.n1565 avdd.n1485 0.0085
R3666 avdd.n1550 avdd.n1506 0.0085
R3667 avdd.n1535 avdd.n1527 0.0085
R3668 avdd.n1186 avdd.n1185 0.0085
R3669 avdd.n1338 avdd 0.0075
R3670 avdd avdd.n1309 0.0075
R3671 avdd avdd.n1294 0.0075
R3672 avdd avdd.n1279 0.0075
R3673 avdd avdd.n1264 0.0075
R3674 avdd avdd.n1249 0.0075
R3675 avdd avdd.n1234 0.0075
R3676 avdd avdd.n1219 0.0075
R3677 avdd avdd.n1204 0.0075
R3678 avdd.n1675 avdd 0.0075
R3679 avdd avdd.n1646 0.0075
R3680 avdd avdd.n1631 0.0075
R3681 avdd avdd.n1616 0.0075
R3682 avdd avdd.n1601 0.0075
R3683 avdd avdd.n1586 0.0075
R3684 avdd avdd.n1571 0.0075
R3685 avdd avdd.n1556 0.0075
R3686 avdd avdd.n1541 0.0075
R3687 avdd avdd.n1176 0.0075
R3688 avdd.n13 avdd.n1 0.00641216
R3689 avdd.n253 avdd.n252 0.00641216
R3690 avdd.n242 avdd.n241 0.00641216
R3691 avdd.n42 avdd.n39 0.00641216
R3692 avdd.n226 avdd.n45 0.00641216
R3693 avdd.n217 avdd.n216 0.00641216
R3694 avdd.n62 avdd.n59 0.00641216
R3695 avdd.n201 avdd.n65 0.00641216
R3696 avdd.n192 avdd.n191 0.00641216
R3697 avdd.n82 avdd.n79 0.00641216
R3698 avdd.n176 avdd.n85 0.00641216
R3699 avdd.n167 avdd.n166 0.00641216
R3700 avdd.n102 avdd.n99 0.00641216
R3701 avdd.n151 avdd.n105 0.00641216
R3702 avdd.n142 avdd.n141 0.00641216
R3703 avdd.n122 avdd.n119 0.00641216
R3704 avdd.n126 avdd.n0 0.00641216
R3705 avdd.n1340 avdd 0.0055
R3706 avdd.n1331 avdd.n1317 0.0055
R3707 avdd.n1307 avdd 0.0055
R3708 avdd.n1300 avdd.n1011 0.0055
R3709 avdd.n1292 avdd 0.0055
R3710 avdd.n1285 avdd.n1032 0.0055
R3711 avdd.n1277 avdd 0.0055
R3712 avdd.n1270 avdd.n1053 0.0055
R3713 avdd.n1262 avdd 0.0055
R3714 avdd.n1255 avdd.n1074 0.0055
R3715 avdd.n1247 avdd 0.0055
R3716 avdd.n1240 avdd.n1095 0.0055
R3717 avdd.n1232 avdd 0.0055
R3718 avdd.n1225 avdd.n1116 0.0055
R3719 avdd.n1217 avdd 0.0055
R3720 avdd.n1210 avdd.n1137 0.0055
R3721 avdd.n1202 avdd 0.0055
R3722 avdd.n1195 avdd.n1158 0.0055
R3723 avdd.n1677 avdd 0.0055
R3724 avdd.n1668 avdd.n1654 0.0055
R3725 avdd.n1644 avdd 0.0055
R3726 avdd.n1637 avdd.n1384 0.0055
R3727 avdd.n1629 avdd 0.0055
R3728 avdd.n1622 avdd.n1405 0.0055
R3729 avdd.n1614 avdd 0.0055
R3730 avdd.n1607 avdd.n1426 0.0055
R3731 avdd.n1599 avdd 0.0055
R3732 avdd.n1592 avdd.n1447 0.0055
R3733 avdd.n1584 avdd 0.0055
R3734 avdd.n1577 avdd.n1468 0.0055
R3735 avdd.n1569 avdd 0.0055
R3736 avdd.n1562 avdd.n1489 0.0055
R3737 avdd.n1554 avdd 0.0055
R3738 avdd.n1547 avdd.n1510 0.0055
R3739 avdd.n1539 avdd 0.0055
R3740 avdd.n1532 avdd.n1531 0.0055
R3741 avdd.n1174 avdd 0.0055
R3742 avdd.n1192 avdd.n1159 0.0055
R3743 avdd.n1341 avdd.n1340 0.004
R3744 avdd.n1317 avdd 0.004
R3745 avdd.n1307 avdd.n996 0.004
R3746 avdd.n1300 avdd 0.004
R3747 avdd.n1292 avdd.n1017 0.004
R3748 avdd.n1285 avdd 0.004
R3749 avdd.n1277 avdd.n1038 0.004
R3750 avdd.n1270 avdd 0.004
R3751 avdd.n1262 avdd.n1059 0.004
R3752 avdd.n1255 avdd 0.004
R3753 avdd.n1247 avdd.n1080 0.004
R3754 avdd.n1240 avdd 0.004
R3755 avdd.n1232 avdd.n1101 0.004
R3756 avdd.n1225 avdd 0.004
R3757 avdd.n1217 avdd.n1122 0.004
R3758 avdd.n1210 avdd 0.004
R3759 avdd.n1202 avdd.n1143 0.004
R3760 avdd.n1195 avdd 0.004
R3761 avdd.n1678 avdd.n1677 0.004
R3762 avdd.n1654 avdd 0.004
R3763 avdd.n1644 avdd.n1369 0.004
R3764 avdd.n1637 avdd 0.004
R3765 avdd.n1629 avdd.n1390 0.004
R3766 avdd.n1622 avdd 0.004
R3767 avdd.n1614 avdd.n1411 0.004
R3768 avdd.n1607 avdd 0.004
R3769 avdd.n1599 avdd.n1432 0.004
R3770 avdd.n1592 avdd 0.004
R3771 avdd.n1584 avdd.n1453 0.004
R3772 avdd.n1577 avdd 0.004
R3773 avdd.n1569 avdd.n1474 0.004
R3774 avdd.n1562 avdd 0.004
R3775 avdd.n1554 avdd.n1495 0.004
R3776 avdd.n1547 avdd 0.004
R3777 avdd.n1539 avdd.n1516 0.004
R3778 avdd.n1532 avdd 0.004
R3779 avdd.n1174 avdd.n1172 0.004
R3780 avdd avdd.n1192 0.004
R3781 avdd.n983 avdd 0.0035
R3782 avdd.n1356 avdd 0.0035
R3783 avdd.n1332 avdd 0.003
R3784 avdd.n1010 avdd 0.003
R3785 avdd.n1031 avdd 0.003
R3786 avdd.n1052 avdd 0.003
R3787 avdd.n1073 avdd 0.003
R3788 avdd.n1094 avdd 0.003
R3789 avdd.n1115 avdd 0.003
R3790 avdd.n1136 avdd 0.003
R3791 avdd.n1157 avdd 0.003
R3792 avdd.n1669 avdd 0.003
R3793 avdd.n1383 avdd 0.003
R3794 avdd.n1404 avdd 0.003
R3795 avdd.n1425 avdd 0.003
R3796 avdd.n1446 avdd 0.003
R3797 avdd.n1467 avdd 0.003
R3798 avdd.n1488 avdd 0.003
R3799 avdd.n1509 avdd 0.003
R3800 avdd.n1530 avdd 0.003
R3801 avdd avdd.n1189 0.003
R3802 avdd.n1689 avdd.n1688 0.0025
R3803 avdd.n1346 avdd.n985 0.001
R3804 avdd avdd.n989 0.001
R3805 avdd.n1303 avdd 0.001
R3806 avdd.n1288 avdd 0.001
R3807 avdd.n1273 avdd 0.001
R3808 avdd.n1258 avdd 0.001
R3809 avdd.n1243 avdd 0.001
R3810 avdd.n1228 avdd 0.001
R3811 avdd.n1213 avdd 0.001
R3812 avdd.n1198 avdd 0.001
R3813 avdd.n1683 avdd.n1358 0.001
R3814 avdd avdd.n1362 0.001
R3815 avdd.n1640 avdd 0.001
R3816 avdd.n1625 avdd 0.001
R3817 avdd.n1610 avdd 0.001
R3818 avdd.n1595 avdd 0.001
R3819 avdd.n1580 avdd 0.001
R3820 avdd.n1565 avdd 0.001
R3821 avdd.n1550 avdd 0.001
R3822 avdd.n1535 avdd 0.001
R3823 avdd.n1185 avdd 0.001
R3824 por_ana_0.ibias_gen_0.vp0.n3 por_ana_0.ibias_gen_0.vp0.n1 57.7416
R3825 por_ana_0.ibias_gen_0.vp0.n8 por_ana_0.ibias_gen_0.vp0.t12 50.9767
R3826 por_ana_0.ibias_gen_0.vp0.t12 por_ana_0.ibias_gen_0.vp0.n6 50.9767
R3827 por_ana_0.ibias_gen_0.vp0.n7 por_ana_0.ibias_gen_0.vp0.t3 49.8109
R3828 por_ana_0.ibias_gen_0.vp0.n0 por_ana_0.ibias_gen_0.vp0.t3 49.7239
R3829 por_ana_0.ibias_gen_0.vp0.t1 por_ana_0.ibias_gen_0.vp0.n9 48.6451
R3830 por_ana_0.ibias_gen_0.vp0.t13 por_ana_0.ibias_gen_0.vp0.n6 48.6451
R3831 por_ana_0.ibias_gen_0.vp0.n10 por_ana_0.ibias_gen_0.vp0.t1 48.6451
R3832 por_ana_0.ibias_gen_0.vp0.n8 por_ana_0.ibias_gen_0.vp0.t13 48.6451
R3833 por_ana_0.ibias_gen_0.vp0.n5 por_ana_0.ibias_gen_0.vp0.n4 42.4505
R3834 por_ana_0.ibias_gen_0.vp0.n3 por_ana_0.ibias_gen_0.vp0.n2 42.4505
R3835 por_ana_0.ibias_gen_0.vp0.n14 por_ana_0.ibias_gen_0.vp0.n13 18.2113
R3836 por_ana_0.ibias_gen_0.vp0.n12 por_ana_0.ibias_gen_0.vp0.n11 17.2812
R3837 por_ana_0.ibias_gen_0.vp0.n10 por_ana_0.ibias_gen_0.vp0.n6 13.7361
R3838 por_ana_0.ibias_gen_0.vp0.n9 por_ana_0.ibias_gen_0.vp0.n8 13.7361
R3839 por_ana_0.ibias_gen_0.vp0.n13 por_ana_0.ibias_gen_0.vp0.n12 13.3639
R3840 por_ana_0.ibias_gen_0.vp0.n4 por_ana_0.ibias_gen_0.vp0.t4 5.5395
R3841 por_ana_0.ibias_gen_0.vp0.n4 por_ana_0.ibias_gen_0.vp0.t2 5.5395
R3842 por_ana_0.ibias_gen_0.vp0.n2 por_ana_0.ibias_gen_0.vp0.t10 5.5395
R3843 por_ana_0.ibias_gen_0.vp0.n2 por_ana_0.ibias_gen_0.vp0.t0 5.5395
R3844 por_ana_0.ibias_gen_0.vp0.n1 por_ana_0.ibias_gen_0.vp0.t9 5.5395
R3845 por_ana_0.ibias_gen_0.vp0.n1 por_ana_0.ibias_gen_0.vp0.t11 5.5395
R3846 por_ana_0.ibias_gen_0.vp0.n13 por_ana_0.ibias_gen_0.vp0.n3 3.97054
R3847 por_ana_0.ibias_gen_0.vp0.n12 por_ana_0.ibias_gen_0.vp0.n0 3.77198
R3848 por_ana_0.ibias_gen_0.vp0.n11 por_ana_0.ibias_gen_0.vp0.t7 3.3065
R3849 por_ana_0.ibias_gen_0.vp0.n11 por_ana_0.ibias_gen_0.vp0.t6 3.3065
R3850 por_ana_0.ibias_gen_0.vp0.n14 por_ana_0.ibias_gen_0.vp0.t8 3.3065
R3851 por_ana_0.ibias_gen_0.vp0.t5 por_ana_0.ibias_gen_0.vp0.n14 3.3065
R3852 por_ana_0.ibias_gen_0.vp0.n7 por_ana_0.ibias_gen_0.vp0.n5 1.47061
R3853 por_ana_0.ibias_gen_0.vp0.n0 por_ana_0.ibias_gen_0.vp0.n10 1.3293
R3854 por_ana_0.ibias_gen_0.vp0.n9 por_ana_0.ibias_gen_0.vp0.n7 1.16626
R3855 por_ana_0.ibias_gen_0.vp0.n0 por_ana_0.ibias_gen_0.vp0.n5 1.13637
R3856 por_ana_0.ibias_gen_0.vn0.n9 por_ana_0.ibias_gen_0.vn0.t19 50.4613
R3857 por_ana_0.ibias_gen_0.vn0.n10 por_ana_0.ibias_gen_0.vn0.t19 50.4344
R3858 por_ana_0.ibias_gen_0.vn0.n1 por_ana_0.ibias_gen_0.vn0.n7 49.6079
R3859 por_ana_0.ibias_gen_0.vn0.n4 por_ana_0.ibias_gen_0.vn0.t2 49.2687
R3860 por_ana_0.ibias_gen_0.vn0.n1 por_ana_0.ibias_gen_0.vn0.t2 49.1817
R3861 por_ana_0.ibias_gen_0.vn0.t4 por_ana_0.ibias_gen_0.vn0.n3 48.1029
R3862 por_ana_0.ibias_gen_0.vn0.t20 por_ana_0.ibias_gen_0.vn0.n9 48.1029
R3863 por_ana_0.ibias_gen_0.vn0.n8 por_ana_0.ibias_gen_0.vn0.t4 48.1029
R3864 por_ana_0.ibias_gen_0.vn0.n10 por_ana_0.ibias_gen_0.vn0.t20 48.1029
R3865 por_ana_0.ibias_gen_0.vn0.n0 por_ana_0.ibias_gen_0.vn0.t14 22.9447
R3866 por_ana_0.ibias_gen_0.Mt4 por_ana_0.ibias_gen_0.vn0.n2 21.105
R3867 por_ana_0.ibias_gen_0.vn0.n0 por_ana_0.ibias_gen_0.vn0.n13 19.6387
R3868 por_ana_0.ibias_gen_0.Mt4 por_ana_0.ibias_gen_0.vn0.n14 19.6387
R3869 por_ana_0.ibias_gen_0.Mt4 por_ana_0.ibias_gen_0.vn0.n15 19.6387
R3870 por_ana_0.ibias_gen_0.Mt4 por_ana_0.ibias_gen_0.vn0.n16 19.6387
R3871 por_ana_0.ibias_gen_0.vn0.n0 por_ana_0.ibias_gen_0.vn0.n12 19.6387
R3872 por_ana_0.ibias_gen_0.vn0.n6 por_ana_0.ibias_gen_0.vn0.n5 13.8791
R3873 por_ana_0.ibias_gen_0.vn0.n9 por_ana_0.ibias_gen_0.vn0.n8 13.7174
R3874 por_ana_0.ibias_gen_0.vn0.n0 por_ana_0.ibias_gen_0.vn0.n11 12.7887
R3875 por_ana_0.ibias_gen_0.vn0.n11 por_ana_0.ibias_gen_0.vn0.n3 7.26784
R3876 por_ana_0.ibias_gen_0.vn0.n11 por_ana_0.ibias_gen_0.vn0.n10 6.45004
R3877 por_ana_0.ibias_gen_0.vn0.n7 por_ana_0.ibias_gen_0.vn0.t0 5.5395
R3878 por_ana_0.ibias_gen_0.vn0.n7 por_ana_0.ibias_gen_0.vn0.t1 5.5395
R3879 por_ana_0.ibias_gen_0.vn0.n5 por_ana_0.ibias_gen_0.vn0.t5 3.3065
R3880 por_ana_0.ibias_gen_0.vn0.n5 por_ana_0.ibias_gen_0.vn0.t3 3.3065
R3881 por_ana_0.ibias_gen_0.vn0.n13 por_ana_0.ibias_gen_0.vn0.t7 3.3065
R3882 por_ana_0.ibias_gen_0.vn0.n13 por_ana_0.ibias_gen_0.vn0.t9 3.3065
R3883 por_ana_0.ibias_gen_0.vn0.n14 por_ana_0.ibias_gen_0.vn0.t12 3.3065
R3884 por_ana_0.ibias_gen_0.vn0.n14 por_ana_0.ibias_gen_0.vn0.t15 3.3065
R3885 por_ana_0.ibias_gen_0.vn0.n15 por_ana_0.ibias_gen_0.vn0.t13 3.3065
R3886 por_ana_0.ibias_gen_0.vn0.n15 por_ana_0.ibias_gen_0.vn0.t10 3.3065
R3887 por_ana_0.ibias_gen_0.vn0.n16 por_ana_0.ibias_gen_0.vn0.t16 3.3065
R3888 por_ana_0.ibias_gen_0.vn0.n16 por_ana_0.ibias_gen_0.vn0.t11 3.3065
R3889 por_ana_0.ibias_gen_0.vn0.n2 por_ana_0.ibias_gen_0.vn0.t18 3.3065
R3890 por_ana_0.ibias_gen_0.vn0.n2 por_ana_0.ibias_gen_0.vn0.t17 3.3065
R3891 por_ana_0.ibias_gen_0.vn0.n12 por_ana_0.ibias_gen_0.vn0.t6 3.3065
R3892 por_ana_0.ibias_gen_0.vn0.n12 por_ana_0.ibias_gen_0.vn0.t8 3.3065
R3893 por_ana_0.ibias_gen_0.Mt4 por_ana_0.ibias_gen_0.vn0.n0 2.11628
R3894 por_ana_0.ibias_gen_0.vn0.n6 por_ana_0.ibias_gen_0.vn0.n4 1.44615
R3895 por_ana_0.ibias_gen_0.vn0.n8 por_ana_0.ibias_gen_0.vn0.n1 1.30001
R3896 por_ana_0.ibias_gen_0.vn0.n4 por_ana_0.ibias_gen_0.vn0.n3 1.16626
R3897 por_ana_0.ibias_gen_0.vn0.n1 por_ana_0.ibias_gen_0.vn0.n6 1.15267
R3898 dvdd.n3109 dvdd.n3107 53399.3
R3899 dvdd.n3111 dvdd.n3107 53399.3
R3900 dvdd.n3111 dvdd.n3110 53399.3
R3901 dvdd.n3110 dvdd.n3109 53399.3
R3902 dvdd.n3108 dvdd.n3106 26464.9
R3903 dvdd.n3112 dvdd.n3106 26464.9
R3904 dvdd.n3112 dvdd.n3104 26464.9
R3905 dvdd.n3108 dvdd.n3104 26464.9
R3906 dvdd.n2935 dvdd.n2933 15977.3
R3907 dvdd.n2937 dvdd.n2933 15974
R3908 dvdd.n2936 dvdd.n2935 15974
R3909 dvdd.n2937 dvdd.n2936 15970.6
R3910 dvdd.n3142 dvdd.n3139 8474.12
R3911 dvdd.n3144 dvdd.n3139 8474.12
R3912 dvdd.n3142 dvdd.n3141 8470.59
R3913 dvdd.n3144 dvdd.n3141 8470.59
R3914 dvdd.n2934 dvdd.n2931 8195.68
R3915 dvdd.n2934 dvdd.n2932 8194.05
R3916 dvdd.n2938 dvdd.n2931 8194.05
R3917 dvdd.n2938 dvdd.n2932 8192.43
R3918 dvdd.n3105 dvdd.n3103 6151.53
R3919 dvdd.n3114 dvdd.n3103 6151.53
R3920 dvdd.n3113 dvdd.n3105 6151.53
R3921 dvdd.n3114 dvdd.n3113 6151.53
R3922 dvdd.n2963 dvdd.n2962 4782.35
R3923 dvdd.n2964 dvdd.n2962 4782.35
R3924 dvdd.n2963 dvdd.n2947 4782.35
R3925 dvdd.n2964 dvdd.n2947 4782.35
R3926 dvdd.n2940 dvdd.n2930 1910.21
R3927 dvdd.n2930 dvdd.n2929 1909.84
R3928 dvdd.n2940 dvdd.n2939 1909.84
R3929 dvdd.n2939 dvdd.n2929 1909.46
R3930 dvdd.t1802 dvdd 1725.39
R3931 dvdd dvdd.t1673 1725.39
R3932 dvdd.t1768 dvdd 1719.47
R3933 dvdd dvdd.t1564 1719.47
R3934 dvdd dvdd.t1745 1719.47
R3935 dvdd.n409 dvdd.n407 1718.5
R3936 dvdd dvdd.t1802 1547.82
R3937 dvdd dvdd.t1768 1547.82
R3938 dvdd.t1564 dvdd 1547.82
R3939 dvdd.t1673 dvdd 1547.82
R3940 dvdd.t1745 dvdd 1547.82
R3941 dvdd.t1623 dvdd 1174.92
R3942 dvdd dvdd.t1623 1003.27
R3943 dvdd.t1537 dvdd 978.534
R3944 dvdd dvdd.t1593 975.178
R3945 dvdd dvdd.t1707 975.178
R3946 dvdd.n3147 dvdd.n3138 903.907
R3947 dvdd.n3145 dvdd.n3140 903.529
R3948 dvdd.n3140 dvdd.n3138 903.529
R3949 dvdd dvdd.t1537 877.827
R3950 dvdd.t1593 dvdd 877.827
R3951 dvdd.t1707 dvdd 877.827
R3952 dvdd.n348 dvdd.t1326 873.438
R3953 dvdd.n2920 dvdd.t712 871.962
R3954 dvdd.n3074 dvdd.t688 871.962
R3955 dvdd.n3017 dvdd.t994 871.962
R3956 dvdd.n2863 dvdd.t692 871.962
R3957 dvdd.n2809 dvdd.t187 871.962
R3958 dvdd.n761 dvdd.t862 871.529
R3959 dvdd.n2031 dvdd.t980 870.355
R3960 dvdd.n3146 dvdd.n3145 857.977
R3961 dvdd.n2352 dvdd.t907 842.716
R3962 dvdd.n2110 dvdd.t306 842.073
R3963 dvdd.n928 dvdd.t887 836.124
R3964 dvdd.n1322 dvdd.t581 836.124
R3965 dvdd.n2127 dvdd.t1322 832.876
R3966 dvdd.n1342 dvdd.t1331 830.703
R3967 dvdd.t24 dvdd.t1807 822.741
R3968 dvdd.n2268 dvdd.t1559 809.372
R3969 dvdd.n2401 dvdd.t1663 809.322
R3970 dvdd.n362 dvdd.t1790 807.567
R3971 dvdd.n643 dvdd.t1689 807.567
R3972 dvdd.n2484 dvdd.t1742 807.548
R3973 dvdd.n432 dvdd.t1782 807.481
R3974 dvdd.n705 dvdd.t1800 807.481
R3975 dvdd.n726 dvdd.t647 806.537
R3976 dvdd.n460 dvdd.t822 806.511
R3977 dvdd.n1007 dvdd.t1078 806.511
R3978 dvdd.n1444 dvdd.t1129 806.511
R3979 dvdd.n1887 dvdd.t227 806.511
R3980 dvdd.n1817 dvdd.t1068 806.511
R3981 dvdd.n2175 dvdd.t1753 806.484
R3982 dvdd.n865 dvdd.t1720 806.423
R3983 dvdd.n222 dvdd.t1675 804.731
R3984 dvdd.n275 dvdd.t1674 804.731
R3985 dvdd.n229 dvdd.t1747 804.731
R3986 dvdd.n223 dvdd.t1746 804.731
R3987 dvdd.n319 dvdd.t1566 804.731
R3988 dvdd.n300 dvdd.t1565 804.731
R3989 dvdd.n156 dvdd.t1804 804.731
R3990 dvdd.n162 dvdd.t1803 804.731
R3991 dvdd.n105 dvdd.t1770 804.731
R3992 dvdd.n100 dvdd.t1769 804.731
R3993 dvdd.n546 dvdd.t1764 804.731
R3994 dvdd.n540 dvdd.t1763 804.731
R3995 dvdd.n546 dvdd.t1595 804.731
R3996 dvdd.n540 dvdd.t1594 804.731
R3997 dvdd.n455 dvdd.t1791 804.731
R3998 dvdd.n431 dvdd.t1651 804.731
R3999 dvdd.n416 dvdd.t1781 804.731
R4000 dvdd.n369 dvdd.t1650 804.731
R4001 dvdd.n370 dvdd.t1539 804.731
R4002 dvdd.n376 dvdd.t1538 804.731
R4003 dvdd.n370 dvdd.t1677 804.731
R4004 dvdd.n376 dvdd.t1676 804.731
R4005 dvdd.n379 dvdd.t1648 804.731
R4006 dvdd.n382 dvdd.t1749 804.731
R4007 dvdd.n537 dvdd.t1697 804.731
R4008 dvdd.n549 dvdd.t1668 804.731
R4009 dvdd.n552 dvdd.t1760 804.731
R4010 dvdd.n650 dvdd.t1688 804.731
R4011 dvdd.n636 dvdd.t1801 804.731
R4012 dvdd.n658 dvdd.t1542 804.731
R4013 dvdd.n662 dvdd.t1686 804.731
R4014 dvdd.n835 dvdd.t1709 804.731
R4015 dvdd.n829 dvdd.t1708 804.731
R4016 dvdd.n835 dvdd.t1793 804.731
R4017 dvdd.n829 dvdd.t1792 804.731
R4018 dvdd.n827 dvdd.t1608 804.731
R4019 dvdd.n879 dvdd.t1719 804.731
R4020 dvdd.n838 dvdd.t1563 804.731
R4021 dvdd.n841 dvdd.t1704 804.731
R4022 dvdd.n956 dvdd.t1744 804.731
R4023 dvdd.n959 dvdd.t1580 804.731
R4024 dvdd.n1125 dvdd.t1756 804.731
R4025 dvdd.n1128 dvdd.t1611 804.731
R4026 dvdd.n1229 dvdd.t1571 804.731
R4027 dvdd.n1236 dvdd.t1570 804.731
R4028 dvdd.n1259 dvdd.t1589 804.731
R4029 dvdd.n1262 dvdd.t1585 804.731
R4030 dvdd.n1416 dvdd.t1627 804.731
R4031 dvdd.n1419 dvdd.t1614 804.731
R4032 dvdd.n1546 dvdd.t1602 804.731
R4033 dvdd.n1550 dvdd.t1788 804.731
R4034 dvdd.n1527 dvdd.t1544 804.731
R4035 dvdd.n1709 dvdd.t1630 804.731
R4036 dvdd.n1712 dvdd.t1806 804.731
R4037 dvdd.n2007 dvdd.t1735 804.731
R4038 dvdd.n2062 dvdd.t1734 804.731
R4039 dvdd.n1864 dvdd.t1639 804.731
R4040 dvdd.n1843 dvdd.t1638 804.731
R4041 dvdd.n1835 dvdd.t1795 804.731
R4042 dvdd.n1838 dvdd.t1723 804.731
R4043 dvdd.n1997 dvdd.t1654 804.731
R4044 dvdd.n2020 dvdd.t1536 804.731
R4045 dvdd.n2023 dvdd.t1739 804.731
R4046 dvdd.n2142 dvdd.t1706 804.731
R4047 dvdd.n2262 dvdd.t1762 804.731
R4048 dvdd.n2235 dvdd.t1761 804.731
R4049 dvdd.n2262 dvdd.t1694 804.731
R4050 dvdd.n2235 dvdd.t1693 804.731
R4051 dvdd.n2238 dvdd.t1558 804.731
R4052 dvdd.n2241 dvdd.t1758 804.731
R4053 dvdd.n2183 dvdd.t1786 804.731
R4054 dvdd.n2180 dvdd.t1754 804.731
R4055 dvdd.n2220 dvdd.t1785 804.731
R4056 dvdd.n2167 dvdd.t1587 804.731
R4057 dvdd.t1716 dvdd.n2169 804.731
R4058 dvdd.n2285 dvdd.t1560 804.731
R4059 dvdd.n2139 dvdd.t1776 804.731
R4060 dvdd.n2291 dvdd.t1736 804.731
R4061 dvdd.n2133 dvdd.t1777 804.731
R4062 dvdd.n2128 dvdd.t1737 804.731
R4063 dvdd.n2132 dvdd.t1567 804.731
R4064 dvdd.n2317 dvdd.t1568 804.731
R4065 dvdd.t1698 dvdd.n2104 804.731
R4066 dvdd.n2109 dvdd.t1524 804.731
R4067 dvdd.n2190 dvdd.t1582 804.731
R4068 dvdd.n2193 dvdd.t1779 804.731
R4069 dvdd.n2467 dvdd.t1741 804.731
R4070 dvdd.n2394 dvdd.t1797 804.731
R4071 dvdd.n2476 dvdd.t1555 804.731
R4072 dvdd.n2513 dvdd.t1775 804.731
R4073 dvdd.n2382 dvdd.t1527 804.731
R4074 dvdd.n2460 dvdd.t1657 804.731
R4075 dvdd.n2441 dvdd.t1662 804.731
R4076 dvdd.n2405 dvdd.t1592 804.731
R4077 dvdd.n2411 dvdd.t1591 804.731
R4078 dvdd.n2414 dvdd.t1772 804.731
R4079 dvdd.n2417 dvdd.t1702 804.731
R4080 dvdd.n2583 dvdd.t1784 804.731
R4081 dvdd.n2586 dvdd.t1712 804.731
R4082 dvdd.n885 dvdd.t1036 804.095
R4083 dvdd.n349 dvdd.t1194 803.572
R4084 dvdd.n1009 dvdd.t922 803.572
R4085 dvdd.n1056 dvdd.t1320 803.572
R4086 dvdd.n1148 dvdd.t992 803.572
R4087 dvdd.n1297 dvdd.t796 803.572
R4088 dvdd.n1390 dvdd.t527 803.572
R4089 dvdd.n1502 dvdd.t1094 803.572
R4090 dvdd.n1735 dvdd.t1510 803.572
R4091 dvdd.n1700 dvdd.t181 803.572
R4092 dvdd.n1966 dvdd.t1123 803.572
R4093 dvdd.n2060 dvdd.t820 803.572
R4094 dvdd.n727 dvdd.t499 783.403
R4095 dvdd.n1381 dvdd.t109 783.403
R4096 dvdd.n1798 dvdd.t149 780.84
R4097 dvdd.n1208 dvdd.t911 770.25
R4098 dvdd.t1544 dvdd.n1526 751.692
R4099 dvdd.t1587 dvdd.n2166 751.692
R4100 dvdd.n2170 dvdd.t1716 751.692
R4101 dvdd.n2153 dvdd.t1698 751.692
R4102 dvdd.t1648 dvdd.n378 725.173
R4103 dvdd.t1749 dvdd.n381 725.173
R4104 dvdd.t1697 dvdd.n536 725.173
R4105 dvdd.t1668 dvdd.n548 725.173
R4106 dvdd.t1760 dvdd.n551 725.173
R4107 dvdd.t1542 dvdd.n657 725.173
R4108 dvdd.t1686 dvdd.n661 725.173
R4109 dvdd.t1608 dvdd.n826 725.173
R4110 dvdd.t1563 dvdd.n837 725.173
R4111 dvdd.t1704 dvdd.n840 725.173
R4112 dvdd.t1744 dvdd.n955 725.173
R4113 dvdd.t1580 dvdd.n958 725.173
R4114 dvdd.t1756 dvdd.n1124 725.173
R4115 dvdd.t1611 dvdd.n1127 725.173
R4116 dvdd.t1589 dvdd.n1258 725.173
R4117 dvdd.t1585 dvdd.n1261 725.173
R4118 dvdd.t1627 dvdd.n1415 725.173
R4119 dvdd.t1614 dvdd.n1418 725.173
R4120 dvdd.t1602 dvdd.n1545 725.173
R4121 dvdd.t1788 dvdd.n1549 725.173
R4122 dvdd.t1630 dvdd.n1708 725.173
R4123 dvdd.t1806 dvdd.n1711 725.173
R4124 dvdd.t1795 dvdd.n1834 725.173
R4125 dvdd.t1723 dvdd.n1837 725.173
R4126 dvdd.t1654 dvdd.n1996 725.173
R4127 dvdd.t1536 dvdd.n2019 725.173
R4128 dvdd.t1739 dvdd.n2022 725.173
R4129 dvdd.t1706 dvdd.n2141 725.173
R4130 dvdd.t1558 dvdd.n2237 725.173
R4131 dvdd.t1758 dvdd.n2240 725.173
R4132 dvdd.t1524 dvdd.n2108 725.173
R4133 dvdd.t1582 dvdd.n2189 725.173
R4134 dvdd.t1779 dvdd.n2192 725.173
R4135 dvdd.t1797 dvdd.n2393 725.173
R4136 dvdd.t1555 dvdd.n2475 725.173
R4137 dvdd.t1775 dvdd.n2512 725.173
R4138 dvdd.t1527 dvdd.n2381 725.173
R4139 dvdd.t1657 dvdd.n2459 725.173
R4140 dvdd.t1772 dvdd.n2413 725.173
R4141 dvdd.t1702 dvdd.n2416 725.173
R4142 dvdd.t1784 dvdd.n2582 725.173
R4143 dvdd.t1712 dvdd.n2585 725.173
R4144 dvdd.n2500 dvdd.n2388 721.278
R4145 dvdd.n2546 dvdd.n2514 721.278
R4146 dvdd.n2550 dvdd.n2504 720.484
R4147 dvdd.n1063 dvdd.n1062 717.729
R4148 dvdd.n1219 dvdd.n1218 717.729
R4149 dvdd.n1288 dvdd.n1243 717.729
R4150 dvdd.n2550 dvdd.n2505 717.729
R4151 dvdd.n466 dvdd.n465 713.462
R4152 dvdd.n1373 dvdd.n1330 713.462
R4153 dvdd.n2012 dvdd.t1182 699.619
R4154 dvdd.t760 dvdd.t1713 689.564
R4155 dvdd.n1102 dvdd.t89 671.408
R4156 dvdd.n1575 dvdd.t1242 671.408
R4157 dvdd dvdd.t1649 669.701
R4158 dvdd.n2536 dvdd.t1441 669.491
R4159 dvdd.n582 dvdd.t7 667.778
R4160 dvdd.n1021 dvdd.t782 667.778
R4161 dvdd.n1023 dvdd.t924 667.778
R4162 dvdd.n1048 dvdd.t517 667.778
R4163 dvdd.n1160 dvdd.t1222 667.778
R4164 dvdd.n1445 dvdd.t1328 667.778
R4165 dvdd.n1669 dvdd.t312 667.778
R4166 dvdd.n1815 dvdd.t663 667.778
R4167 dvdd.n604 dvdd.t371 667.751
R4168 dvdd.n1080 dvdd.t1151 667.751
R4169 dvdd.n1120 dvdd.t720 667.751
R4170 dvdd.n1507 dvdd.t1412 667.751
R4171 dvdd.n1747 dvdd.t1098 667.751
R4172 dvdd.n1720 dvdd.t1086 667.751
R4173 dvdd.n1882 dvdd.t1211 667.751
R4174 dvdd.n2489 dvdd.t680 667.672
R4175 dvdd.n1433 dvdd.t1190 666.774
R4176 dvdd.n1290 dvdd.t1137 666.254
R4177 dvdd.n2547 dvdd.t747 666.206
R4178 dvdd.n2068 dvdd.t909 665.715
R4179 dvdd.t1765 dvdd 664.664
R4180 dvdd.n447 dvdd.t1508 664.455
R4181 dvdd.n715 dvdd.t571 664.455
R4182 dvdd.n905 dvdd.t637 664.455
R4183 dvdd.n993 dvdd.t792 664.455
R4184 dvdd.n1000 dvdd.t521 664.455
R4185 dvdd.n1467 dvdd.t639 664.455
R4186 dvdd.n1453 dvdd.t807 664.455
R4187 dvdd.n1875 dvdd.t97 664.455
R4188 dvdd.n1933 dvdd.t318 664.455
R4189 dvdd.n514 dvdd.t573 663.426
R4190 dvdd.n629 dvdd.t525 663.426
R4191 dvdd.n872 dvdd.t324 663.426
R4192 dvdd.n1310 dvdd.t1300 663.426
R4193 dvdd.n1691 dvdd.t529 663.426
R4194 dvdd.n1722 dvdd.t1020 663.426
R4195 dvdd.n1813 dvdd.t1008 663.426
R4196 dvdd.n1951 dvdd.t1486 663.426
R4197 dvdd.n2048 dvdd.t1016 663.426
R4198 dvdd.n1274 dvdd.t505 662.841
R4199 dvdd.n1593 dvdd.t1147 661.644
R4200 dvdd.n777 dvdd.t1164 659.593
R4201 dvdd.n795 dvdd.n760 629.801
R4202 dvdd.n1380 dvdd.n1327 620.338
R4203 dvdd.n2548 dvdd.n2506 615.659
R4204 dvdd.n2494 dvdd.n2491 613.89
R4205 dvdd.n1069 dvdd.n1065 611.646
R4206 dvdd.n1221 dvdd.n1220 611.178
R4207 dvdd.n1290 dvdd.n1240 611.178
R4208 dvdd.n2548 dvdd.n2508 611.149
R4209 dvdd.n1371 dvdd.n1331 611.122
R4210 dvdd.n1369 dvdd.n1335 611.122
R4211 dvdd.n1946 dvdd.n1945 611.122
R4212 dvdd.n1794 dvdd.n1793 611.122
R4213 dvdd.n737 dvdd.n736 610.861
R4214 dvdd.n745 dvdd.n744 610.861
R4215 dvdd.n1380 dvdd.n1378 610.098
R4216 dvdd.n2081 dvdd.n1796 610.098
R4217 dvdd.n511 dvdd.n469 609.847
R4218 dvdd.n731 dvdd.n730 609.847
R4219 dvdd.n1367 dvdd.n1339 609.615
R4220 dvdd.n1357 dvdd.n1344 609.615
R4221 dvdd.n1941 dvdd.n1940 609.615
R4222 dvdd.n1959 dvdd.n1944 609.615
R4223 dvdd.n85 dvdd.n84 608.631
R4224 dvdd.n1195 dvdd.n921 608.631
R4225 dvdd.n1255 dvdd.n1254 608.631
R4226 dvdd.n2113 dvdd.n2112 607.155
R4227 dvdd.n2561 dvdd.n2560 607.155
R4228 dvdd.n2626 dvdd.n2562 607.155
R4229 dvdd.n739 dvdd.n631 606.42
R4230 dvdd.n1374 dvdd.n1329 606.42
R4231 dvdd.n1952 dvdd.n1948 606.42
R4232 dvdd.n1322 dvdd.n1223 606.299
R4233 dvdd.n748 dvdd.n747 605.186
R4234 dvdd.n627 dvdd.n626 605.186
R4235 dvdd.n755 dvdd.n754 605.186
R4236 dvdd.n1362 dvdd.n1341 605.186
R4237 dvdd.n1968 dvdd.n1939 605.186
R4238 dvdd.n603 dvdd.n338 604.457
R4239 dvdd.n602 dvdd.n339 604.457
R4240 dvdd.n621 dvdd.n620 604.457
R4241 dvdd.n1003 dvdd.n1002 604.457
R4242 dvdd.n1082 dvdd.n1059 604.457
R4243 dvdd.n1139 dvdd.n1119 604.457
R4244 dvdd.n1291 dvdd.n1237 604.457
R4245 dvdd.n1394 dvdd.n1393 604.457
R4246 dvdd.n1621 dvdd.n1506 604.457
R4247 dvdd.n1820 dvdd.n1819 604.457
R4248 dvdd.n577 dvdd.n534 604.394
R4249 dvdd.n933 dvdd.n932 604.394
R4250 dvdd.n1165 dvdd.n1110 604.394
R4251 dvdd.n1316 dvdd.n1228 604.394
R4252 dvdd.n1428 dvdd.n1408 604.394
R4253 dvdd.n1749 dvdd.n1690 604.394
R4254 dvdd.n1706 dvdd.n1705 604.394
R4255 dvdd.n1913 dvdd.n1912 604.394
R4256 dvdd.n2082 dvdd.n1795 604.394
R4257 dvdd.n1368 dvdd.n1338 604.076
R4258 dvdd.n2541 dvdd.n2519 603.38
R4259 dvdd.n492 dvdd.n478 603.231
R4260 dvdd.n986 dvdd.n947 603.015
R4261 dvdd.n1426 dvdd.n1409 603.015
R4262 dvdd.n1646 dvdd.n1645 603.015
R4263 dvdd.n2332 dvdd.n2119 603.015
R4264 dvdd.n818 dvdd.n817 601.907
R4265 dvdd.n1069 dvdd.n1066 601.732
R4266 dvdd.n729 dvdd.n634 601.679
R4267 dvdd.n1016 dvdd.n1015 601.679
R4268 dvdd.n1890 dvdd.n1889 601.679
R4269 dvdd.n1898 dvdd.n1897 601.679
R4270 dvdd.n1961 dvdd.n1943 601.679
R4271 dvdd.n471 dvdd.n470 601.097
R4272 dvdd.n749 dvdd.n746 601.097
R4273 dvdd.n824 dvdd.n823 601.097
R4274 dvdd.n1401 dvdd.n1400 601.097
R4275 dvdd.n1906 dvdd.n1905 601.097
R4276 dvdd.n1998 dvdd.n1994 601.004
R4277 dvdd.n1514 dvdd.n1513 600.322
R4278 dvdd.n453 dvdd.n356 600.105
R4279 dvdd.n336 dvdd.n335 600.105
R4280 dvdd.n639 dvdd.n638 600.105
R4281 dvdd.n999 dvdd.n942 600.105
R4282 dvdd.n1216 dvdd.n1215 600.105
R4283 dvdd.n1742 dvdd.n1693 600.105
R4284 dvdd.n1704 dvdd.n1703 600.105
R4285 dvdd.n1880 dvdd.n1822 600.105
R4286 dvdd.n1974 dvdd.n1935 600.105
R4287 dvdd.n1433 dvdd.n1405 599.966
R4288 dvdd.n2341 dvdd.n2115 599.966
R4289 dvdd.n1213 dvdd.n1212 599.933
R4290 dvdd.n1276 dvdd.n1251 599.74
R4291 dvdd.n1990 dvdd.n1989 599.203
R4292 dvdd.n677 dvdd.n676 598.986
R4293 dvdd.n1530 dvdd.n1528 598.986
R4294 dvdd.n1765 dvdd.n1498 598.986
R4295 dvdd.n1919 dvdd.n1810 598.986
R4296 dvdd.n1249 dvdd.n1248 598.965
R4297 dvdd.n1638 dvdd.n1637 598.572
R4298 dvdd.n351 dvdd.n350 598.383
R4299 dvdd.n527 dvdd.n526 598.383
R4300 dvdd.n938 dvdd.n937 598.383
R4301 dvdd.n1094 dvdd.n1054 598.383
R4302 dvdd.n1115 dvdd.n1114 598.383
R4303 dvdd.n1303 dvdd.n1233 598.383
R4304 dvdd.n1452 dvdd.n1392 598.383
R4305 dvdd.n1402 dvdd.n1399 598.383
R4306 dvdd.n1629 dvdd.n1628 598.383
R4307 dvdd.n1734 dvdd.n1696 598.383
R4308 dvdd.n1698 dvdd.n1697 598.383
R4309 dvdd.n2003 dvdd.n2002 598.383
R4310 dvdd.n2367 dvdd.n2365 596.97
R4311 dvdd.n687 dvdd.n649 596.619
R4312 dvdd.n978 dvdd.n977 596.619
R4313 dvdd.n1779 dvdd.n1493 596.619
R4314 dvdd.n1587 dvdd.n1585 596.619
R4315 dvdd.n770 dvdd.n767 596.442
R4316 dvdd.n1662 dvdd.n1661 595.303
R4317 dvdd.n2530 dvdd.n2526 594.144
R4318 dvdd.n2525 dvdd.n2524 594.144
R4319 dvdd.n2370 dvdd.n2369 594.144
R4320 dvdd.n2573 dvdd.n2572 594.144
R4321 dvdd.n2571 dvdd.n2569 594.144
R4322 dvdd.n2010 dvdd.n2009 592.04
R4323 dvdd.n1030 dvdd.n1029 591.601
R4324 dvdd.n1041 dvdd.n1040 591.601
R4325 dvdd dvdd.t1618 588.942
R4326 dvdd.n1518 dvdd.n1516 585
R4327 dvdd.n1517 dvdd.n1516 585
R4328 dvdd.n2517 dvdd.n2516 585
R4329 dvdd.n2521 dvdd.n2520 585
R4330 dvdd.n2615 dvdd.n2614 585
R4331 dvdd.t1780 dvdd 568.994
R4332 dvdd.t1531 dvdd.n193 544.548
R4333 dvdd.t1546 dvdd 515.284
R4334 dvdd.n2965 dvdd.n2961 510.118
R4335 dvdd.n2966 dvdd.n2965 510.118
R4336 dvdd.n2966 dvdd.n2946 510.118
R4337 dvdd.n2961 dvdd.n2946 510.118
R4338 dvdd dvdd.t1640 494.238
R4339 dvdd dvdd.t1583 493.464
R4340 dvdd.t1807 dvdd 458.724
R4341 dvdd.t1015 dvdd.t815 448.146
R4342 dvdd.n1030 dvdd.n1028 428.8
R4343 dvdd.n1041 dvdd.n930 428.8
R4344 dvdd.t797 dvdd 424.647
R4345 dvdd.n282 dvdd.t1474 417.291
R4346 dvdd dvdd.t1590 414.577
R4347 dvdd.t934 dvdd 412.899
R4348 dvdd.n670 dvdd.t1726 396.406
R4349 dvdd.n654 dvdd.t1725 391.005
R4350 dvdd.n2150 dvdd.t1699 390.875
R4351 dvdd.n1825 dvdd.t1548 390.062
R4352 dvdd.n2172 dvdd.t1717 389.195
R4353 dvdd.n506 dvdd.t1616 388.656
R4354 dvdd.n500 dvdd.t1617 388.656
R4355 dvdd.n651 dvdd.t1574 388.656
R4356 dvdd.n655 dvdd.t1573 388.656
R4357 dvdd.n964 dvdd.t1683 388.656
R4358 dvdd.n968 dvdd.t1684 388.656
R4359 dvdd.n1032 dvdd.t1635 388.656
R4360 dvdd.n1039 dvdd.t1636 388.656
R4361 dvdd.n1112 dvdd.t1659 388.656
R4362 dvdd.n1117 dvdd.t1660 388.656
R4363 dvdd.n1601 dvdd.t1731 388.656
R4364 dvdd.n1610 dvdd.t1732 388.656
R4365 dvdd.n1586 dvdd.t1545 388.656
R4366 dvdd.n1918 dvdd.t1632 388.656
R4367 dvdd.n1922 dvdd.t1633 388.656
R4368 dvdd.n1857 dvdd.t1547 388.656
R4369 dvdd.n1927 dvdd.t1604 388.656
R4370 dvdd.n1929 dvdd.t1605 388.656
R4371 dvdd.n2322 dvdd.t1664 388.656
R4372 dvdd.n2326 dvdd.t1665 388.656
R4373 dvdd.n2426 dvdd.t1766 388.656
R4374 dvdd.n2407 dvdd.t1767 388.656
R4375 dvdd.n2570 dvdd.t1691 388.656
R4376 dvdd.n2602 dvdd.t1692 388.656
R4377 dvdd.n209 dvdd.t1808 388.656
R4378 dvdd.n212 dvdd.t1809 388.656
R4379 dvdd.n135 dvdd.t1625 388.656
R4380 dvdd.n92 dvdd.t1624 388.656
R4381 dvdd.n694 dvdd.t1728 388.656
R4382 dvdd.n700 dvdd.t1729 388.656
R4383 dvdd.n768 dvdd.t1751 388.656
R4384 dvdd.n778 dvdd.t1752 388.656
R4385 dvdd.n892 dvdd.t1576 388.656
R4386 dvdd.n624 dvdd.t1577 388.656
R4387 dvdd.n2076 dvdd.t1644 388.656
R4388 dvdd.n2070 dvdd.t1645 388.656
R4389 dvdd.n2576 dvdd.t1529 388.656
R4390 dvdd.n2590 dvdd.t1530 388.656
R4391 dvdd.n2163 dvdd.t1586 385.026
R4392 dvdd.n2391 dvdd.t1798 382.673
R4393 dvdd.n230 dvdd.t1641 381.443
R4394 dvdd.n294 dvdd.t1714 381.443
R4395 dvdd.n83 dvdd.t1715 381.443
R4396 dvdd.n90 dvdd.t1532 381.443
R4397 dvdd.n151 dvdd.t1533 381.443
R4398 dvdd.n164 dvdd.t1619 381.443
R4399 dvdd.n165 dvdd.t1620 381.443
R4400 dvdd.n2335 dvdd.t1621 381.443
R4401 dvdd.n2116 dvdd.t1622 381.443
R4402 dvdd.n233 dvdd.t1642 381.443
R4403 dvdd.n377 dvdd.t1647 380.193
R4404 dvdd.n380 dvdd.t1748 380.193
R4405 dvdd.n535 dvdd.t1696 380.193
R4406 dvdd.n547 dvdd.t1667 380.193
R4407 dvdd.n550 dvdd.t1759 380.193
R4408 dvdd.n656 dvdd.t1541 380.193
R4409 dvdd.n660 dvdd.t1685 380.193
R4410 dvdd.n825 dvdd.t1607 380.193
R4411 dvdd.n836 dvdd.t1562 380.193
R4412 dvdd.n839 dvdd.t1703 380.193
R4413 dvdd.n954 dvdd.t1743 380.193
R4414 dvdd.n957 dvdd.t1579 380.193
R4415 dvdd.n1123 dvdd.t1755 380.193
R4416 dvdd.n1126 dvdd.t1610 380.193
R4417 dvdd.n1257 dvdd.t1588 380.193
R4418 dvdd.n1260 dvdd.t1584 380.193
R4419 dvdd.n1414 dvdd.t1626 380.193
R4420 dvdd.n1417 dvdd.t1613 380.193
R4421 dvdd.n1544 dvdd.t1601 380.193
R4422 dvdd.n1548 dvdd.t1787 380.193
R4423 dvdd.n1707 dvdd.t1629 380.193
R4424 dvdd.n1710 dvdd.t1805 380.193
R4425 dvdd.n1833 dvdd.t1794 380.193
R4426 dvdd.n1836 dvdd.t1722 380.193
R4427 dvdd.n1995 dvdd.t1653 380.193
R4428 dvdd.n2018 dvdd.t1535 380.193
R4429 dvdd.n2021 dvdd.t1738 380.193
R4430 dvdd.n2140 dvdd.t1705 380.193
R4431 dvdd.n2236 dvdd.t1557 380.193
R4432 dvdd.n2239 dvdd.t1757 380.193
R4433 dvdd.n2107 dvdd.t1523 380.193
R4434 dvdd.n2188 dvdd.t1581 380.193
R4435 dvdd.n2191 dvdd.t1778 380.193
R4436 dvdd.n2474 dvdd.t1554 380.193
R4437 dvdd.n2511 dvdd.t1774 380.193
R4438 dvdd.n2380 dvdd.t1526 380.193
R4439 dvdd.n2458 dvdd.t1656 380.193
R4440 dvdd.n2412 dvdd.t1771 380.193
R4441 dvdd.n2415 dvdd.t1701 380.193
R4442 dvdd.n2581 dvdd.t1783 380.193
R4443 dvdd.n2584 dvdd.t1711 380.193
R4444 dvdd.t556 dvdd.n2963 369.05
R4445 dvdd.n2964 dvdd.t560 369.05
R4446 dvdd.t1543 dvdd.t1099 364.224
R4447 dvdd.n3128 dvdd.t1284 360.925
R4448 dvdd.t1724 dvdd 360.866
R4449 dvdd.n3126 dvdd.t1292 360.795
R4450 dvdd.n1754 dvdd.t986 353.774
R4451 dvdd.n354 dvdd.t943 353.774
R4452 dvdd.n1083 dvdd.t941 353.774
R4453 dvdd.n1081 dvdd.t939 353.774
R4454 dvdd.n1273 dvdd.t1298 353.774
R4455 dvdd.n438 dvdd.t461 350.582
R4456 dvdd dvdd.t186 350
R4457 dvdd dvdd.t691 350
R4458 dvdd.n2821 dvdd.t291 349.238
R4459 dvdd.n2887 dvdd.t215 348.805
R4460 dvdd.n3041 dvdd.t978 348.755
R4461 dvdd.n2984 dvdd.t39 348.755
R4462 dvdd.n446 dvdd.t469 347.572
R4463 dvdd.n1061 dvdd.t327 343.579
R4464 dvdd.n1616 dvdd.t1226 343.579
R4465 dvdd.n1824 dvdd.t257 343.579
R4466 dvdd.n619 dvdd.t1072 343.577
R4467 dvdd.n991 dvdd.t716 343.577
R4468 dvdd.n1289 dvdd.t1052 343.577
R4469 dvdd.n1209 dvdd.t641 343.577
R4470 dvdd.n1706 dvdd.t1342 343.308
R4471 dvdd.n1749 dvdd.t397 343.308
R4472 dvdd.n1766 dvdd.t83 342.841
R4473 dvdd.t1643 dvdd.t148 342.404
R4474 dvdd dvdd.t687 341.488
R4475 dvdd dvdd.t993 341.488
R4476 dvdd.n1652 dvdd.t1401 340.301
R4477 dvdd.n1340 dvdd.t1046 340.243
R4478 dvdd.n1479 dvdd.t776 340.211
R4479 dvdd.n992 dvdd.t233 340.012
R4480 dvdd.n1133 dvdd.t1345 340.012
R4481 dvdd.n1391 dvdd.t1040 340.012
R4482 dvdd.n1930 dvdd.t450 340.012
R4483 dvdd.n484 dvdd.t1266 340.01
R4484 dvdd.n708 dvdd.t881 340.01
R4485 dvdd.n1823 dvdd.t1203 340.01
R4486 dvdd.n1806 dvdd.t316 340.01
R4487 dvdd.n2333 dvdd.t739 337.952
R4488 dvdd.n1630 dvdd.t75 337.372
R4489 dvdd dvdd.t1578 337.368
R4490 dvdd dvdd.t711 336.933
R4491 dvdd.n530 dvdd.t513 336.567
R4492 dvdd.n1111 dvdd.t459 336.567
R4493 dvdd.n794 dvdd.t1455 336.524
R4494 dvdd.n1931 dvdd.t1463 336.522
R4495 dvdd.n904 dvdd.t1162 336.416
R4496 dvdd.n1173 dvdd.t930 336.416
R4497 dvdd.n1282 dvdd.t1388 334.784
R4498 dvdd.n575 dvdd.t269 334.634
R4499 dvdd.n1626 dvdd.t749 334.497
R4500 dvdd dvdd.t1646 334.012
R4501 dvdd dvdd.t1540 334.012
R4502 dvdd dvdd.t1600 334.012
R4503 dvdd dvdd.t1721 334.012
R4504 dvdd dvdd.t1700 334.012
R4505 dvdd.n1576 dvdd.t866 333.8
R4506 dvdd.n1595 dvdd.t1246 333.798
R4507 dvdd.n925 dvdd.t1333 333.368
R4508 dvdd.n1562 dvdd.t101 333.368
R4509 dvdd.t356 dvdd.t991 330.654
R4510 dvdd.t795 dvdd.t340 330.654
R4511 dvdd.t819 dvdd.t336 330.654
R4512 dvdd.n2297 dvdd.t1876 328.005
R4513 dvdd.t468 dvdd.t1507 327.298
R4514 dvdd.n2351 dvdd.n2105 325.639
R4515 dvdd.n2157 dvdd.n2152 324.74
R4516 dvdd.n619 dvdd.n618 324.543
R4517 dvdd.n360 dvdd.n359 323.988
R4518 dvdd dvdd.t1531 322.587
R4519 dvdd.t1713 dvdd 322.587
R4520 dvdd.t1640 dvdd 322.587
R4521 dvdd.n1179 dvdd.n927 322.329
R4522 dvdd.n1534 dvdd.n1533 322.329
R4523 dvdd.n480 dvdd.n479 320.976
R4524 dvdd.n1105 dvdd.n1104 320.976
R4525 dvdd.n2925 dvdd.n2874 320.976
R4526 dvdd.n2914 dvdd.n2878 320.976
R4527 dvdd.n2880 dvdd.n2879 320.976
R4528 dvdd.n2906 dvdd.n2882 320.976
R4529 dvdd.n2900 dvdd.n2899 320.976
R4530 dvdd.n2897 dvdd.n2885 320.976
R4531 dvdd.n2891 dvdd.n2890 320.976
R4532 dvdd.n2889 dvdd.n2888 320.976
R4533 dvdd.n3079 dvdd.n3028 320.976
R4534 dvdd.n3068 dvdd.n3032 320.976
R4535 dvdd.n3034 dvdd.n3033 320.976
R4536 dvdd.n3060 dvdd.n3036 320.976
R4537 dvdd.n3054 dvdd.n3053 320.976
R4538 dvdd.n3051 dvdd.n3039 320.976
R4539 dvdd.n3045 dvdd.n3044 320.976
R4540 dvdd.n3043 dvdd.n3042 320.976
R4541 dvdd.n3022 dvdd.n2971 320.976
R4542 dvdd.n3011 dvdd.n2975 320.976
R4543 dvdd.n2977 dvdd.n2976 320.976
R4544 dvdd.n3003 dvdd.n2979 320.976
R4545 dvdd.n2997 dvdd.n2996 320.976
R4546 dvdd.n2994 dvdd.n2982 320.976
R4547 dvdd.n2988 dvdd.n2987 320.976
R4548 dvdd.n2986 dvdd.n2985 320.976
R4549 dvdd.n2858 dvdd.n2808 320.976
R4550 dvdd.n2868 dvdd.n2804 320.976
R4551 dvdd.n2848 dvdd.n2812 320.976
R4552 dvdd.n2814 dvdd.n2813 320.976
R4553 dvdd.n2840 dvdd.n2816 320.976
R4554 dvdd.n2834 dvdd.n2833 320.976
R4555 dvdd.n2831 dvdd.n2819 320.976
R4556 dvdd.n2825 dvdd.n2824 320.976
R4557 dvdd.n2823 dvdd.n2822 320.976
R4558 dvdd.n1647 dvdd.n1642 320.976
R4559 dvdd.n2014 dvdd.n2013 317.943
R4560 dvdd.t252 dvdd.t1054 317.226
R4561 dvdd.n2031 dvdd.n2016 317.103
R4562 dvdd.n1759 dvdd.n1685 316.974
R4563 dvdd.n1616 dvdd.n1509 316.693
R4564 dvdd.n282 dvdd 316.668
R4565 dvdd.n281 dvdd 316.668
R4566 dvdd.n758 dvdd.n757 315.334
R4567 dvdd.n1350 dvdd.n1349 315.334
R4568 dvdd.n1937 dvdd.n1936 315.334
R4569 dvdd.n803 dvdd.n802 315.089
R4570 dvdd.n787 dvdd.n763 313.591
R4571 dvdd.n2274 dvdd.t1824 312.89
R4572 dvdd.n1320 dvdd.n1225 312.829
R4573 dvdd.n1047 dvdd.n1046 312.827
R4574 dvdd.t1413 dvdd.t458 312.192
R4575 dvdd.n107 dvdd.n106 312.053
R4576 dvdd.n1425 dvdd.n1412 312.053
R4577 dvdd.n2012 dvdd.n2011 312.053
R4578 dvdd.n2186 dvdd.n2185 312.053
R4579 dvdd.n2186 dvdd.n2184 312.051
R4580 dvdd.n2565 dvdd.n2564 312.051
R4581 dvdd.n969 dvdd.n967 312.005
R4582 dvdd.n1849 dvdd.n1831 312.005
R4583 dvdd.n1370 dvdd.n1334 311.659
R4584 dvdd.n2367 dvdd.n2366 311.582
R4585 dvdd.n1976 dvdd.n1934 311.149
R4586 dvdd.n1347 dvdd.n1346 310.902
R4587 dvdd.n498 dvdd.n474 310.502
R4588 dvdd.n493 dvdd.n477 310.502
R4589 dvdd.n2473 dvdd.t1879 309.962
R4590 dvdd.n532 dvdd.n531 309.726
R4591 dvdd.n923 dvdd.n922 309.726
R4592 dvdd.n1166 dvdd.n1107 309.724
R4593 dvdd.n2557 dvdd.n2385 309.7
R4594 dvdd.n2316 dvdd.n2126 309.531
R4595 dvdd.t1649 dvdd.t1780 308.834
R4596 dvdd.t1687 dvdd.t1727 308.834
R4597 dvdd.t1305 dvdd 308.834
R4598 dvdd.n2324 dvdd.n2123 308.755
R4599 dvdd.n2493 dvdd.n2492 308.755
R4600 dvdd.n2482 dvdd.n2397 308.755
R4601 dvdd.n2466 dvdd.n2465 308.755
R4602 dvdd.n2454 dvdd.n2403 308.755
R4603 dvdd.n1134 dvdd.n1122 308.755
R4604 dvdd.n1539 dvdd.n1538 308.755
R4605 dvdd.n1554 dvdd.n1542 308.755
R4606 dvdd.n2182 dvdd.n2181 308.755
R4607 dvdd.n2591 dvdd.n2580 308.755
R4608 dvdd.n3092 dvdd.n3084 307.762
R4609 dvdd.n2800 dvdd.n3 307.762
R4610 dvdd.n2796 dvdd.n10 307.762
R4611 dvdd.n2792 dvdd.n17 307.762
R4612 dvdd.n2788 dvdd.n24 307.762
R4613 dvdd.n2784 dvdd.n31 307.762
R4614 dvdd.n2780 dvdd.n38 307.762
R4615 dvdd.n2776 dvdd.n45 307.762
R4616 dvdd.n2772 dvdd.n52 307.762
R4617 dvdd.n2768 dvdd.n59 307.762
R4618 dvdd.n2718 dvdd.n2716 307.762
R4619 dvdd.n2722 dvdd.n2709 307.762
R4620 dvdd.n2726 dvdd.n2702 307.762
R4621 dvdd.n2730 dvdd.n2695 307.762
R4622 dvdd.n2734 dvdd.n2688 307.762
R4623 dvdd.n2738 dvdd.n2681 307.762
R4624 dvdd.n2742 dvdd.n2674 307.762
R4625 dvdd.n2746 dvdd.n2667 307.762
R4626 dvdd.n2750 dvdd.n2660 307.762
R4627 dvdd.n1281 dvdd.n1247 307.204
R4628 dvdd.n1778 dvdd.n1494 307.204
R4629 dvdd.n785 dvdd.n764 307.204
R4630 dvdd.n225 dvdd.t1848 306.735
R4631 dvdd.n219 dvdd.t1810 306.735
R4632 dvdd.n307 dvdd.t1884 306.735
R4633 dvdd.n101 dvdd.t1857 306.735
R4634 dvdd.n160 dvdd.t1866 306.735
R4635 dvdd.n374 dvdd.t1839 306.735
R4636 dvdd.n374 dvdd.t1892 306.735
R4637 dvdd.n417 dvdd.t1822 306.735
R4638 dvdd.n423 dvdd.t1880 306.735
R4639 dvdd.n440 dvdd.t1875 306.735
R4640 dvdd.n542 dvdd.t1814 306.735
R4641 dvdd.n542 dvdd.t1871 306.735
R4642 dvdd.n709 dvdd.t1817 306.735
R4643 dvdd.n688 dvdd.t1836 306.735
R4644 dvdd.n821 dvdd.t1885 306.735
R4645 dvdd.n831 dvdd.t1816 306.735
R4646 dvdd.n831 dvdd.t1846 306.735
R4647 dvdd.n1234 dvdd.t1907 306.735
R4648 dvdd.n1851 dvdd.t1827 306.735
R4649 dvdd.n2004 dvdd.t1863 306.735
R4650 dvdd.n2233 dvdd.t1852 306.735
R4651 dvdd.n2233 dvdd.t1893 306.735
R4652 dvdd.n2130 dvdd.t1813 306.735
R4653 dvdd.n2137 dvdd.t1882 306.735
R4654 dvdd.n2219 dvdd.t1889 306.735
R4655 dvdd.n2178 dvdd.t1890 306.735
R4656 dvdd.n2429 dvdd.t1819 306.735
R4657 dvdd.n2447 dvdd.t1853 306.735
R4658 dvdd.n1623 dvdd.n1504 306.541
R4659 dvdd.n588 dvdd.n529 306.428
R4660 dvdd.n1556 dvdd.n1555 306.428
R4661 dvdd.t880 dvdd.t1799 305.478
R4662 dvdd.n1657 dvdd.n1656 292.5
R4663 dvdd.n1659 dvdd.n1658 292.5
R4664 dvdd.t1442 dvdd.t1690 288.693
R4665 dvdd.n2145 dvdd.t70 284.029
R4666 dvdd.t323 dvdd.t1718 283.658
R4667 dvdd.t1472 dvdd.t1428 281.154
R4668 dvdd dvdd.t460 280.3
R4669 dvdd dvdd.t1666 280.3
R4670 dvdd dvdd.t1606 280.3
R4671 dvdd dvdd.t1561 280.3
R4672 dvdd dvdd.t1609 280.3
R4673 dvdd dvdd.t1628 280.3
R4674 dvdd dvdd.t1655 280.3
R4675 dvdd dvdd.t1553 280.3
R4676 dvdd dvdd.t1796 280.3
R4677 dvdd dvdd.t1710 280.3
R4678 dvdd.n2229 dvdd.n2228 278.93
R4679 dvdd.n2228 dvdd.n2227 278.858
R4680 dvdd dvdd.t1612 278.623
R4681 dvdd dvdd.t1534 278.623
R4682 dvdd.t1387 dvdd.t1370 276.943
R4683 dvdd.n1520 dvdd.n1519 275.348
R4684 dvdd.n1355 dvdd.n1345 274.346
R4685 dvdd.n2146 dvdd.n2145 269.485
R4686 dvdd.n2227 dvdd.n2147 269.485
R4687 dvdd.n2229 dvdd.n2147 269.483
R4688 dvdd.n646 dvdd.t853 266.873
R4689 dvdd.t554 dvdd.t556 264.262
R4690 dvdd.t552 dvdd.t554 264.262
R4691 dvdd.t1290 dvdd.t552 264.262
R4692 dvdd.t713 dvdd.t1290 264.262
R4693 dvdd.t703 dvdd.t713 264.262
R4694 dvdd.t701 dvdd.t703 264.262
R4695 dvdd.t568 dvdd.t701 264.262
R4696 dvdd.t566 dvdd.t568 264.262
R4697 dvdd.t562 dvdd.t566 264.262
R4698 dvdd.t558 dvdd.t562 264.262
R4699 dvdd.t564 dvdd.t558 264.262
R4700 dvdd.t560 dvdd.t564 264.262
R4701 dvdd.t538 dvdd.t760 263.397
R4702 dvdd.t1128 dvdd.t401 261.837
R4703 dvdd.t1727 dvdd 260.159
R4704 dvdd.t985 dvdd 260.159
R4705 dvdd dvdd.t1546 260.159
R4706 dvdd.t1631 dvdd 260.159
R4707 dvdd.n1499 dvdd.t91 257.474
R4708 dvdd dvdd.t315 256.803
R4709 dvdd.n472 dvdd.t1168 255.976
R4710 dvdd.n2600 dvdd.t1125 255.904
R4711 dvdd.t1158 dvdd.t538 254.518
R4712 dvdd.n2876 dvdd.t213 250.785
R4713 dvdd.n3030 dvdd.t976 250.785
R4714 dvdd.n2973 dvdd.t37 250.785
R4715 dvdd.n2810 dvdd.t277 250.785
R4716 dvdd.n1608 dvdd.t139 250.724
R4717 dvdd.n487 dvdd.t1279 249.901
R4718 dvdd.n1687 dvdd.t1228 249.901
R4719 dvdd.n197 dvdd.t25 249.363
R4720 dvdd.n87 dvdd.t1475 249.363
R4721 dvdd.n771 dvdd.t770 249.363
R4722 dvdd.n1167 dvdd.t1492 249.363
R4723 dvdd.n1413 dvdd.t722 249.363
R4724 dvdd.n2196 dvdd.t1518 249.363
R4725 dvdd.n2490 dvdd.t1410 249.363
R4726 dvdd.n2639 dvdd.t1133 249.363
R4727 dvdd.n987 dvdd.t856 249.362
R4728 dvdd.n984 dvdd.t503 249.362
R4729 dvdd.n1172 dvdd.t607 249.362
R4730 dvdd.n1567 dvdd.t456 249.362
R4731 dvdd.n1552 dvdd.t1004 249.362
R4732 dvdd.n1644 dvdd.t392 249.362
R4733 dvdd.n1869 dvdd.t812 249.362
R4734 dvdd.n2196 dvdd.t1398 249.362
R4735 dvdd.n2613 dvdd.t3 249.362
R4736 dvdd.n2124 dvdd.t1220 248.929
R4737 dvdd.t1474 dvdd.t1472 248.599
R4738 dvdd.t1430 dvdd.t24 248.599
R4739 dvdd.t1515 dvdd 248.411
R4740 dvdd.n1609 dvdd.t145 248.219
R4741 dvdd.n2577 dvdd.t1127 248.219
R4742 dvdd.n2393 dvdd.t1894 247.744
R4743 dvdd.n2464 dvdd.t1218 247.542
R4744 dvdd.n322 dvdd.t1431 247.394
R4745 dvdd.n985 dvdd.t1296 247.394
R4746 dvdd.n950 dvdd.t1110 247.394
R4747 dvdd.n1168 dvdd.t1488 247.394
R4748 dvdd.t1142 dvdd.t1132 246.732
R4749 dvdd.n707 dvdd.t879 246.111
R4750 dvdd.n71 dvdd.t1059 246.106
R4751 dvdd.n2652 dvdd.t625 246.106
R4752 dvdd.n378 dvdd.t1821 245.667
R4753 dvdd.n381 dvdd.t1868 245.667
R4754 dvdd.n536 dvdd.t1841 245.667
R4755 dvdd.n548 dvdd.t1831 245.667
R4756 dvdd.n551 dvdd.t1873 245.667
R4757 dvdd.n657 dvdd.t1895 245.667
R4758 dvdd.n661 dvdd.t1870 245.667
R4759 dvdd.n826 dvdd.t1908 245.667
R4760 dvdd.n837 dvdd.t1903 245.667
R4761 dvdd.n840 dvdd.t1874 245.667
R4762 dvdd.n955 dvdd.t1865 245.667
R4763 dvdd.n958 dvdd.t1845 245.667
R4764 dvdd.n1124 dvdd.t1872 245.667
R4765 dvdd.n1127 dvdd.t1851 245.667
R4766 dvdd.n1258 dvdd.t1838 245.667
R4767 dvdd.n1261 dvdd.t1811 245.667
R4768 dvdd.n1415 dvdd.t1847 245.667
R4769 dvdd.n1418 dvdd.t1818 245.667
R4770 dvdd.n1545 dvdd.t1842 245.667
R4771 dvdd.n1549 dvdd.t1883 245.667
R4772 dvdd.n1708 dvdd.t1849 245.667
R4773 dvdd.n1711 dvdd.t1891 245.667
R4774 dvdd.n1834 dvdd.t1909 245.667
R4775 dvdd.n1837 dvdd.t1859 245.667
R4776 dvdd.n1996 dvdd.t1834 245.667
R4777 dvdd.n2019 dvdd.t1815 245.667
R4778 dvdd.n2022 dvdd.t1864 245.667
R4779 dvdd.n2141 dvdd.t1858 245.667
R4780 dvdd.n2237 dvdd.t1823 245.667
R4781 dvdd.n2240 dvdd.t1877 245.667
R4782 dvdd.n2108 dvdd.t1900 245.667
R4783 dvdd.n2189 dvdd.t1832 245.667
R4784 dvdd.n2192 dvdd.t1887 245.667
R4785 dvdd.n2475 dvdd.t1911 245.667
R4786 dvdd.n2512 dvdd.t1881 245.667
R4787 dvdd.n2381 dvdd.t1910 245.667
R4788 dvdd.n2459 dvdd.t1837 245.667
R4789 dvdd.n2413 dvdd.t1897 245.667
R4790 dvdd.n2416 dvdd.t1855 245.667
R4791 dvdd.n2582 dvdd.t1904 245.667
R4792 dvdd.n2585 dvdd.t1860 245.667
R4793 dvdd.n2399 dvdd.t657 245.178
R4794 dvdd.n2379 dvdd.t852 245.178
R4795 dvdd.n2446 dvdd.t1314 245.178
R4796 dvdd.n1052 dvdd.t73 245.178
R4797 dvdd.t376 dvdd.t727 245.054
R4798 dvdd.n2927 dvdd.t710 244.737
R4799 dvdd.n3081 dvdd.t686 244.737
R4800 dvdd.n3024 dvdd.t996 244.737
R4801 dvdd.n2870 dvdd.t690 244.737
R4802 dvdd.n2806 dvdd.t193 244.737
R4803 dvdd.n1759 dvdd.t79 244.192
R4804 dvdd.n1075 dvdd.t310 244.191
R4805 dvdd.n1268 dvdd.t1506 244.191
R4806 dvdd.n1315 dvdd.t753 243.512
R4807 dvdd.n1055 dvdd.t611 243.508
R4808 dvdd.n1874 dvdd.t81 243.508
R4809 dvdd.n1600 dvdd.t1055 243.127
R4810 dvdd.n232 dvdd.t1905 242.282
R4811 dvdd.n295 dvdd.t1830 242.282
R4812 dvdd.n91 dvdd.t1869 242.282
R4813 dvdd.n166 dvdd.t1898 242.282
R4814 dvdd.n2336 dvdd.t1828 242.282
R4815 dvdd.n3121 dvdd.t1287 241.409
R4816 dvdd.n462 dvdd.t1014 240.792
R4817 dvdd.n1088 dvdd.t659 240.792
R4818 dvdd.n3134 dvdd.t1282 240.538
R4819 dvdd.n2945 dvdd.t1289 240.488
R4820 dvdd.n976 dvdd.t85 240.214
R4821 dvdd.t666 dvdd 238.339
R4822 dvdd dvdd.t498 236.661
R4823 dvdd.n2448 dvdd.t1313 236.661
R4824 dvdd.n808 dvdd.n753 235.248
R4825 dvdd.t440 dvdd.t1323 234.982
R4826 dvdd.t1021 dvdd.t1033 234.982
R4827 dvdd.t1416 dvdd.t1280 234.982
R4828 dvdd.t1134 dvdd.t432 234.982
R4829 dvdd.t1299 dvdd 234.982
R4830 dvdd.t785 dvdd.t16 234.982
R4831 dvdd.t632 dvdd.n2555 234.982
R4832 dvdd.t1039 dvdd.t330 229.947
R4833 dvdd.n2944 dvdd.t561 228.669
R4834 dvdd.t622 dvdd.t502 226.59
R4835 dvdd.t1358 dvdd.n3142 224.668
R4836 dvdd.n920 dvdd.n919 223.869
R4837 dvdd.n488 dvdd.n482 223.868
R4838 dvdd.t1362 dvdd.t1360 223.429
R4839 dvdd.t1352 dvdd.t1362 223.429
R4840 dvdd.t1618 dvdd 221.964
R4841 dvdd.n193 dvdd 221.964
R4842 dvdd dvdd.n281 221.964
R4843 dvdd.t1379 dvdd.t1191 221.555
R4844 dvdd.t1183 dvdd.t1733 221.555
R4845 dvdd.t286 dvdd.t290 221.054
R4846 dvdd.t280 dvdd.t286 221.054
R4847 dvdd.t292 dvdd.t280 221.054
R4848 dvdd.t282 dvdd.t292 221.054
R4849 dvdd.t294 dvdd.t282 221.054
R4850 dvdd.t272 dvdd.t294 221.054
R4851 dvdd.t284 dvdd.t272 221.054
R4852 dvdd.t296 dvdd.t284 221.054
R4853 dvdd.t288 dvdd.t296 221.054
R4854 dvdd.t300 dvdd.t288 221.054
R4855 dvdd.t278 dvdd.t300 221.054
R4856 dvdd.t274 dvdd.t278 221.054
R4857 dvdd.t302 dvdd.t298 221.054
R4858 dvdd.t298 dvdd.t276 221.054
R4859 dvdd.t186 dvdd.t190 221.054
R4860 dvdd.t190 dvdd.t188 221.054
R4861 dvdd.t188 dvdd.t192 221.054
R4862 dvdd.t691 dvdd.t699 221.054
R4863 dvdd.t699 dvdd.t683 221.054
R4864 dvdd.t683 dvdd.t689 221.054
R4865 dvdd dvdd.t878 219.876
R4866 dvdd.t1185 dvdd.t586 219.876
R4867 dvdd.t1400 dvdd 219.876
R4868 dvdd.t12 dvdd.t1097 219.876
R4869 dvdd.t1085 dvdd.t21 219.876
R4870 dvdd.n1465 dvdd.n1214 219.517
R4871 dvdd.t853 dvdd.t934 218.198
R4872 dvdd.t270 dvdd.t134 218.198
R4873 dvdd.t1187 dvdd.t1185 218.198
R4874 dvdd dvdd.t584 216.519
R4875 dvdd.t951 dvdd.t977 215.677
R4876 dvdd.t947 dvdd.t951 215.677
R4877 dvdd.t959 dvdd.t947 215.677
R4878 dvdd.t953 dvdd.t959 215.677
R4879 dvdd.t949 dvdd.t953 215.677
R4880 dvdd.t961 dvdd.t949 215.677
R4881 dvdd.t955 dvdd.t961 215.677
R4882 dvdd.t969 dvdd.t955 215.677
R4883 dvdd.t965 dvdd.t969 215.677
R4884 dvdd.t971 dvdd.t965 215.677
R4885 dvdd.t963 dvdd.t957 215.677
R4886 dvdd.t957 dvdd.t973 215.677
R4887 dvdd.t973 dvdd.t967 215.677
R4888 dvdd.t967 dvdd.t975 215.677
R4889 dvdd.t687 dvdd.t695 215.677
R4890 dvdd.t695 dvdd.t697 215.677
R4891 dvdd.t697 dvdd.t685 215.677
R4892 dvdd.t44 dvdd.t38 215.677
R4893 dvdd.t40 dvdd.t44 215.677
R4894 dvdd.t52 dvdd.t40 215.677
R4895 dvdd.t46 dvdd.t52 215.677
R4896 dvdd.t42 dvdd.t46 215.677
R4897 dvdd.t54 dvdd.t42 215.677
R4898 dvdd.t48 dvdd.t54 215.677
R4899 dvdd.t62 dvdd.t48 215.677
R4900 dvdd.t58 dvdd.t62 215.677
R4901 dvdd.t64 dvdd.t58 215.677
R4902 dvdd.t56 dvdd.t50 215.677
R4903 dvdd.t50 dvdd.t66 215.677
R4904 dvdd.t66 dvdd.t60 215.677
R4905 dvdd.t60 dvdd.t36 215.677
R4906 dvdd.t993 dvdd.t999 215.677
R4907 dvdd.t999 dvdd.t997 215.677
R4908 dvdd.t997 dvdd.t995 215.677
R4909 dvdd.t540 dvdd 213.163
R4910 dvdd dvdd.t433 213.163
R4911 dvdd dvdd.t1063 213.163
R4912 dvdd.n1100 dvdd.n1099 213.119
R4913 dvdd.n1386 dvdd.n1385 213.119
R4914 dvdd.n1992 dvdd.n1991 213.119
R4915 dvdd.n281 dvdd.n280 213.119
R4916 dvdd.n283 dvdd.n282 213.119
R4917 dvdd.n193 dvdd.n192 213.119
R4918 dvdd.n945 dvdd.n944 213.119
R4919 dvdd.n1245 dvdd.n1244 213.119
R4920 dvdd.n1460 dvdd.n1387 213.119
R4921 dvdd.n1760 dvdd.n1684 213.119
R4922 dvdd.t220 dvdd.t214 212.8
R4923 dvdd.t216 dvdd.t220 212.8
R4924 dvdd.t196 dvdd.t216 212.8
R4925 dvdd.t222 dvdd.t196 212.8
R4926 dvdd.t218 dvdd.t222 212.8
R4927 dvdd.t198 dvdd.t218 212.8
R4928 dvdd.t224 dvdd.t198 212.8
R4929 dvdd.t206 dvdd.t224 212.8
R4930 dvdd.t202 dvdd.t206 212.8
R4931 dvdd.t208 dvdd.t202 212.8
R4932 dvdd.t200 dvdd.t194 212.8
R4933 dvdd.t194 dvdd.t210 212.8
R4934 dvdd.t210 dvdd.t204 212.8
R4935 dvdd.t204 dvdd.t212 212.8
R4936 dvdd.t711 dvdd.t705 212.8
R4937 dvdd.t705 dvdd.t707 212.8
R4938 dvdd.t707 dvdd.t709 212.8
R4939 dvdd.n1868 dvdd.n1826 211.732
R4940 dvdd dvdd.t912 211.484
R4941 dvdd.n210 dvdd.t1867 210.964
R4942 dvdd.n505 dvdd.t1812 210.964
R4943 dvdd.n645 dvdd.t1888 210.964
R4944 dvdd.n654 dvdd.t1886 210.964
R4945 dvdd.n769 dvdd.t1901 210.964
R4946 dvdd.n891 dvdd.t1844 210.964
R4947 dvdd.n965 dvdd.t1840 210.964
R4948 dvdd.n1031 dvdd.t1820 210.964
R4949 dvdd.n1920 dvdd.t1850 210.964
R4950 dvdd.n1928 dvdd.t1843 210.964
R4951 dvdd.n2075 dvdd.t1829 210.964
R4952 dvdd.n2323 dvdd.t1856 210.964
R4953 dvdd dvdd.t232 209.806
R4954 dvdd dvdd.t1479 209.806
R4955 dvdd.n2557 dvdd.n2556 209.486
R4956 dvdd.n593 dvdd.n525 209.368
R4957 dvdd.n524 dvdd.n523 209.368
R4958 dvdd.n884 dvdd.n814 209.368
R4959 dvdd.n813 dvdd.n812 209.368
R4960 dvdd.n693 dvdd.n646 209.368
R4961 dvdd.n1177 dvdd.n1101 209.368
R4962 dvdd.n1530 dvdd.n1529 209.368
R4963 dvdd.n1683 dvdd.n1682 209.368
R4964 dvdd.n2067 dvdd.n1993 209.368
R4965 dvdd.n2449 dvdd.n2448 209.368
R4966 dvdd.t1265 dvdd 208.127
R4967 dvdd dvdd.t1225 206.45
R4968 dvdd dvdd.t256 206.45
R4969 dvdd.n2764 dvdd.n66 205.5
R4970 dvdd.n2754 dvdd.n2653 205.5
R4971 dvdd.t276 dvdd 205.263
R4972 dvdd.t1099 dvdd 204.77
R4973 dvdd.t1615 dvdd 203.093
R4974 dvdd.n144 dvdd.n94 202.66
R4975 dvdd.n3123 dvdd.n3117 200.31
R4976 dvdd.n3132 dvdd.n3129 200.31
R4977 dvdd.n3131 dvdd.n3130 200.31
R4978 dvdd.n3122 dvdd.n3118 200.31
R4979 dvdd.n3120 dvdd.n3119 200.31
R4980 dvdd.n3098 dvdd.n3097 200.31
R4981 dvdd.t975 dvdd 200.27
R4982 dvdd.t36 dvdd 200.27
R4983 dvdd.n3153 dvdd.n3152 200.173
R4984 dvdd.n3126 dvdd.n3125 200.115
R4985 dvdd.n2957 dvdd.n2956 200.105
R4986 dvdd.n2958 dvdd.n2955 200.105
R4987 dvdd.n2959 dvdd.n2954 200.105
R4988 dvdd.n2953 dvdd.n2948 200.105
R4989 dvdd.n2952 dvdd.n2949 200.105
R4990 dvdd.n2951 dvdd.n2950 200.105
R4991 dvdd.n3126 dvdd.n3124 200.095
R4992 dvdd.n3128 dvdd.n3127 200.034
R4993 dvdd.t612 dvdd.t1115 199.736
R4994 dvdd.t1243 dvdd.t793 199.736
R4995 dvdd.t262 dvdd.t925 199.736
R4996 dvdd.t1229 dvdd.t1375 199.736
R4997 dvdd.t746 dvdd 199.736
R4998 dvdd.t212 dvdd 197.601
R4999 dvdd.t192 dvdd 197.369
R5000 dvdd.t689 dvdd 197.369
R5001 dvdd dvdd.t268 196.379
R5002 dvdd.t68 dvdd.n1992 196.379
R5003 dvdd.t1350 dvdd.t927 194.701
R5004 dvdd.t764 dvdd.t1351 193.022
R5005 dvdd.t685 dvdd 192.569
R5006 dvdd.t995 dvdd 192.569
R5007 dvdd.t108 dvdd.t1468 191.344
R5008 dvdd.t1393 dvdd.t1497 191.344
R5009 dvdd.n143 dvdd.n142 190.165
R5010 dvdd.t709 dvdd 190
R5011 dvdd.t1603 dvdd.t68 189.665
R5012 dvdd.t669 dvdd 187.987
R5013 dvdd.n409 dvdd.n408 186.894
R5014 dvdd.n3088 dvdd.n3085 185
R5015 dvdd.n3089 dvdd.n3088 185
R5016 dvdd.n7 dvdd.n4 185
R5017 dvdd.n8 dvdd.n7 185
R5018 dvdd.n14 dvdd.n11 185
R5019 dvdd.n15 dvdd.n14 185
R5020 dvdd.n21 dvdd.n18 185
R5021 dvdd.n22 dvdd.n21 185
R5022 dvdd.n28 dvdd.n25 185
R5023 dvdd.n29 dvdd.n28 185
R5024 dvdd.n35 dvdd.n32 185
R5025 dvdd.n36 dvdd.n35 185
R5026 dvdd.n42 dvdd.n39 185
R5027 dvdd.n43 dvdd.n42 185
R5028 dvdd.n49 dvdd.n46 185
R5029 dvdd.n50 dvdd.n49 185
R5030 dvdd.n56 dvdd.n53 185
R5031 dvdd.n57 dvdd.n56 185
R5032 dvdd.n63 dvdd.n60 185
R5033 dvdd.n64 dvdd.n63 185
R5034 dvdd.n2713 dvdd.n2710 185
R5035 dvdd.n2714 dvdd.n2713 185
R5036 dvdd.n2706 dvdd.n2703 185
R5037 dvdd.n2707 dvdd.n2706 185
R5038 dvdd.n2699 dvdd.n2696 185
R5039 dvdd.n2700 dvdd.n2699 185
R5040 dvdd.n2692 dvdd.n2689 185
R5041 dvdd.n2693 dvdd.n2692 185
R5042 dvdd.n2685 dvdd.n2682 185
R5043 dvdd.n2686 dvdd.n2685 185
R5044 dvdd.n2678 dvdd.n2675 185
R5045 dvdd.n2679 dvdd.n2678 185
R5046 dvdd.n2671 dvdd.n2668 185
R5047 dvdd.n2672 dvdd.n2671 185
R5048 dvdd.n2664 dvdd.n2661 185
R5049 dvdd.n2665 dvdd.n2664 185
R5050 dvdd.n2657 dvdd.n2654 185
R5051 dvdd.n2658 dvdd.n2657 185
R5052 dvdd.n1244 dvdd 184.63
R5053 dvdd.t1666 dvdd 182.952
R5054 dvdd.t1606 dvdd 182.952
R5055 dvdd.t1561 dvdd 182.952
R5056 dvdd.t1609 dvdd 182.952
R5057 dvdd.t1612 dvdd 182.952
R5058 dvdd.n1529 dvdd 182.952
R5059 dvdd.t1628 dvdd 182.952
R5060 dvdd.t1534 dvdd 182.952
R5061 dvdd.t1655 dvdd 182.952
R5062 dvdd.t1553 dvdd 182.952
R5063 dvdd.t1710 dvdd 182.952
R5064 dvdd.t354 dvdd.t466 181.273
R5065 dvdd.t348 dvdd.t882 181.273
R5066 dvdd.t805 dvdd.t938 181.273
R5067 dvdd.t1346 dvdd.t334 181.273
R5068 dvdd.t247 dvdd.t249 181.273
R5069 dvdd.t843 dvdd.t254 181.273
R5070 dvdd.t364 dvdd.t313 181.273
R5071 dvdd.t1360 dvdd.t1288 180.129
R5072 dvdd.n408 dvdd 179.595
R5073 dvdd dvdd.n1683 179.595
R5074 dvdd dvdd.t77 177.916
R5075 dvdd.n3144 dvdd.t1423 175.306
R5076 dvdd.t532 dvdd.t378 174.559
R5077 dvdd.t242 dvdd.n3143 174.066
R5078 dvdd dvdd.t328 171.202
R5079 dvdd.n2846 dvdd.t274 171.054
R5080 dvdd.t88 dvdd 169.524
R5081 dvdd.t931 dvdd 169.524
R5082 dvdd.t892 dvdd.t92 169.524
R5083 dvdd.t832 dvdd.t520 167.845
R5084 dvdd.t630 dvdd.t1493 167.845
R5085 dvdd.t981 dvdd.t266 167.845
R5086 dvdd.t989 dvdd 167.845
R5087 dvdd.t374 dvdd.t614 166.167
R5088 dvdd.t872 dvdd.t646 166.167
R5089 dvdd.t1035 dvdd.t1034 166.167
R5090 dvdd.t1033 dvdd.t1018 166.167
R5091 dvdd.t650 dvdd.t921 166.167
R5092 dvdd.t408 dvdd.t1416 166.167
R5093 dvdd.t431 dvdd.t795 166.167
R5094 dvdd.t432 dvdd.t436 166.167
R5095 dvdd.t585 dvdd.t1128 166.167
R5096 dvdd.t23 dvdd.t1509 166.167
R5097 dvdd.t180 dvdd.t14 166.167
R5098 dvdd.t17 dvdd.t226 166.167
R5099 dvdd.t1066 dvdd.t1080 166.167
R5100 dvdd.t817 dvdd.t819 166.167
R5101 dvdd.t818 dvdd.t1521 166.167
R5102 dvdd.t1718 dvdd.t1031 164.488
R5103 dvdd.t1118 dvdd.t510 162.81
R5104 dvdd.t826 dvdd.t578 162.81
R5105 dvdd.t991 dvdd 162.81
R5106 dvdd.t1087 dvdd.t1173 162.81
R5107 dvdd.t1177 dvdd.t1511 162.81
R5108 dvdd.t810 dvdd.t1305 162.81
R5109 dvdd.t336 dvdd.t1183 162.81
R5110 dvdd.t1272 dvdd.t1265 161.131
R5111 dvdd.t548 dvdd.t1272 161.131
R5112 dvdd.t1161 dvdd.t542 161.131
R5113 dvdd.t608 dvdd.t387 161.131
R5114 dvdd.t1730 dvdd.t138 161.131
R5115 dvdd.t1252 dvdd.t1400 161.131
R5116 dvdd.t771 dvdd.t884 159.452
R5117 dvdd.t1489 dvdd.t1029 159.452
R5118 dvdd.t82 dvdd.t1350 159.452
R5119 dvdd.t1215 dvdd.t634 159.452
R5120 dvdd.t1740 dvdd.t656 159.452
R5121 dvdd.t654 dvdd.t660 159.452
R5122 dvdd.t742 dvdd.t1336 159.452
R5123 dvdd.t1438 dvdd.t632 159.452
R5124 dvdd.t1476 dvdd.t849 159.452
R5125 dvdd.t1513 dvdd.t1442 159.452
R5126 dvdd.t1023 dvdd.t989 159.452
R5127 dvdd.t1054 dvdd.t1730 157.774
R5128 dvdd.t1173 dvdd.t1177 157.774
R5129 dvdd.t449 dvdd.t1603 157.774
R5130 dvdd.t1528 dvdd.t588 157.774
R5131 dvdd.n70 dvdd.t1058 157.446
R5132 dvdd.n2651 dvdd.t624 157.446
R5133 dvdd.t544 dvdd.t767 156.095
R5134 dvdd.n525 dvdd.t342 156.095
R5135 dvdd.n814 dvdd.t352 156.095
R5136 dvdd.t1372 dvdd.t1113 156.095
R5137 dvdd.t679 dvdd.t1409 156.095
R5138 dvdd.t681 dvdd.t1438 156.095
R5139 dvdd.t1572 dvdd.t1724 154.417
R5140 dvdd.t1018 dvdd.t323 154.417
R5141 dvdd.t781 dvdd.t9 154.417
R5142 dvdd.t9 dvdd.t923 154.417
R5143 dvdd.t1221 dvdd.t408 154.417
R5144 dvdd.t1384 dvdd.t76 154.417
R5145 dvdd.t626 dvdd.t1051 154.417
R5146 dvdd.t436 dvdd.t1299 154.417
R5147 dvdd.t1312 dvdd.t1189 154.417
R5148 dvdd.t830 dvdd.t750 154.417
R5149 dvdd.t1090 dvdd.t764 154.417
R5150 dvdd.t1521 dvdd.t1015 154.417
R5151 dvdd.t1590 dvdd.t1765 154.417
R5152 dvdd.t437 dvdd.t616 154.417
R5153 dvdd.t894 dvdd.t735 154.417
R5154 dvdd.t404 dvdd.t824 154.417
R5155 dvdd.n145 dvdd.n144 152
R5156 dvdd.t1163 dvdd.t1750 151.06
R5157 dvdd.t1225 dvdd.t140 151.06
R5158 dvdd.t1661 dvdd.t574 151.06
R5159 dvdd.t762 dvdd.t26 149.382
R5160 dvdd.t86 dvdd.t1025 147.703
R5161 dvdd.t1479 dvdd.t1103 147.703
R5162 dvdd.t979 dvdd.t797 147.703
R5163 dvdd.t1130 dvdd.t857 147.703
R5164 dvdd.t588 dvdd.t1101 147.703
R5165 dvdd.n3062 dvdd.t963 146.351
R5166 dvdd.n3005 dvdd.t56 146.351
R5167 dvdd.n1633 dvdd.n1632 146.25
R5168 dvdd.t578 dvdd.t836 146.025
R5169 dvdd.t1421 dvdd.t1283 145.488
R5170 dvdd.t912 dvdd.t664 144.346
R5171 dvdd.t873 dvdd.t872 144.346
R5172 dvdd.t484 dvdd.t494 144.346
R5173 dvdd.t478 dvdd.t488 144.346
R5174 dvdd.t470 dvdd.t490 144.346
R5175 dvdd.t1452 dvdd.t1460 144.346
R5176 dvdd.t378 dvdd.t1274 144.346
R5177 dvdd.t915 dvdd.t1073 144.346
R5178 dvdd.t1319 dvdd 144.346
R5179 dvdd.t1470 dvdd.t630 144.346
R5180 dvdd.t1415 dvdd.t409 144.346
R5181 dvdd.t903 dvdd.t508 144.346
R5182 dvdd.t435 dvdd.t431 144.346
R5183 dvdd.t120 dvdd.t106 144.346
R5184 dvdd.t132 dvdd.t124 144.346
R5185 dvdd.t104 dvdd.t130 144.346
R5186 dvdd.t775 dvdd.t779 144.346
R5187 dvdd.t100 dvdd.t729 144.346
R5188 dvdd.t867 dvdd.t252 144.346
R5189 dvdd.t1079 dvdd.t1065 144.346
R5190 dvdd.t174 dvdd.t162 144.346
R5191 dvdd.t158 dvdd.t174 144.346
R5192 dvdd.t168 dvdd.t158 144.346
R5193 dvdd.t178 dvdd.t164 144.346
R5194 dvdd.t160 dvdd.t178 144.346
R5195 dvdd.t172 dvdd.t160 144.346
R5196 dvdd.t1417 dvdd 144.346
R5197 dvdd.n2042 dvdd.n2010 142.934
R5198 dvdd.t1334 dvdd.t726 142.668
R5199 dvdd.t488 dvdd.t476 142.668
R5200 dvdd.t496 dvdd.n813 142.668
R5201 dvdd.t1077 dvdd.t650 142.668
R5202 dvdd.t914 dvdd.t651 142.668
R5203 dvdd.t1382 dvdd.t1307 142.668
R5204 dvdd.t140 dvdd.t99 142.668
R5205 dvdd.t662 dvdd.t1066 142.668
R5206 dvdd.t1485 dvdd.t152 142.668
R5207 dvdd.n2908 dvdd.t200 141.868
R5208 dvdd.t460 dvdd.t464 140.989
R5209 dvdd.t464 dvdd.t462 140.989
R5210 dvdd.t1507 dvdd.t354 140.989
R5211 dvdd.t466 dvdd.t518 140.989
R5212 dvdd.t1159 dvdd.t544 140.989
R5213 dvdd.t1165 dvdd.t1167 140.989
R5214 dvdd.t615 dvdd.t1267 140.989
R5215 dvdd.t878 dvdd.t880 140.989
R5216 dvdd.t570 dvdd.t348 140.989
R5217 dvdd.t882 dvdd.t873 140.989
R5218 dvdd.t758 dvdd.t861 140.989
R5219 dvdd.t1269 dvdd.t769 140.989
R5220 dvdd.t358 dvdd.t636 140.989
R5221 dvdd.t1017 dvdd.t1069 140.989
R5222 dvdd.t1031 dvdd.t596 140.989
R5223 dvdd.t502 dvdd.t1109 140.989
R5224 dvdd.t791 dvdd.t832 140.989
R5225 dvdd.t230 dvdd.t8 140.989
R5226 dvdd.t1074 dvdd.t590 140.989
R5227 dvdd.t652 dvdd.t592 140.989
R5228 dvdd.t1150 dvdd.t366 140.989
R5229 dvdd.t929 dvdd.t606 140.989
R5230 dvdd.t334 dvdd.t719 140.989
R5231 dvdd.t1113 dvdd.t506 140.989
R5232 dvdd.t1049 dvdd.t435 140.989
R5233 dvdd.t582 dvdd.t580 140.989
R5234 dvdd.t102 dvdd.t1263 140.989
R5235 dvdd.t586 dvdd.t414 140.989
R5236 dvdd.t723 dvdd.t721 140.989
R5237 dvdd.t1001 dvdd.t1003 140.989
R5238 dvdd.t863 dvdd 140.989
R5239 dvdd.t138 dvdd.t144 140.989
R5240 dvdd.t1223 dvdd.t802 140.989
R5241 dvdd.t98 dvdd.t1390 140.989
R5242 dvdd.t396 dvdd.t12 140.989
R5243 dvdd.t1097 dvdd.t1179 140.989
R5244 dvdd.t1175 dvdd.t1085 140.989
R5245 dvdd.t21 dvdd.t425 140.989
R5246 dvdd.t256 dvdd.t80 140.989
R5247 dvdd.t254 dvdd.t1210 140.989
R5248 dvdd.t1210 dvdd.t847 140.989
R5249 dvdd.t1200 dvdd.t1079 140.989
R5250 dvdd.t1313 dvdd.t1315 140.989
R5251 dvdd.t1217 dvdd.t1215 140.989
R5252 dvdd.t656 dvdd.t654 140.989
R5253 dvdd.t1409 dvdd.t1407 140.989
R5254 dvdd.t1391 dvdd.t1444 140.989
R5255 dvdd.t92 dvdd.t677 140.989
R5256 dvdd.t1197 dvdd.t1449 140.989
R5257 dvdd.t675 dvdd.t944 140.989
R5258 dvdd.t4 dvdd.t2 140.989
R5259 dvdd.t1124 dvdd.t1126 140.989
R5260 dvdd.t803 dvdd.t1276 139.311
R5261 dvdd dvdd.t1021 139.311
R5262 dvdd.t923 dvdd.t1074 139.311
R5263 dvdd.t1405 dvdd.t393 139.311
R5264 dvdd.t1053 dvdd.t1245 139.311
R5265 dvdd.t1080 dvdd.t18 139.311
R5266 dvdd.t936 dvdd 139.311
R5267 dvdd.t767 dvdd.t572 137.633
R5268 dvdd.t1233 dvdd.t728 137.633
R5269 dvdd.t733 dvdd.t671 137.633
R5270 dvdd.n1569 dvdd.n1536 136.882
R5271 dvdd.t1356 dvdd.t1358 136.828
R5272 dvdd.t1354 dvdd.t1356 136.828
R5273 dvdd.t445 dvdd.t1354 136.828
R5274 dvdd.t443 dvdd.t445 136.828
R5275 dvdd.t447 dvdd.t443 136.828
R5276 dvdd.t1288 dvdd.t447 136.828
R5277 dvdd.t236 dvdd.t242 136.828
R5278 dvdd.t234 dvdd.t236 136.828
R5279 dvdd.t240 dvdd.t234 136.828
R5280 dvdd.t244 dvdd.t240 136.828
R5281 dvdd.t238 dvdd.t244 136.828
R5282 dvdd.t1440 dvdd.t892 135.954
R5283 dvdd.t871 dvdd.t480 134.276
R5284 dvdd dvdd.t1346 134.276
R5285 dvdd.t74 dvdd.t801 134.276
R5286 dvdd.t875 dvdd.t519 132.597
R5287 dvdd.t886 dvdd.t1318 132.597
R5288 dvdd.t1366 dvdd.t1111 132.597
R5289 dvdd.t756 dvdd.t122 132.597
R5290 dvdd.t142 dvdd.t406 132.597
R5291 dvdd.t834 dvdd.t1067 132.597
R5292 dvdd.t1652 dvdd.t1520 132.597
R5293 dvdd.t1169 dvdd.t546 130.919
R5294 dvdd.t372 dvdd.t725 130.919
R5295 dvdd.t534 dvdd.t474 130.919
R5296 dvdd.t330 dvdd.t806 130.919
R5297 dvdd.t828 dvdd 130.919
R5298 dvdd.t1121 dvdd.t166 130.919
R5299 dvdd.t156 dvdd.t1083 130.919
R5300 dvdd dvdd.t1447 130.919
R5301 dvdd.t1204 dvdd.n3087 129.546
R5302 dvdd.t919 dvdd.n6 129.546
R5303 dvdd.t1231 dvdd.n13 129.546
R5304 dvdd.t1212 dvdd.n20 129.546
R5305 dvdd.t1140 dvdd.n27 129.546
R5306 dvdd.t1250 dvdd.n34 129.546
R5307 dvdd.t1385 dvdd.n41 129.546
R5308 dvdd.t429 dvdd.n48 129.546
R5309 dvdd.t576 dvdd.n55 129.546
R5310 dvdd.t34 dvdd.n62 129.546
R5311 dvdd.t917 dvdd.n2712 129.546
R5312 dvdd.t787 dvdd.n2705 129.546
R5313 dvdd.t1261 dvdd.n2698 129.546
R5314 dvdd.t1138 dvdd.n2691 129.546
R5315 dvdd.t410 dvdd.n2684 129.546
R5316 dvdd.t1483 dvdd.n2677 129.546
R5317 dvdd.t514 dvdd.n2670 129.546
R5318 dvdd.t228 dvdd.n2663 129.546
R5319 dvdd.t94 dvdd.n2656 129.546
R5320 dvdd.n1512 dvdd.t1878 129.344
R5321 dvdd.n1828 dvdd.t1826 129.344
R5322 dvdd.n2596 dvdd.t1902 129.344
R5323 dvdd.n2608 dvdd.t1862 129.344
R5324 dvdd.n525 dvdd 129.24
R5325 dvdd.t1460 dvdd.t766 129.24
R5326 dvdd.t1317 dvdd.t457 129.24
R5327 dvdd.t1132 dvdd.t673 129.24
R5328 dvdd.t1061 dvdd.n67 127.638
R5329 dvdd.t899 dvdd.n2648 127.638
R5330 dvdd.t821 dvdd.t877 127.562
R5331 dvdd.n524 dvdd 127.562
R5332 dvdd.t542 dvdd.t1071 127.562
R5333 dvdd.t717 dvdd.t845 127.562
R5334 dvdd.t740 dvdd.t731 127.562
R5335 dvdd.t1646 dvdd 125.883
R5336 dvdd.n408 dvdd 125.883
R5337 dvdd.t1540 dvdd 125.883
R5338 dvdd.n814 dvdd 125.883
R5339 dvdd.t1578 dvdd 125.883
R5340 dvdd.n944 dvdd 125.883
R5341 dvdd dvdd.t28 125.883
R5342 dvdd.n1101 dvdd 125.883
R5343 dvdd.t1583 dvdd 125.883
R5344 dvdd.t362 dvdd.t403 125.883
R5345 dvdd.t1600 dvdd 125.883
R5346 dvdd.n1529 dvdd 125.883
R5347 dvdd.n1684 dvdd 125.883
R5348 dvdd.t1721 dvdd 125.883
R5349 dvdd.n1826 dvdd 125.883
R5350 dvdd.t1007 dvdd.t412 125.883
R5351 dvdd.t154 dvdd.t789 125.883
R5352 dvdd dvdd.t170 125.883
R5353 dvdd.t1700 dvdd 125.883
R5354 dvdd.n2448 dvdd 125.883
R5355 dvdd.n2556 dvdd 125.883
R5356 dvdd dvdd.t482 124.206
R5357 dvdd.t387 dvdd.t640 124.206
R5358 dvdd.t1311 dvdd.t1327 124.206
R5359 dvdd.t1411 dvdd.t1389 124.206
R5360 dvdd.t799 dvdd.t1481 124.206
R5361 dvdd.n2555 dvdd 124.206
R5362 dvdd.n753 dvdd.t535 123.507
R5363 dvdd.t614 dvdd.t512 122.526
R5364 dvdd.n1244 dvdd 122.526
R5365 dvdd dvdd.t102 122.526
R5366 dvdd.n1387 dvdd.t400 122.526
R5367 dvdd.t1146 dvdd.t247 122.526
R5368 dvdd.t877 dvdd.t1013 120.849
R5369 dvdd.t1069 dvdd 120.849
R5370 dvdd.t1117 dvdd 120.849
R5371 dvdd.t84 dvdd.t1381 120.849
R5372 dvdd.t309 dvdd.t805 120.849
R5373 dvdd.t389 dvdd.t1487 120.849
R5374 dvdd dvdd.t1049 120.849
R5375 dvdd.t752 dvdd.t1235 120.849
R5376 dvdd.t32 dvdd.t110 120.849
R5377 dvdd.t77 dvdd.t810 120.849
R5378 dvdd.t1009 dvdd.t1010 120.849
R5379 dvdd.n356 dvdd.t467 119.608
R5380 dvdd.n339 dvdd.t1268 119.608
R5381 dvdd.n638 dvdd.t883 119.608
R5382 dvdd.n620 dvdd.t1070 119.608
R5383 dvdd.n942 dvdd.t718 119.608
R5384 dvdd.n1002 dvdd.t231 119.608
R5385 dvdd.n1059 dvdd.t329 119.608
R5386 dvdd.n1119 dvdd.t1347 119.608
R5387 dvdd.n1237 dvdd.t1050 119.608
R5388 dvdd.n1215 dvdd.t643 119.608
R5389 dvdd.n1393 dvdd.t1038 119.608
R5390 dvdd.n1506 dvdd.t1224 119.608
R5391 dvdd.n1693 dvdd.t399 119.608
R5392 dvdd.n1703 dvdd.t1341 119.608
R5393 dvdd.n1822 dvdd.t255 119.608
R5394 dvdd.n1819 dvdd.t1201 119.608
R5395 dvdd.n1935 dvdd.t452 119.608
R5396 dvdd.n1994 dvdd.t314 119.608
R5397 dvdd.t884 dvdd.t516 119.171
R5398 dvdd.t1152 dvdd 119.171
R5399 dvdd.t904 dvdd.t1107 119.171
R5400 dvdd dvdd.t1504 119.171
R5401 dvdd.n1993 dvdd.t364 119.171
R5402 dvdd.n2170 dvdd.t1861 119.007
R5403 dvdd.n1526 dvdd.t1825 118.853
R5404 dvdd.n2153 dvdd.t1854 118.853
R5405 dvdd.t1293 dvdd.t1421 117.776
R5406 dvdd dvdd.t610 117.492
R5407 dvdd.t1259 dvdd.t983 117.492
R5408 dvdd.t80 dvdd 117.492
R5409 dvdd.n764 dvdd.t1275 117.451
R5410 dvdd.n1247 dvdd.t1371 117.451
R5411 dvdd.n668 dvdd.t1906 117.294
R5412 dvdd.n1155 dvdd.t1833 117.294
R5413 dvdd.n2428 dvdd.t1896 117.294
R5414 dvdd.n927 dvdd.t1240 116.341
R5415 dvdd.n1533 dvdd.t143 116.341
R5416 dvdd.t1207 dvdd 115.814
R5417 dvdd dvdd.t1206 115.814
R5418 dvdd.t1502 dvdd.t1393 115.814
R5419 dvdd.n2165 dvdd.t1835 115.109
R5420 dvdd.t754 dvdd.t381 114.135
R5421 dvdd.t260 dvdd.t1349 114.135
R5422 dvdd.t439 dvdd.t942 112.457
R5423 dvdd.t874 dvdd.t492 112.457
R5424 dvdd.t1404 dvdd.t1489 112.457
R5425 dvdd.t458 dvdd 112.457
R5426 dvdd dvdd.t1056 112.457
R5427 dvdd.t128 dvdd.t1395 112.457
R5428 dvdd.t721 dvdd 112.457
R5429 dvdd.t144 dvdd 112.457
R5430 dvdd.t1126 dvdd 112.457
R5431 dvdd.t1271 dvdd.t540 110.778
R5432 dvdd.t1239 dvdd.t1332 110.778
R5433 dvdd dvdd.t30 110.778
R5434 dvdd.t1037 dvdd.t860 110.778
R5435 dvdd dvdd.t455 110.778
R5436 dvdd.t1336 dvdd 110.778
R5437 dvdd.t1285 dvdd.t238 109.983
R5438 dvdd.t1283 dvdd.t823 109.983
R5439 dvdd dvdd.t602 109.1
R5440 dvdd.t594 dvdd 109.1
R5441 dvdd dvdd.t1163 109.1
R5442 dvdd.t596 dvdd 109.1
R5443 dvdd dvdd.t855 109.1
R5444 dvdd.t590 dvdd 109.1
R5445 dvdd.t592 dvdd 109.1
R5446 dvdd dvdd.t385 109.1
R5447 dvdd dvdd.t1470 109.1
R5448 dvdd.t1103 dvdd 109.1
R5449 dvdd dvdd.t1297 109.1
R5450 dvdd.t321 dvdd.t104 109.1
R5451 dvdd dvdd.t526 109.1
R5452 dvdd.t1148 dvdd.t362 109.1
R5453 dvdd dvdd.t865 109.1
R5454 dvdd dvdd.t420 109.1
R5455 dvdd.t425 dvdd 109.1
R5456 dvdd.t412 dvdd 109.1
R5457 dvdd.t418 dvdd 109.1
R5458 dvdd.t1081 dvdd.t154 109.1
R5459 dvdd dvdd.t427 109.1
R5460 dvdd.t416 dvdd 109.1
R5461 dvdd.t574 dvdd 109.1
R5462 dvdd.t634 dvdd 109.1
R5463 dvdd.t660 dvdd 109.1
R5464 dvdd.t1338 dvdd 109.1
R5465 dvdd dvdd.t851 109.1
R5466 dvdd.t1101 dvdd 109.1
R5467 dvdd dvdd.t1278 107.421
R5468 dvdd.t1193 dvdd 107.421
R5469 dvdd dvdd.t86 107.421
R5470 dvdd dvdd.t309 107.421
R5471 dvdd.t1491 dvdd 107.421
R5472 dvdd.t1235 dvdd 107.421
R5473 dvdd.t905 dvdd.t332 107.421
R5474 dvdd dvdd.t250 107.421
R5475 dvdd dvdd.t391 107.421
R5476 dvdd dvdd.t90 107.421
R5477 dvdd.t1227 dvdd 107.421
R5478 dvdd.n2555 dvdd.n2554 106.559
R5479 dvdd dvdd.t1430 106.543
R5480 dvdd dvdd.t1572 105.743
R5481 dvdd.t1634 dvdd 105.743
R5482 dvdd.t1209 dvdd.t658 105.743
R5483 dvdd.t26 dvdd 105.743
R5484 dvdd.t859 dvdd 105.743
R5485 dvdd dvdd.t628 105.743
R5486 dvdd dvdd.t783 105.743
R5487 dvdd.t462 dvdd.t1789 104.064
R5488 dvdd.t1368 dvdd.t1295 104.064
R5489 dvdd dvdd.t604 104.064
R5490 dvdd dvdd.t1093 104.064
R5491 dvdd.t0 dvdd.t932 104.064
R5492 dvdd.t1500 dvdd 104.064
R5493 dvdd dvdd.t1377 104.064
R5494 dvdd.t908 dvdd 104.064
R5495 dvdd dvdd.t1158 103.584
R5496 dvdd.t1156 dvdd.t370 102.385
R5497 dvdd.t380 dvdd.t346 102.385
R5498 dvdd.t524 dvdd.t478 102.385
R5499 dvdd.t598 dvdd 102.385
R5500 dvdd.n1100 dvdd.t1318 102.385
R5501 dvdd.t1005 dvdd.t813 102.385
R5502 dvdd.t1426 dvdd 102.385
R5503 dvdd.t1402 dvdd 102.385
R5504 dvdd.t319 dvdd.t118 102.385
R5505 dvdd.t910 dvdd.t773 102.385
R5506 dvdd.t1011 dvdd 102.385
R5507 dvdd.t136 dvdd.t1502 102.385
R5508 dvdd dvdd.t1637 102.385
R5509 dvdd dvdd.t96 102.385
R5510 dvdd.t96 dvdd.t1202 102.385
R5511 dvdd dvdd.t449 102.385
R5512 dvdd.t1122 dvdd.t150 102.385
R5513 dvdd.t1171 dvdd 102.385
R5514 dvdd.t1181 dvdd 102.385
R5515 dvdd.n3090 dvdd.n3085 101.644
R5516 dvdd.n9 dvdd.n4 101.644
R5517 dvdd.n16 dvdd.n11 101.644
R5518 dvdd.n23 dvdd.n18 101.644
R5519 dvdd.n30 dvdd.n25 101.644
R5520 dvdd.n37 dvdd.n32 101.644
R5521 dvdd.n44 dvdd.n39 101.644
R5522 dvdd.n51 dvdd.n46 101.644
R5523 dvdd.n58 dvdd.n53 101.644
R5524 dvdd.n65 dvdd.n60 101.644
R5525 dvdd.n2715 dvdd.n2710 101.644
R5526 dvdd.n2708 dvdd.n2703 101.644
R5527 dvdd.n2701 dvdd.n2696 101.644
R5528 dvdd.n2694 dvdd.n2689 101.644
R5529 dvdd.n2687 dvdd.n2682 101.644
R5530 dvdd.n2680 dvdd.n2675 101.644
R5531 dvdd.n2673 dvdd.n2668 101.644
R5532 dvdd.n2666 dvdd.n2661 101.644
R5533 dvdd.n2659 dvdd.n2654 101.644
R5534 dvdd.t526 dvdd.t1039 100.707
R5535 dvdd.t1351 dvdd.t311 100.707
R5536 dvdd.t264 dvdd.t1090 100.707
R5537 dvdd.t838 dvdd.t1374 100.707
R5538 dvdd.t338 dvdd.t472 99.0288
R5539 dvdd.t1575 dvdd.t1017 99.0288
R5540 dvdd.t715 dvdd 99.0288
R5541 dvdd.t748 dvdd.t828 99.0288
R5542 dvdd.n2016 dvdd.t1482 98.5005
R5543 dvdd.t550 dvdd.t383 97.3503
R5544 dvdd.t987 dvdd 97.3503
R5545 dvdd.t1301 dvdd 97.3503
R5546 dvdd dvdd.t453 97.3503
R5547 dvdd.t1063 dvdd 97.3503
R5548 dvdd.t1450 dvdd.t841 97.3503
R5549 dvdd.n763 dvdd.t87 96.1553
R5550 dvdd.n967 dvdd.t511 96.1553
R5551 dvdd.n1831 dvdd.t811 96.1553
R5552 dvdd.n2013 dvdd.t147 96.1553
R5553 dvdd.n2112 dvdd.t738 96.1553
R5554 dvdd.n2560 dvdd.t1448 96.1553
R5555 dvdd.n2562 dvdd.t670 96.1553
R5556 dvdd.n2763 dvdd.n67 95.8438
R5557 dvdd.n2755 dvdd.n2648 95.8438
R5558 dvdd dvdd.t441 95.6719
R5559 dvdd.t1325 dvdd.t615 95.6719
R5560 dvdd.t1144 dvdd 95.6719
R5561 dvdd.t932 dvdd.t394 95.6719
R5562 dvdd.t815 dvdd 95.6719
R5563 dvdd.n1658 dvdd.n1657 94.5605
R5564 dvdd dvdd.t439 93.9934
R5565 dvdd dvdd.t440 93.9934
R5566 dvdd.t114 dvdd.t1043 93.9934
R5567 dvdd.t126 dvdd.t1047 93.9934
R5568 dvdd.t112 dvdd.t1041 93.9934
R5569 dvdd.t124 dvdd.t1045 93.9934
R5570 dvdd.t584 dvdd 93.9934
R5571 dvdd.t528 dvdd.t398 93.9934
R5572 dvdd.t1340 dvdd.t1019 93.9934
R5573 dvdd.t1456 dvdd.t317 93.9934
R5574 dvdd dvdd.t817 93.9934
R5575 dvdd.n350 dvdd.t1324 93.81
R5576 dvdd.n465 dvdd.t768 93.81
R5577 dvdd.n526 dvdd.t897 93.81
R5578 dvdd.n634 dvdd.t649 93.81
R5579 dvdd.n817 dvdd.t1022 93.81
R5580 dvdd.n937 dvdd.t579 93.81
R5581 dvdd.n1015 dvdd.t305 93.81
R5582 dvdd.n1054 dvdd.t1153 93.81
R5583 dvdd.n1062 dvdd.t1490 93.81
R5584 dvdd.n1114 dvdd.t1281 93.81
R5585 dvdd.n1218 dvdd.t31 93.81
R5586 dvdd.n1233 dvdd.t1135 93.81
R5587 dvdd.n1243 dvdd.t1373 93.81
R5588 dvdd.n1330 dvdd.t757 93.81
R5589 dvdd.n1392 dvdd.t1149 93.81
R5590 dvdd.n1399 dvdd.t1310 93.81
R5591 dvdd.n1628 dvdd.t809 93.81
R5592 dvdd.n1696 dvdd.t1088 93.81
R5593 dvdd.n1697 dvdd.t1512 93.81
R5594 dvdd.n1889 dvdd.t786 93.81
R5595 dvdd.n1897 dvdd.t1304 93.81
R5596 dvdd.n1943 dvdd.t790 93.81
R5597 dvdd.n2002 dvdd.t1184 93.81
R5598 dvdd.n2388 dvdd.t743 93.81
R5599 dvdd.n2505 dvdd.t1439 93.81
R5600 dvdd.n2504 dvdd.t1446 93.81
R5601 dvdd.n2514 dvdd.t736 93.81
R5602 dvdd.n3090 dvdd.n3089 92.5005
R5603 dvdd.n69 dvdd.n68 92.5005
R5604 dvdd.n9 dvdd.n8 92.5005
R5605 dvdd.n16 dvdd.n15 92.5005
R5606 dvdd.n23 dvdd.n22 92.5005
R5607 dvdd.n30 dvdd.n29 92.5005
R5608 dvdd.n37 dvdd.n36 92.5005
R5609 dvdd.n44 dvdd.n43 92.5005
R5610 dvdd.n51 dvdd.n50 92.5005
R5611 dvdd.n58 dvdd.n57 92.5005
R5612 dvdd.n65 dvdd.n64 92.5005
R5613 dvdd.n2650 dvdd.n2649 92.5005
R5614 dvdd.n2715 dvdd.n2714 92.5005
R5615 dvdd.n2708 dvdd.n2707 92.5005
R5616 dvdd.n2701 dvdd.n2700 92.5005
R5617 dvdd.n2694 dvdd.n2693 92.5005
R5618 dvdd.n2687 dvdd.n2686 92.5005
R5619 dvdd.n2680 dvdd.n2679 92.5005
R5620 dvdd.n2673 dvdd.n2672 92.5005
R5621 dvdd.n2666 dvdd.n2665 92.5005
R5622 dvdd.n2659 dvdd.n2658 92.5005
R5623 dvdd.t1195 dvdd.t496 92.315
R5624 dvdd.t304 dvdd.t914 92.315
R5625 dvdd.t1241 dvdd.t246 92.315
R5626 dvdd.t802 dvdd.t258 92.315
R5627 dvdd.t1303 dvdd.t662 92.315
R5628 dvdd.t1428 dvdd 91.745
R5629 dvdd.t72 dvdd.t1152 90.6365
R5630 dvdd dvdd.t360 90.6365
R5631 dvdd.t423 dvdd.t1309 90.6365
R5632 dvdd dvdd.t1092 90.6365
R5633 dvdd.t1115 dvdd 88.9581
R5634 dvdd.t600 dvdd.t500 88.9581
R5635 dvdd.t836 dvdd.t1076 88.9581
R5636 dvdd.t328 dvdd.t940 88.9581
R5637 dvdd dvdd.t1243 88.9581
R5638 dvdd dvdd.t1229 88.9581
R5639 dvdd.t1095 dvdd.t644 88.9581
R5640 dvdd.t1280 dvdd.t1658 87.2797
R5641 dvdd.t1569 dvdd.t1134 87.2797
R5642 dvdd.n1386 dvdd.t1257 87.2797
R5643 dvdd.t1179 dvdd.t528 87.2797
R5644 dvdd.t1019 dvdd.t1175 87.2797
R5645 dvdd.t1690 dvdd.t1023 87.2797
R5646 dvdd.n760 dvdd.t621 86.7743
R5647 dvdd.n767 dvdd.t379 86.7743
R5648 dvdd.n767 dvdd.t533 86.7743
R5649 dvdd.n1251 dvdd.t1112 86.7743
R5650 dvdd.n1251 dvdd.t814 86.7743
R5651 dvdd.t869 dvdd.t486 85.6012
R5652 dvdd.t1478 dvdd.t1452 85.6012
R5653 dvdd.t1329 dvdd.t777 85.6012
R5654 dvdd.t945 dvdd.t15 85.6012
R5655 dvdd.t20 dvdd.t10 85.6012
R5656 dvdd.t342 dvdd.t1154 83.9228
R5657 dvdd.t268 dvdd.t1695 83.9228
R5658 dvdd.t451 dvdd.t1450 83.9228
R5659 dvdd dvdd.t744 83.9228
R5660 dvdd.t823 dvdd.t1285 83.1363
R5661 dvdd.n69 dvdd.n67 82.3534
R5662 dvdd.n2650 dvdd.n2648 82.3534
R5663 dvdd.t1013 dvdd.t350 82.2443
R5664 dvdd.t1454 dvdd.t620 82.2443
R5665 dvdd.t1682 dvdd.t1117 82.2443
R5666 dvdd dvdd.t775 82.2443
R5667 dvdd.t1495 dvdd.t638 82.2443
R5668 dvdd.t6 dvdd 80.5659
R5669 dvdd.t648 dvdd.t484 80.5659
R5670 dvdd.n944 dvdd.t715 80.5659
R5671 dvdd.n1684 dvdd.t1500 80.5659
R5672 dvdd.t11 dvdd.t945 80.5659
R5673 dvdd.t10 dvdd.t946 80.5659
R5674 dvdd.t1120 dvdd.t1458 80.5659
R5675 dvdd.t1082 dvdd.t176 80.5659
R5676 dvdd.t1773 dvdd.t746 80.5659
R5677 dvdd.t1525 dvdd.t1476 80.5659
R5678 dvdd.t1267 dvdd.t380 78.8874
R5679 dvdd.t1154 dvdd.t896 78.8874
R5680 dvdd.t536 dvdd.t1454 78.8874
R5681 dvdd.t925 dvdd.t82 78.8874
R5682 dvdd.t1423 dvdd.t1293 78.8063
R5683 dvdd.n2614 dvdd.t1516 77.3934
R5684 dvdd.n2520 dvdd.t745 77.3934
R5685 dvdd.n2516 dvdd.t895 77.3934
R5686 dvdd.n2526 dvdd.t784 77.3934
R5687 dvdd.n2524 dvdd.t1096 77.3934
R5688 dvdd.n2365 dvdd.t674 77.3934
R5689 dvdd.n2369 dvdd.t1418 77.3934
R5690 dvdd.n2572 dvdd.t990 77.3934
R5691 dvdd.n2569 dvdd.t1443 77.3934
R5692 dvdd.n646 dvdd.t1687 77.209
R5693 dvdd.t1390 dvdd.t808 77.209
R5694 dvdd.n3087 dvdd.n3086 77.057
R5695 dvdd.n6 dvdd.n5 77.057
R5696 dvdd.n13 dvdd.n12 77.057
R5697 dvdd.n20 dvdd.n19 77.057
R5698 dvdd.n27 dvdd.n26 77.057
R5699 dvdd.n34 dvdd.n33 77.057
R5700 dvdd.n41 dvdd.n40 77.057
R5701 dvdd.n48 dvdd.n47 77.057
R5702 dvdd.n55 dvdd.n54 77.057
R5703 dvdd.n62 dvdd.n61 77.057
R5704 dvdd.n2712 dvdd.n2711 77.057
R5705 dvdd.n2705 dvdd.n2704 77.057
R5706 dvdd.n2698 dvdd.n2697 77.057
R5707 dvdd.n2691 dvdd.n2690 77.057
R5708 dvdd.n2684 dvdd.n2683 77.057
R5709 dvdd.n2677 dvdd.n2676 77.057
R5710 dvdd.n2670 dvdd.n2669 77.057
R5711 dvdd.n2663 dvdd.n2662 77.057
R5712 dvdd.n2656 dvdd.n2655 77.057
R5713 dvdd.n2145 dvdd.n2124 76.0729
R5714 dvdd.t1658 dvdd.t356 75.5305
R5715 dvdd.t340 dvdd.t1569 75.5305
R5716 dvdd.t638 dvdd.t608 75.5305
R5717 dvdd.t801 dvdd 75.5305
R5718 dvdd.n649 dvdd.t935 75.0481
R5719 dvdd.n977 dvdd.t271 75.0481
R5720 dvdd.n1405 dvdd.t1186 75.0481
R5721 dvdd.n1493 dvdd.t928 75.0481
R5722 dvdd.n1637 dvdd.t137 75.0481
R5723 dvdd.n1585 dvdd.t1100 75.0481
R5724 dvdd.n1989 dvdd.t1378 75.0481
R5725 dvdd.n2115 dvdd.t326 75.0481
R5726 dvdd.n2267 dvdd.n2229 74.7537
R5727 dvdd.t1076 dvdd.t304 73.8521
R5728 dvdd.t642 dvdd.t905 73.8521
R5729 dvdd.n2227 dvdd.n2226 73.3193
R5730 dvdd.t519 dvdd 72.1736
R5731 dvdd.t636 dvdd.t1161 72.1736
R5732 dvdd.t368 dvdd.t72 72.1736
R5733 dvdd dvdd.t108 72.1736
R5734 dvdd.t344 dvdd.t423 72.1736
R5735 dvdd dvdd.t1312 72.1736
R5736 dvdd.t414 dvdd.t1198 72.1736
R5737 dvdd.n2908 dvdd.t208 70.9338
R5738 dvdd.t1332 dvdd.t376 70.4952
R5739 dvdd.t644 dvdd.t936 70.4952
R5740 dvdd.t783 dvdd.t1095 70.4952
R5741 dvdd.n474 dvdd.t541 69.9355
R5742 dvdd.n1504 dvdd.t751 69.9355
R5743 dvdd.n3062 dvdd.t971 69.3248
R5744 dvdd.n3005 dvdd.t64 69.3248
R5745 dvdd.t610 dvdd.t368 68.8168
R5746 dvdd.t30 dvdd.n1386 68.8168
R5747 dvdd.t401 dvdd.t344 68.8168
R5748 dvdd.t793 dvdd.t1543 68.8168
R5749 dvdd.t1375 dvdd.t1631 68.8168
R5750 dvdd.n1345 dvdd.t320 68.6784
R5751 dvdd.n1345 dvdd.t322 68.6784
R5752 dvdd.n760 dvdd.t537 68.0124
R5753 dvdd.n3088 dvdd.t1204 67.8576
R5754 dvdd.n7 dvdd.t919 67.8576
R5755 dvdd.n14 dvdd.t1231 67.8576
R5756 dvdd.n21 dvdd.t1212 67.8576
R5757 dvdd.n28 dvdd.t1140 67.8576
R5758 dvdd.n35 dvdd.t1250 67.8576
R5759 dvdd.n42 dvdd.t1385 67.8576
R5760 dvdd.n49 dvdd.t429 67.8576
R5761 dvdd.n56 dvdd.t576 67.8576
R5762 dvdd.n63 dvdd.t34 67.8576
R5763 dvdd.n2713 dvdd.t917 67.8576
R5764 dvdd.n2706 dvdd.t787 67.8576
R5765 dvdd.n2699 dvdd.t1261 67.8576
R5766 dvdd.n2692 dvdd.t1138 67.8576
R5767 dvdd.n2685 dvdd.t410 67.8576
R5768 dvdd.n2678 dvdd.t1483 67.8576
R5769 dvdd.n2671 dvdd.t514 67.8576
R5770 dvdd.n2664 dvdd.t228 67.8576
R5771 dvdd.n2657 dvdd.t94 67.8576
R5772 dvdd.t99 dvdd.t1411 67.1383
R5773 dvdd.t851 dvdd.t1417 67.1383
R5774 dvdd dvdd.t1513 67.1383
R5775 dvdd.t896 dvdd.t1334 65.4599
R5776 dvdd.t134 dvdd.t84 65.4599
R5777 dvdd dvdd.t929 65.4599
R5778 dvdd.t1330 dvdd 65.4599
R5779 dvdd.t16 dvdd.t838 65.4599
R5780 dvdd.t383 dvdd.t1169 63.7814
R5781 dvdd.t472 dvdd.t648 63.7814
R5782 dvdd.t1206 dvdd.n1100 63.7814
R5783 dvdd.t808 dvdd.t748 63.7814
R5784 dvdd.t176 dvdd.t1120 63.7814
R5785 dvdd.t150 dvdd.t1082 63.7814
R5786 dvdd.n356 dvdd.t355 63.3219
R5787 dvdd.n350 dvdd.t351 63.3219
R5788 dvdd.n469 dvdd.t545 63.3219
R5789 dvdd.n469 dvdd.t1160 63.3219
R5790 dvdd.n339 dvdd.t347 63.3219
R5791 dvdd.n526 dvdd.t343 63.3219
R5792 dvdd.n634 dvdd.t339 63.3219
R5793 dvdd.n638 dvdd.t349 63.3219
R5794 dvdd.n676 dvdd.t1116 63.3219
R5795 dvdd.n676 dvdd.t613 63.3219
R5796 dvdd.n620 dvdd.t359 63.3219
R5797 dvdd.n817 dvdd.t353 63.3219
R5798 dvdd.n947 dvdd.t623 63.3219
R5799 dvdd.n947 dvdd.t1369 63.3219
R5800 dvdd.n942 dvdd.t833 63.3219
R5801 dvdd.n1002 dvdd.t846 63.3219
R5802 dvdd.n937 dvdd.t827 63.3219
R5803 dvdd.n1015 dvdd.t837 63.3219
R5804 dvdd.n1054 dvdd.t369 63.3219
R5805 dvdd.n1059 dvdd.t367 63.3219
R5806 dvdd.n1065 dvdd.t984 63.3219
R5807 dvdd.n1065 dvdd.t386 63.3219
R5808 dvdd.n1114 dvdd.t357 63.3219
R5809 dvdd.n1119 dvdd.t335 63.3219
R5810 dvdd.n1220 dvdd.t1403 63.3219
R5811 dvdd.n1220 dvdd.t1258 63.3219
R5812 dvdd.n1233 dvdd.t341 63.3219
R5813 dvdd.n1237 dvdd.t361 63.3219
R5814 dvdd.n1240 dvdd.t1114 63.3219
R5815 dvdd.n1240 dvdd.t507 63.3219
R5816 dvdd.n1327 dvdd.t1256 63.3219
R5817 dvdd.n1327 dvdd.t33 63.3219
R5818 dvdd.n1215 dvdd.t333 63.3219
R5819 dvdd.n1392 dvdd.t331 63.3219
R5820 dvdd.n1393 dvdd.t363 63.3219
R5821 dvdd.n1399 dvdd.t345 63.3219
R5822 dvdd.n1409 dvdd.t1199 63.3219
R5823 dvdd.n1409 dvdd.t1344 63.3219
R5824 dvdd.n1528 dvdd.t1244 63.3219
R5825 dvdd.n1528 dvdd.t794 63.3219
R5826 dvdd.n1498 dvdd.t926 63.3219
R5827 dvdd.n1498 dvdd.t263 63.3219
R5828 dvdd.n1645 dvdd.t395 63.3219
R5829 dvdd.n1645 dvdd.t1 63.3219
R5830 dvdd.n1628 dvdd.t829 63.3219
R5831 dvdd.n1506 dvdd.t831 63.3219
R5832 dvdd.n1693 dvdd.t1180 63.3219
R5833 dvdd.n1696 dvdd.t1174 63.3219
R5834 dvdd.n1697 dvdd.t1178 63.3219
R5835 dvdd.n1703 dvdd.t1176 63.3219
R5836 dvdd.n1822 dvdd.t844 63.3219
R5837 dvdd.n1819 dvdd.t848 63.3219
R5838 dvdd.n1889 dvdd.t835 63.3219
R5839 dvdd.n1897 dvdd.t839 63.3219
R5840 dvdd.n1810 dvdd.t1230 63.3219
R5841 dvdd.n1810 dvdd.t1376 63.3219
R5842 dvdd.n1935 dvdd.t842 63.3219
R5843 dvdd.n1943 dvdd.t840 63.3219
R5844 dvdd.n1994 dvdd.t365 63.3219
R5845 dvdd.n2002 dvdd.t337 63.3219
R5846 dvdd.n2119 dvdd.t1499 63.3219
R5847 dvdd.n2119 dvdd.t916 63.3219
R5848 dvdd.n2491 dvdd.t1392 63.3219
R5849 dvdd.n2491 dvdd.t1445 63.3219
R5850 dvdd.n2506 dvdd.t672 63.3219
R5851 dvdd.n2506 dvdd.t629 63.3219
R5852 dvdd.n2508 dvdd.t682 63.3219
R5853 dvdd.n2508 dvdd.t734 63.3219
R5854 dvdd.n2519 dvdd.t678 63.3219
R5855 dvdd.n2519 dvdd.t93 63.3219
R5856 dvdd dvdd.t1165 62.103
R5857 dvdd.t620 dvdd.t1464 62.103
R5858 dvdd.t1089 dvdd 62.103
R5859 dvdd.t1374 dvdd.t1303 62.103
R5860 dvdd.n474 dvdd.t1166 62.0555
R5861 dvdd.n1536 dvdd.t1192 60.9739
R5862 dvdd dvdd.t358 60.4245
R5863 dvdd.t1109 dvdd 60.4245
R5864 dvdd.t1295 dvdd 60.4245
R5865 dvdd.t360 dvdd 60.4245
R5866 dvdd.t865 dvdd.t1241 60.4245
R5867 dvdd.t398 dvdd.t11 60.4245
R5868 dvdd.t946 dvdd.t1340 60.4245
R5869 dvdd.t1458 dvdd.t451 60.4245
R5870 dvdd.n1632 dvdd.t765 60.0855
R5871 dvdd.n1632 dvdd.t265 60.0855
R5872 dvdd.n1536 dvdd.t407 59.9892
R5873 dvdd dvdd.t375 58.7461
R5874 dvdd.t476 dvdd.t869 58.7461
R5875 dvdd.t1464 dvdd.t1478 58.7461
R5876 dvdd dvdd.t1118 58.7461
R5877 dvdd dvdd.t652 58.7461
R5878 dvdd.t938 dvdd.t1150 58.7461
R5879 dvdd dvdd.t1301 58.7461
R5880 dvdd.t506 dvdd.t1136 58.7461
R5881 dvdd.t773 dvdd.t1329 58.7461
R5882 dvdd.t332 dvdd.t1495 58.7461
R5883 dvdd.t1191 dvdd 58.7461
R5884 dvdd dvdd.t1144 58.7461
R5885 dvdd.t15 dvdd.t23 58.7461
R5886 dvdd.t14 dvdd.t20 58.7461
R5887 dvdd dvdd.t1124 58.7461
R5888 dvdd.t1167 dvdd.t1615 57.0676
R5889 dvdd dvdd.t582 57.0676
R5890 dvdd.t400 dvdd 57.0676
R5891 dvdd dvdd.t723 57.0676
R5892 dvdd.t1003 dvdd 57.0676
R5893 dvdd.n68 dvdd.t1061 55.9594
R5894 dvdd.n68 dvdd.t1058 55.9594
R5895 dvdd.n2649 dvdd.t899 55.9594
R5896 dvdd.n2649 dvdd.t624 55.9594
R5897 dvdd.n106 dvdd.t1429 55.4067
R5898 dvdd.n1412 dvdd.t1012 55.4067
R5899 dvdd.n1538 dvdd.t730 55.4067
R5900 dvdd.n1542 dvdd.t1383 55.4067
R5901 dvdd.n2123 dvdd.t619 55.4067
R5902 dvdd.n2184 dvdd.t523 55.4067
R5903 dvdd.n2185 dvdd.t1517 55.4067
R5904 dvdd.n2492 dvdd.t1339 55.4067
R5905 dvdd.n2397 dvdd.t661 55.4067
R5906 dvdd.n2465 dvdd.t635 55.4067
R5907 dvdd.n2366 dvdd.t889 55.4067
R5908 dvdd.n2385 dvdd.t1477 55.4067
R5909 dvdd.n2403 dvdd.t575 55.4067
R5910 dvdd.n2564 dvdd.t405 55.4067
R5911 dvdd.t1799 dvdd.t570 55.3892
R5912 dvdd.t486 dvdd.t600 55.3892
R5913 dvdd.t1029 dvdd 55.3892
R5914 dvdd.t403 dvdd.t1037 55.3892
R5915 dvdd.t942 dvdd.t821 53.7107
R5916 dvdd.t861 dvdd 53.7107
R5917 dvdd dvdd.t771 53.7107
R5918 dvdd dvdd.t1426 53.7107
R5919 dvdd.t1462 dvdd 53.7107
R5920 dvdd dvdd.t1217 53.7107
R5921 dvdd.n1504 dvdd.t259 53.1905
R5922 dvdd.t232 dvdd.t791 52.0323
R5923 dvdd dvdd.t598 52.0323
R5924 dvdd.t940 dvdd.t1317 52.0323
R5925 dvdd.t504 dvdd 52.0323
R5926 dvdd.t1255 dvdd 52.0323
R5927 dvdd.t729 dvdd 52.0323
R5928 dvdd dvdd.t1146 52.0323
R5929 dvdd.t258 dvdd.t1089 52.0323
R5930 dvdd dvdd.t396 52.0323
R5931 dvdd dvdd.t1171 52.0323
R5932 dvdd.t616 dvdd 52.0323
R5933 dvdd.t888 dvdd 52.0323
R5934 dvdd dvdd.t1528 52.0323
R5935 dvdd.n143 dvdd.t1899 50.5057
R5936 dvdd.t518 dvdd 50.3539
R5937 dvdd.t769 dvdd 50.3539
R5938 dvdd.t1381 dvdd 50.3539
R5939 dvdd.t658 dvdd 50.3539
R5940 dvdd.t1505 dvdd 50.3539
R5941 dvdd dvdd.t626 50.3539
R5942 dvdd.t1136 dvdd 50.3539
R5943 dvdd.t1047 dvdd.t114 50.3539
R5944 dvdd.t1041 dvdd.t126 50.3539
R5945 dvdd.t1045 dvdd.t112 50.3539
R5946 dvdd dvdd.t78 50.3539
R5947 dvdd.t317 dvdd.t1462 50.3539
R5948 dvdd.t1520 dvdd 50.3539
R5949 dvdd dvdd.t146 50.3539
R5950 dvdd dvdd.t679 50.3539
R5951 dvdd dvdd.t404 50.3539
R5952 dvdd.n2846 dvdd.t302 50.0005
R5953 dvdd.t375 dvdd.t1325 48.6754
R5954 dvdd.t646 dvdd 48.6754
R5955 dvdd dvdd.t1035 48.6754
R5956 dvdd dvdd.t1634 48.6754
R5957 dvdd.t1468 dvdd 48.6754
R5958 dvdd.t1043 dvdd.t128 48.6754
R5959 dvdd.t406 dvdd.t1379 48.6754
R5960 dvdd.t246 dvdd.t142 48.6754
R5961 dvdd.t1637 dvdd 48.6754
R5962 dvdd dvdd.t1740 48.6754
R5963 dvdd.n3087 dvdd.t693 47.2949
R5964 dvdd.n6 dvdd.t184 47.2949
R5965 dvdd.n13 dvdd.t1432 47.2949
R5966 dvdd.n20 dvdd.t1436 47.2949
R5967 dvdd.n27 dvdd.t1419 47.2949
R5968 dvdd.n34 dvdd.t1551 47.2949
R5969 dvdd.n41 dvdd.t1671 47.2949
R5970 dvdd.n48 dvdd.t1680 47.2949
R5971 dvdd.n55 dvdd.t1598 47.2949
R5972 dvdd.n62 dvdd.t1466 47.2949
R5973 dvdd.n2712 dvdd.t1105 47.2949
R5974 dvdd.n2705 dvdd.t1364 47.2949
R5975 dvdd.n2698 dvdd.t1248 47.2949
R5976 dvdd.n2691 dvdd.t1434 47.2949
R5977 dvdd.n2684 dvdd.t1549 47.2949
R5978 dvdd.n2677 dvdd.t1669 47.2949
R5979 dvdd.n2670 dvdd.t1678 47.2949
R5980 dvdd.n2663 dvdd.t1596 47.2949
R5981 dvdd.n2656 dvdd.t890 47.2949
R5982 dvdd dvdd.t901 46.997
R5983 dvdd.t1497 dvdd 46.997
R5984 dvdd.t266 dvdd.t666 46.997
R5985 dvdd dvdd.t985 46.997
R5986 dvdd.t841 dvdd.t1456 46.997
R5987 dvdd.n2965 dvdd.n2964 46.2505
R5988 dvdd.n2963 dvdd.n2946 46.2505
R5989 dvdd.n3147 dvdd.n3146 45.9299
R5990 dvdd.t602 dvdd 45.3185
R5991 dvdd dvdd.t1193 45.3185
R5992 dvdd.t498 dvdd.t338 45.3185
R5993 dvdd.t1034 dvdd.t1575 45.3185
R5994 dvdd.t1493 dvdd 45.3185
R5995 dvdd.t394 dvdd.t1252 45.3185
R5996 dvdd dvdd.t416 45.3185
R5997 dvdd dvdd.t530 45.3185
R5998 dvdd.t381 dvdd.t550 43.6401
R5999 dvdd.t983 dvdd.t1404 43.6401
R6000 dvdd dvdd.t1491 43.6401
R6001 dvdd.t1343 dvdd.t1011 43.6401
R6002 dvdd.t455 dvdd 43.6401
R6003 dvdd dvdd.t418 43.6401
R6004 dvdd.n649 dvdd.t854 43.3874
R6005 dvdd.n977 dvdd.t135 43.3874
R6006 dvdd.n1405 dvdd.t1188 43.3874
R6007 dvdd.n1493 dvdd.t667 43.3874
R6008 dvdd.n1637 dvdd.t1394 43.3874
R6009 dvdd.n1585 dvdd.t864 43.3874
R6010 dvdd.n1989 dvdd.t69 43.3874
R6011 dvdd.n2115 dvdd.t71 43.3874
R6012 dvdd.n477 dvdd.t547 42.3555
R6013 dvdd.n477 dvdd.t384 42.3555
R6014 dvdd.n764 dvdd.t1026 42.3555
R6015 dvdd.n1247 dvdd.t1057 42.3555
R6016 dvdd.t492 dvdd.t524 41.9616
R6017 dvdd.t813 dvdd.t1366 41.9616
R6018 dvdd.t1370 dvdd.t1005 41.9616
R6019 dvdd.t130 dvdd.t319 41.9616
R6020 dvdd.t779 dvdd.t910 41.9616
R6021 dvdd.t162 dvdd.t1122 41.9616
R6022 dvdd.n470 dvdd.t442 41.5552
R6023 dvdd.n470 dvdd.t603 41.5552
R6024 dvdd.n534 dvdd.t373 41.5552
R6025 dvdd.n534 dvdd.t595 41.5552
R6026 dvdd.n746 dvdd.t870 41.5552
R6027 dvdd.n746 dvdd.t601 41.5552
R6028 dvdd.n823 dvdd.t1032 41.5552
R6029 dvdd.n823 dvdd.t597 41.5552
R6030 dvdd.n1040 dvdd.t599 41.5552
R6031 dvdd.n1040 dvdd.t1208 41.5552
R6032 dvdd.n932 dvdd.t1075 41.5552
R6033 dvdd.n932 dvdd.t591 41.5552
R6034 dvdd.n1029 dvdd.t653 41.5552
R6035 dvdd.n1029 dvdd.t593 41.5552
R6036 dvdd.n1110 dvdd.t1234 41.5552
R6037 dvdd.n1110 dvdd.t1414 41.5552
R6038 dvdd.n1228 dvdd.t434 41.5552
R6039 dvdd.n1228 dvdd.t1236 41.5552
R6040 dvdd.n1400 dvdd.t402 41.5552
R6041 dvdd.n1400 dvdd.t424 41.5552
R6042 dvdd.n1408 dvdd.t587 41.5552
R6043 dvdd.n1408 dvdd.t415 41.5552
R6044 dvdd.n1661 dvdd.t1091 41.5552
R6045 dvdd.n1661 dvdd.t421 41.5552
R6046 dvdd.n1690 dvdd.t422 41.5552
R6047 dvdd.n1690 dvdd.t13 41.5552
R6048 dvdd.n1705 dvdd.t22 41.5552
R6049 dvdd.n1705 dvdd.t426 41.5552
R6050 dvdd.n2009 dvdd.t816 41.5552
R6051 dvdd.n2009 dvdd.t417 41.5552
R6052 dvdd.n1905 dvdd.t19 41.5552
R6053 dvdd.n1905 dvdd.t413 41.5552
R6054 dvdd.n1912 dvdd.t1064 41.5552
R6055 dvdd.n1912 dvdd.t419 41.5552
R6056 dvdd.n1795 dvdd.t1084 41.5552
R6057 dvdd.n1795 dvdd.t428 41.5552
R6058 dvdd.n2614 dvdd.t825 41.0422
R6059 dvdd.n2520 dvdd.t893 41.0422
R6060 dvdd.n2516 dvdd.t438 41.0422
R6061 dvdd.n2526 dvdd.t645 41.0422
R6062 dvdd.n2524 dvdd.t937 41.0422
R6063 dvdd.n2365 dvdd.t858 41.0422
R6064 dvdd.n2369 dvdd.t1143 41.0422
R6065 dvdd.n2572 dvdd.t1024 41.0422
R6066 dvdd.n2569 dvdd.t1514 41.0422
R6067 dvdd dvdd.t132 40.2832
R6068 dvdd.t420 dvdd.t264 40.2832
R6069 dvdd dvdd.t742 40.2832
R6070 dvdd.n3116 dvdd.n3115 38.8029
R6071 dvdd.t370 dvdd.t548 38.6047
R6072 dvdd.t346 dvdd.t1156 38.6047
R6073 dvdd.t510 dvdd.t1682 38.6047
R6074 dvdd dvdd.t1207 38.6047
R6075 dvdd dvdd.t1254 38.6047
R6076 dvdd dvdd.t1257 38.6047
R6077 dvdd.t118 dvdd.t1330 38.6047
R6078 dvdd.t1202 dvdd.t843 38.6047
R6079 dvdd.n1685 dvdd.t1501 38.4155
R6080 dvdd.n1334 dvdd.t1044 37.4305
R6081 dvdd.t1789 dvdd.t468 36.9263
R6082 dvdd.t855 dvdd.t1368 36.9263
R6083 dvdd.t640 dvdd.t931 36.9263
R6084 dvdd.t1198 dvdd 36.9263
R6085 dvdd.t391 dvdd.t0 36.9263
R6086 dvdd.t90 dvdd.t262 36.9263
R6087 dvdd.n1046 dvdd.t885 36.4455
R6088 dvdd.n1225 dvdd.t583 36.4455
R6089 dvdd.n2126 dvdd.t1321 36.4455
R6090 dvdd.n1122 dvdd.t1480 36.1587
R6091 dvdd.n1122 dvdd.t1104 36.1587
R6092 dvdd.n2011 dvdd.t1172 36.1587
R6093 dvdd.n2011 dvdd.t531 36.1587
R6094 dvdd.n2181 dvdd.t1348 36.1587
R6095 dvdd.n2181 dvdd.t1028 36.1587
R6096 dvdd.n2580 dvdd.t589 36.1587
R6097 dvdd.n2580 dvdd.t1102 36.1587
R6098 dvdd dvdd.t622 35.2479
R6099 dvdd.t777 dvdd.t321 35.2479
R6100 dvdd dvdd.t642 35.2479
R6101 dvdd.t1504 dvdd 35.2479
R6102 dvdd.t166 dvdd.t1081 35.2479
R6103 dvdd.t1010 dvdd.t799 35.2479
R6104 dvdd.n1135 dvdd.n1134 34.6358
R6105 dvdd.n1283 dvdd.n1282 34.6358
R6106 dvdd.n287 dvdd.n86 34.6358
R6107 dvdd.n288 dvdd.n287 34.6358
R6108 dvdd.n523 dvdd.n352 34.6358
R6109 dvdd.n519 dvdd.n352 34.6358
R6110 dvdd.n519 dvdd.n518 34.6358
R6111 dvdd.n513 dvdd.n512 34.6358
R6112 dvdd.n497 dvdd.n475 34.6358
R6113 dvdd.n597 dvdd.n596 34.6358
R6114 dvdd.n593 dvdd.n592 34.6358
R6115 dvdd.n587 dvdd.n586 34.6358
R6116 dvdd.n793 dvdd.n792 34.6358
R6117 dvdd.n884 dvdd.n815 34.6358
R6118 dvdd.n975 dvdd.n974 34.6358
R6119 dvdd.n998 dvdd.n943 34.6358
R6120 dvdd.n1010 dvdd.n1008 34.6358
R6121 dvdd.n1014 dvdd.n1013 34.6358
R6122 dvdd.n1017 dvdd.n935 34.6358
R6123 dvdd.n1093 dvdd.n1092 34.6358
R6124 dvdd.n1087 dvdd.n1057 34.6358
R6125 dvdd.n1070 dvdd.n1069 34.6358
R6126 dvdd.n1184 dvdd.n1183 34.6358
R6127 dvdd.n1178 dvdd.n1177 34.6358
R6128 dvdd.n1319 dvdd.n1226 34.6358
R6129 dvdd.n1267 dvdd.n1256 34.6358
R6130 dvdd.n1459 dvdd.n1388 34.6358
R6131 dvdd.n1455 dvdd.n1454 34.6358
R6132 dvdd.n1447 dvdd.n1446 34.6358
R6133 dvdd.n1443 dvdd.n1398 34.6358
R6134 dvdd.n1439 dvdd.n1438 34.6358
R6135 dvdd.n1438 dvdd.n1403 34.6358
R6136 dvdd.n1434 dvdd.n1403 34.6358
R6137 dvdd.n1432 dvdd.n1406 34.6358
R6138 dvdd.n1574 dvdd.n1573 34.6358
R6139 dvdd.n1561 dvdd.n1540 34.6358
R6140 dvdd.n1777 dvdd.n1495 34.6358
R6141 dvdd.n1767 dvdd.n1495 34.6358
R6142 dvdd.n1780 dvdd.n1492 34.6358
R6143 dvdd.n1648 dvdd.n1640 34.6358
R6144 dvdd.n1675 dvdd.n1674 34.6358
R6145 dvdd.n1674 dvdd.n1673 34.6358
R6146 dvdd.n1679 dvdd.n1678 34.6358
R6147 dvdd.n1682 dvdd.n1501 34.6358
R6148 dvdd.n1596 dvdd.n1594 34.6358
R6149 dvdd.n1753 dvdd.n1688 34.6358
R6150 dvdd.n1741 dvdd.n1740 34.6358
R6151 dvdd.n1740 dvdd.n1694 34.6358
R6152 dvdd.n1736 dvdd.n1694 34.6358
R6153 dvdd.n1733 dvdd.n1732 34.6358
R6154 dvdd.n1729 dvdd.n1728 34.6358
R6155 dvdd.n1728 dvdd.n1727 34.6358
R6156 dvdd.n1727 dvdd.n1701 34.6358
R6157 dvdd.n1891 dvdd.n1888 34.6358
R6158 dvdd.n1896 dvdd.n1895 34.6358
R6159 dvdd.n1904 dvdd.n1903 34.6358
R6160 dvdd.n1907 dvdd.n1904 34.6358
R6161 dvdd.n1911 dvdd.n1910 34.6358
R6162 dvdd.n2037 dvdd.n2036 34.6358
R6163 dvdd.n2030 dvdd.n2017 34.6358
R6164 dvdd.n2026 dvdd.n2017 34.6358
R6165 dvdd.n2346 dvdd.n2345 34.6358
R6166 dvdd.n2347 dvdd.n2346 34.6358
R6167 dvdd.n2499 dvdd.n2389 34.6358
R6168 dvdd.n2535 dvdd.n2522 34.6358
R6169 dvdd.n2529 dvdd.n2528 34.6358
R6170 dvdd.n2635 dvdd.n2634 34.6358
R6171 dvdd.n2632 dvdd.n2558 34.6358
R6172 dvdd.n2628 dvdd.n2627 34.6358
R6173 dvdd.n2625 dvdd.n2563 34.6358
R6174 dvdd.n2621 dvdd.n2563 34.6358
R6175 dvdd.n2621 dvdd.n2620 34.6358
R6176 dvdd.n482 dvdd.t755 34.4755
R6177 dvdd.n919 dvdd.t1238 34.4755
R6178 dvdd.n1214 dvdd.t1496 34.4755
R6179 dvdd.n1494 dvdd.t267 34.4755
R6180 dvdd.n1494 dvdd.t982 34.4755
R6181 dvdd.n1519 dvdd.n1518 34.3087
R6182 dvdd.n1519 dvdd.n1517 34.3087
R6183 dvdd.n1663 dvdd.n1662 34.3045
R6184 dvdd.n1183 dvdd.n925 34.2593
R6185 dvdd.n1562 dvdd.n1561 34.2593
R6186 dvdd.n106 dvdd.t1473 34.0906
R6187 dvdd.n1412 dvdd.t724 34.0906
R6188 dvdd.n1538 dvdd.t454 34.0906
R6189 dvdd.n1542 dvdd.t1002 34.0906
R6190 dvdd.n2123 dvdd.t1219 34.0906
R6191 dvdd.n2184 dvdd.t1399 34.0906
R6192 dvdd.n2185 dvdd.t1519 34.0906
R6193 dvdd.n2492 dvdd.t1408 34.0906
R6194 dvdd.n2397 dvdd.t655 34.0906
R6195 dvdd.n2465 dvdd.t1216 34.0906
R6196 dvdd.n2366 dvdd.t1131 34.0906
R6197 dvdd.n2385 dvdd.t850 34.0906
R6198 dvdd.n2403 dvdd.t1316 34.0906
R6199 dvdd.n2564 dvdd.t5 34.0906
R6200 dvdd.n588 dvdd.n587 33.8829
R6201 dvdd.n1556 dvdd.n1540 33.8829
R6202 dvdd.n1761 dvdd.n1499 33.8829
R6203 dvdd.n2549 dvdd.n2548 33.8829
R6204 dvdd.n750 dvdd.n745 33.6462
R6205 dvdd.n812 dvdd.n625 33.6462
R6206 dvdd.n1374 dvdd.n1326 33.6462
R6207 dvdd.n1958 dvdd.n1946 33.6462
R6208 dvdd.n1954 dvdd.n1953 33.6462
R6209 dvdd.t727 dvdd 33.5694
R6210 dvdd.t1065 dvdd.t834 33.5694
R6211 dvdd.n788 dvdd.n787 33.5064
R6212 dvdd.n1098 dvdd.n1052 33.5064
R6213 dvdd.n482 dvdd.t804 33.4905
R6214 dvdd.n919 dvdd.t1406 33.4905
R6215 dvdd.n1214 dvdd.t906 33.4905
R6216 dvdd.n71 dvdd.n70 33.4807
R6217 dvdd.n2652 dvdd.n2651 33.4807
R6218 dvdd.n1358 dvdd.n1342 33.2805
R6219 dvdd.n462 dvdd.n461 33.1299
R6220 dvdd.n486 dvdd.n484 33.1299
R6221 dvdd.n1088 dvdd.n1087 33.1299
R6222 dvdd.n1876 dvdd.n1823 33.1299
R6223 dvdd.n2530 dvdd.n2529 33.1299
R6224 dvdd.n605 dvdd.n336 33.1299
R6225 dvdd.n809 dvdd.n808 32.9148
R6226 dvdd.n3084 dvdd.t1205 32.8338
R6227 dvdd.n3084 dvdd.t694 32.8338
R6228 dvdd.n3 dvdd.t920 32.8338
R6229 dvdd.n3 dvdd.t185 32.8338
R6230 dvdd.n10 dvdd.t1232 32.8338
R6231 dvdd.n10 dvdd.t1433 32.8338
R6232 dvdd.n17 dvdd.t1213 32.8338
R6233 dvdd.n17 dvdd.t1437 32.8338
R6234 dvdd.n24 dvdd.t1141 32.8338
R6235 dvdd.n24 dvdd.t1420 32.8338
R6236 dvdd.n31 dvdd.t1251 32.8338
R6237 dvdd.n31 dvdd.t1552 32.8338
R6238 dvdd.n38 dvdd.t1386 32.8338
R6239 dvdd.n38 dvdd.t1672 32.8338
R6240 dvdd.n45 dvdd.t430 32.8338
R6241 dvdd.n45 dvdd.t1681 32.8338
R6242 dvdd.n52 dvdd.t577 32.8338
R6243 dvdd.n52 dvdd.t1599 32.8338
R6244 dvdd.n59 dvdd.t35 32.8338
R6245 dvdd.n59 dvdd.t1467 32.8338
R6246 dvdd.n2716 dvdd.t918 32.8338
R6247 dvdd.n2716 dvdd.t1106 32.8338
R6248 dvdd.n2709 dvdd.t788 32.8338
R6249 dvdd.n2709 dvdd.t1365 32.8338
R6250 dvdd.n2702 dvdd.t1262 32.8338
R6251 dvdd.n2702 dvdd.t1249 32.8338
R6252 dvdd.n2695 dvdd.t1139 32.8338
R6253 dvdd.n2695 dvdd.t1435 32.8338
R6254 dvdd.n2688 dvdd.t411 32.8338
R6255 dvdd.n2688 dvdd.t1550 32.8338
R6256 dvdd.n2681 dvdd.t1484 32.8338
R6257 dvdd.n2681 dvdd.t1670 32.8338
R6258 dvdd.n2674 dvdd.t515 32.8338
R6259 dvdd.n2674 dvdd.t1679 32.8338
R6260 dvdd.n2667 dvdd.t229 32.8338
R6261 dvdd.n2667 dvdd.t1597 32.8338
R6262 dvdd.n2660 dvdd.t95 32.8338
R6263 dvdd.n2660 dvdd.t891 32.8338
R6264 dvdd.n1133 dvdd.n1132 32.7534
R6265 dvdd.n478 dvdd.t1170 32.5055
R6266 dvdd.n478 dvdd.t551 32.5055
R6267 dvdd.n335 dvdd.t1425 32.5055
R6268 dvdd.n335 dvdd.t1273 32.5055
R6269 dvdd.n1066 dvdd.t1260 32.5055
R6270 dvdd.n1066 dvdd.t29 32.5055
R6271 dvdd.n1212 dvdd.t388 32.5055
R6272 dvdd.n1212 dvdd.t609 32.5055
R6273 dvdd.n976 dvdd.n975 32.377
R6274 dvdd.n1021 dvdd.n935 32.377
R6275 dvdd.n1023 dvdd.n1022 32.377
R6276 dvdd.n1446 dvdd.n1445 32.377
R6277 dvdd.n1596 dvdd.n1595 32.377
R6278 dvdd.n1899 dvdd.n1815 32.377
R6279 dvdd.n518 dvdd.n466 32.377
R6280 dvdd.n1466 dvdd.n1465 32.377
R6281 dvdd.n1977 dvdd.n1976 32.377
R6282 dvdd.n1007 dvdd.n940 32.0005
R6283 dvdd.n1566 dvdd.n1539 32.0005
R6284 dvdd.n1554 dvdd.n1553 32.0005
R6285 dvdd.n2332 dvdd.n2331 32.0005
R6286 dvdd.t512 dvdd.t6 31.891
R6287 dvdd.t480 dvdd.t874 31.891
R6288 dvdd.t1237 dvdd 31.891
R6289 dvdd.t1395 dvdd.t116 31.891
R6290 dvdd.t806 dvdd.t1148 31.891
R6291 dvdd.t849 dvdd 31.891
R6292 dvdd.n3102 dvdd.n3100 31.8331
R6293 dvdd.n1373 dvdd.n1372 31.0862
R6294 dvdd.n3089 dvdd.n3086 30.8889
R6295 dvdd.n3086 dvdd.n3085 30.8889
R6296 dvdd.n8 dvdd.n5 30.8889
R6297 dvdd.n5 dvdd.n4 30.8889
R6298 dvdd.n15 dvdd.n12 30.8889
R6299 dvdd.n12 dvdd.n11 30.8889
R6300 dvdd.n22 dvdd.n19 30.8889
R6301 dvdd.n19 dvdd.n18 30.8889
R6302 dvdd.n29 dvdd.n26 30.8889
R6303 dvdd.n26 dvdd.n25 30.8889
R6304 dvdd.n36 dvdd.n33 30.8889
R6305 dvdd.n33 dvdd.n32 30.8889
R6306 dvdd.n43 dvdd.n40 30.8889
R6307 dvdd.n40 dvdd.n39 30.8889
R6308 dvdd.n50 dvdd.n47 30.8889
R6309 dvdd.n47 dvdd.n46 30.8889
R6310 dvdd.n57 dvdd.n54 30.8889
R6311 dvdd.n54 dvdd.n53 30.8889
R6312 dvdd.n64 dvdd.n61 30.8889
R6313 dvdd.n61 dvdd.n60 30.8889
R6314 dvdd.n2714 dvdd.n2711 30.8889
R6315 dvdd.n2711 dvdd.n2710 30.8889
R6316 dvdd.n2707 dvdd.n2704 30.8889
R6317 dvdd.n2704 dvdd.n2703 30.8889
R6318 dvdd.n2700 dvdd.n2697 30.8889
R6319 dvdd.n2697 dvdd.n2696 30.8889
R6320 dvdd.n2693 dvdd.n2690 30.8889
R6321 dvdd.n2690 dvdd.n2689 30.8889
R6322 dvdd.n2686 dvdd.n2683 30.8889
R6323 dvdd.n2683 dvdd.n2682 30.8889
R6324 dvdd.n2679 dvdd.n2676 30.8889
R6325 dvdd.n2676 dvdd.n2675 30.8889
R6326 dvdd.n2672 dvdd.n2669 30.8889
R6327 dvdd.n2669 dvdd.n2668 30.8889
R6328 dvdd.n2665 dvdd.n2662 30.8889
R6329 dvdd.n2662 dvdd.n2661 30.8889
R6330 dvdd.n2658 dvdd.n2655 30.8889
R6331 dvdd.n2655 dvdd.n2654 30.8889
R6332 dvdd.n1434 dvdd.n1433 30.8711
R6333 dvdd.n2342 dvdd.n2341 30.8711
R6334 dvdd.n804 dvdd.n803 30.7205
R6335 dvdd.n1969 dvdd.n1937 30.7205
R6336 dvdd.n84 dvdd.t761 30.5355
R6337 dvdd.n921 dvdd.t1494 30.5355
R6338 dvdd.n1223 dvdd.t763 30.5355
R6339 dvdd.n1254 dvdd.t1108 30.5355
R6340 dvdd.t546 dvdd.t1271 30.2125
R6341 dvdd.t508 dvdd.t904 30.2125
R6342 dvdd.t860 dvdd.t1311 30.2125
R6343 dvdd.t1067 dvdd.t785 30.2125
R6344 dvdd.n903 dvdd.n621 30.1181
R6345 dvdd.n1003 dvdd.n1001 30.1181
R6346 dvdd.n1139 dvdd.n1138 30.1181
R6347 dvdd.n1451 dvdd.n1394 30.1181
R6348 dvdd.n1621 dvdd.n1620 30.1181
R6349 dvdd.n1883 dvdd.n1820 30.1181
R6350 dvdd.n1366 dvdd.n1340 29.9891
R6351 dvdd.n1461 dvdd.n1216 29.7417
R6352 dvdd.n1742 dvdd.n1741 29.7417
R6353 dvdd.n1704 dvdd.n1701 29.7417
R6354 dvdd.n1881 dvdd.n1880 29.7417
R6355 dvdd.n1974 dvdd.n1973 29.7417
R6356 dvdd.n1509 dvdd.t1247 29.5505
R6357 dvdd.n1509 dvdd.t141 29.5505
R6358 dvdd.n3127 dvdd.t1286 29.5505
R6359 dvdd.n785 dvdd.n784 29.3652
R6360 dvdd.n1281 dvdd.n1280 29.3652
R6361 dvdd.n739 dvdd.n738 29.2576
R6362 dvdd.n2081 dvdd.n2080 28.9887
R6363 dvdd.n753 dvdd.t1196 28.752
R6364 dvdd.n1657 dvdd.t1503 28.5655
R6365 dvdd.n1517 dvdd.t1145 28.5655
R6366 dvdd.n2956 dvdd.t559 28.5655
R6367 dvdd.n2956 dvdd.t565 28.5655
R6368 dvdd.n2955 dvdd.t567 28.5655
R6369 dvdd.n2955 dvdd.t563 28.5655
R6370 dvdd.n2954 dvdd.t702 28.5655
R6371 dvdd.n2954 dvdd.t569 28.5655
R6372 dvdd.n2948 dvdd.t714 28.5655
R6373 dvdd.n2948 dvdd.t704 28.5655
R6374 dvdd.n2949 dvdd.t553 28.5655
R6375 dvdd.n2949 dvdd.t1291 28.5655
R6376 dvdd.n2950 dvdd.t557 28.5655
R6377 dvdd.n2950 dvdd.t555 28.5655
R6378 dvdd.n3117 dvdd.t1353 28.5655
R6379 dvdd.n3117 dvdd.t243 28.5655
R6380 dvdd.n3125 dvdd.t1294 28.5655
R6381 dvdd.n3125 dvdd.t1424 28.5655
R6382 dvdd.n3124 dvdd.t1422 28.5655
R6383 dvdd.t1294 dvdd.n3124 28.5655
R6384 dvdd.n3127 dvdd.t239 28.5655
R6385 dvdd.n3129 dvdd.t241 28.5655
R6386 dvdd.n3129 dvdd.t245 28.5655
R6387 dvdd.n3130 dvdd.t237 28.5655
R6388 dvdd.n3130 dvdd.t235 28.5655
R6389 dvdd.n3118 dvdd.t1361 28.5655
R6390 dvdd.n3118 dvdd.t1363 28.5655
R6391 dvdd.n3119 dvdd.t444 28.5655
R6392 dvdd.n3119 dvdd.t448 28.5655
R6393 dvdd.n3097 dvdd.t1355 28.5655
R6394 dvdd.n3097 dvdd.t446 28.5655
R6395 dvdd.n3152 dvdd.t1359 28.5655
R6396 dvdd.n3152 dvdd.t1357 28.5655
R6397 dvdd.t1695 dvdd 28.5341
R6398 dvdd.t474 dvdd 28.5341
R6399 dvdd.t28 dvdd 28.5341
R6400 dvdd.n1826 dvdd 28.5341
R6401 dvdd.t1796 dvdd 28.5341
R6402 dvdd dvdd.t1525 28.5341
R6403 dvdd.n2556 dvdd 28.5341
R6404 dvdd.n2388 dvdd.t1337 28.5169
R6405 dvdd.n2504 dvdd.t633 28.5169
R6406 dvdd.n2514 dvdd.t617 28.5169
R6407 dvdd.n927 dvdd.t377 28.4453
R6408 dvdd.n1533 dvdd.t1380 28.4453
R6409 dvdd.n292 dvdd.n85 28.2358
R6410 dvdd.n1195 dvdd.n1194 28.2358
R6411 dvdd.n1276 dvdd.n1275 28.2358
R6412 dvdd.n1623 dvdd.n1501 28.2358
R6413 dvdd.n2350 dvdd.n2110 27.8593
R6414 dvdd.n70 dvdd.n69 27.7986
R6415 dvdd.n2651 dvdd.n2650 27.7986
R6416 dvdd.n84 dvdd.t539 27.5805
R6417 dvdd.n529 dvdd.t1155 27.5805
R6418 dvdd.n529 dvdd.t1335 27.5805
R6419 dvdd.n531 dvdd.t913 27.5805
R6420 dvdd.n531 dvdd.t665 27.5805
R6421 dvdd.n802 dvdd.t471 27.5805
R6422 dvdd.n802 dvdd.t1461 27.5805
R6423 dvdd.n730 dvdd.t473 27.5805
R6424 dvdd.n730 dvdd.t485 27.5805
R6425 dvdd.n736 dvdd.t495 27.5805
R6426 dvdd.n736 dvdd.t481 27.5805
R6427 dvdd.n631 dvdd.t493 27.5805
R6428 dvdd.n631 dvdd.t479 27.5805
R6429 dvdd.n744 dvdd.t477 27.5805
R6430 dvdd.n747 dvdd.t487 27.5805
R6431 dvdd.n747 dvdd.t501 27.5805
R6432 dvdd.n626 dvdd.t483 27.5805
R6433 dvdd.n626 dvdd.t497 27.5805
R6434 dvdd.n754 dvdd.t475 27.5805
R6435 dvdd.n754 dvdd.t491 27.5805
R6436 dvdd.n757 dvdd.t1453 27.5805
R6437 dvdd.n757 dvdd.t1465 27.5805
R6438 dvdd.n1046 dvdd.t772 27.5805
R6439 dvdd.n921 dvdd.t605 27.5805
R6440 dvdd.n922 dvdd.t631 27.5805
R6441 dvdd.n922 dvdd.t1471 27.5805
R6442 dvdd.n1107 dvdd.t1302 27.5805
R6443 dvdd.n1107 dvdd.t902 27.5805
R6444 dvdd.n1329 dvdd.t107 27.5805
R6445 dvdd.n1329 dvdd.t121 27.5805
R6446 dvdd.n1223 dvdd.t27 27.5805
R6447 dvdd.n1225 dvdd.t1427 27.5805
R6448 dvdd.n1248 dvdd.t1367 27.5805
R6449 dvdd.n1248 dvdd.t1006 27.5805
R6450 dvdd.n1254 dvdd.t509 27.5805
R6451 dvdd.n1378 dvdd.t111 27.5805
R6452 dvdd.n1378 dvdd.t123 27.5805
R6453 dvdd.n1331 dvdd.t103 27.5805
R6454 dvdd.n1331 dvdd.t117 27.5805
R6455 dvdd.n1334 dvdd.t1396 27.5805
R6456 dvdd.n1335 dvdd.t115 27.5805
R6457 dvdd.n1338 dvdd.t1048 27.5805
R6458 dvdd.n1338 dvdd.t1042 27.5805
R6459 dvdd.n1339 dvdd.t127 27.5805
R6460 dvdd.n1339 dvdd.t113 27.5805
R6461 dvdd.n1341 dvdd.t125 27.5805
R6462 dvdd.n1341 dvdd.t133 27.5805
R6463 dvdd.n1344 dvdd.t119 27.5805
R6464 dvdd.n1344 dvdd.t131 27.5805
R6465 dvdd.n1346 dvdd.t105 27.5805
R6466 dvdd.n1346 dvdd.t778 27.5805
R6467 dvdd.n1349 dvdd.t774 27.5805
R6468 dvdd.n1349 dvdd.t780 27.5805
R6469 dvdd.n1555 dvdd.t1308 27.5805
R6470 dvdd.n1555 dvdd.t251 27.5805
R6471 dvdd.n1658 dvdd.t1498 27.5805
R6472 dvdd.n1513 dvdd.t868 27.5805
R6473 dvdd.n1513 dvdd.t253 27.5805
R6474 dvdd.n1518 dvdd.t248 27.5805
R6475 dvdd.n1934 dvdd.t1457 27.5805
R6476 dvdd.n1934 dvdd.t1451 27.5805
R6477 dvdd.n1936 dvdd.t1459 27.5805
R6478 dvdd.n1936 dvdd.t177 27.5805
R6479 dvdd.n1939 dvdd.t151 27.5805
R6480 dvdd.n1939 dvdd.t163 27.5805
R6481 dvdd.n1940 dvdd.t175 27.5805
R6482 dvdd.n1940 dvdd.t159 27.5805
R6483 dvdd.n1944 dvdd.t169 27.5805
R6484 dvdd.n1944 dvdd.t155 27.5805
R6485 dvdd.n1945 dvdd.t167 27.5805
R6486 dvdd.n1948 dvdd.t165 27.5805
R6487 dvdd.n1948 dvdd.t179 27.5805
R6488 dvdd.n1793 dvdd.t161 27.5805
R6489 dvdd.n1793 dvdd.t173 27.5805
R6490 dvdd.n1796 dvdd.t157 27.5805
R6491 dvdd.n1796 dvdd.t171 27.5805
R6492 dvdd.n2126 dvdd.t1397 27.5805
R6493 dvdd.n1351 dvdd.n1347 27.5797
R6494 dvdd.n492 dvdd.n491 27.4829
R6495 dvdd.n597 dvdd.n348 27.4829
R6496 dvdd.n1070 dvdd.n1063 27.4829
R6497 dvdd.n2500 dvdd.n2499 27.4829
R6498 dvdd.n2550 dvdd.n2549 27.4829
R6499 dvdd.n514 dvdd.n513 27.4829
R6500 dvdd.n1746 dvdd.n1691 27.4829
R6501 dvdd.n1722 dvdd.n1721 27.4829
R6502 dvdd.n1910 dvdd.n1813 27.4829
R6503 dvdd.n2112 dvdd.t676 27.3647
R6504 dvdd.n2560 dvdd.t741 27.3647
R6505 dvdd.n2562 dvdd.t732 27.3647
R6506 dvdd.n800 dvdd.n758 27.1064
R6507 dvdd.n1351 dvdd.n1350 27.1064
R6508 dvdd.n276 dvdd.n194 27.0566
R6509 dvdd.n172 dvdd.n171 27.0566
R6510 dvdd.n1844 dvdd.n1842 27.0566
R6511 dvdd.n2422 dvdd.n2421 27.0566
R6512 dvdd.n465 dvdd.t876 26.9729
R6513 dvdd.n1062 dvdd.t1030 26.9729
R6514 dvdd.n1218 dvdd.t1469 26.9729
R6515 dvdd.n1243 dvdd.t627 26.9729
R6516 dvdd.n1330 dvdd.t1264 26.9729
R6517 dvdd.n2505 dvdd.t1214 26.9729
R6518 dvdd.t1276 dvdd.t754 26.8556
R6519 dvdd.t726 dvdd.t374 26.8556
R6520 dvdd.t393 dvdd.t1237 26.8556
R6521 dvdd.t750 dvdd.t1223 26.8556
R6522 dvdd.t1349 dvdd.t1227 26.8556
R6523 dvdd dvdd.t1773 26.8556
R6524 dvdd.n114 dvdd.n113 26.7859
R6525 dvdd.n2202 dvdd.n2201 26.7859
R6526 dvdd.n792 dvdd.n761 26.7299
R6527 dvdd.n743 dvdd.n629 26.6976
R6528 dvdd.n1951 dvdd.n1950 26.6976
R6529 dvdd.n359 dvdd.t465 26.5955
R6530 dvdd.n359 dvdd.t463 26.5955
R6531 dvdd.n479 dvdd.t382 26.5955
R6532 dvdd.n479 dvdd.t1277 26.5955
R6533 dvdd.n338 dvdd.t549 26.5955
R6534 dvdd.n338 dvdd.t1157 26.5955
R6535 dvdd.n744 dvdd.t489 26.5955
R6536 dvdd.n618 dvdd.t1270 26.5955
R6537 dvdd.n618 dvdd.t543 26.5955
R6538 dvdd.n1104 dvdd.t390 26.5955
R6539 dvdd.n1104 dvdd.t988 26.5955
R6540 dvdd.n1335 dvdd.t129 26.5955
R6541 dvdd.n1642 dvdd.t1253 26.5955
R6542 dvdd.n1642 dvdd.t933 26.5955
R6543 dvdd.n1685 dvdd.t261 26.5955
R6544 dvdd.n1945 dvdd.t153 26.5955
R6545 dvdd.n2152 dvdd.t308 26.5955
R6546 dvdd.n2152 dvdd.t307 26.5955
R6547 dvdd.n2105 dvdd.t183 26.5955
R6548 dvdd.n2105 dvdd.t182 26.5955
R6549 dvdd.n2874 dvdd.t706 26.5955
R6550 dvdd.n2874 dvdd.t708 26.5955
R6551 dvdd.n2878 dvdd.t211 26.5955
R6552 dvdd.n2878 dvdd.t205 26.5955
R6553 dvdd.n2879 dvdd.t201 26.5955
R6554 dvdd.n2879 dvdd.t195 26.5955
R6555 dvdd.n2882 dvdd.t203 26.5955
R6556 dvdd.n2882 dvdd.t209 26.5955
R6557 dvdd.n2899 dvdd.t225 26.5955
R6558 dvdd.n2899 dvdd.t207 26.5955
R6559 dvdd.n2885 dvdd.t219 26.5955
R6560 dvdd.n2885 dvdd.t199 26.5955
R6561 dvdd.n2890 dvdd.t197 26.5955
R6562 dvdd.n2890 dvdd.t223 26.5955
R6563 dvdd.n2888 dvdd.t221 26.5955
R6564 dvdd.n2888 dvdd.t217 26.5955
R6565 dvdd.n3028 dvdd.t696 26.5955
R6566 dvdd.n3028 dvdd.t698 26.5955
R6567 dvdd.n3032 dvdd.t974 26.5955
R6568 dvdd.n3032 dvdd.t968 26.5955
R6569 dvdd.n3033 dvdd.t964 26.5955
R6570 dvdd.n3033 dvdd.t958 26.5955
R6571 dvdd.n3036 dvdd.t966 26.5955
R6572 dvdd.n3036 dvdd.t972 26.5955
R6573 dvdd.n3053 dvdd.t956 26.5955
R6574 dvdd.n3053 dvdd.t970 26.5955
R6575 dvdd.n3039 dvdd.t950 26.5955
R6576 dvdd.n3039 dvdd.t962 26.5955
R6577 dvdd.n3044 dvdd.t960 26.5955
R6578 dvdd.n3044 dvdd.t954 26.5955
R6579 dvdd.n3042 dvdd.t952 26.5955
R6580 dvdd.n3042 dvdd.t948 26.5955
R6581 dvdd.n2971 dvdd.t1000 26.5955
R6582 dvdd.n2971 dvdd.t998 26.5955
R6583 dvdd.n2975 dvdd.t67 26.5955
R6584 dvdd.n2975 dvdd.t61 26.5955
R6585 dvdd.n2976 dvdd.t57 26.5955
R6586 dvdd.n2976 dvdd.t51 26.5955
R6587 dvdd.n2979 dvdd.t59 26.5955
R6588 dvdd.n2979 dvdd.t65 26.5955
R6589 dvdd.n2996 dvdd.t49 26.5955
R6590 dvdd.n2996 dvdd.t63 26.5955
R6591 dvdd.n2982 dvdd.t43 26.5955
R6592 dvdd.n2982 dvdd.t55 26.5955
R6593 dvdd.n2987 dvdd.t53 26.5955
R6594 dvdd.n2987 dvdd.t47 26.5955
R6595 dvdd.n2985 dvdd.t45 26.5955
R6596 dvdd.n2985 dvdd.t41 26.5955
R6597 dvdd.n2808 dvdd.t191 26.5955
R6598 dvdd.n2808 dvdd.t189 26.5955
R6599 dvdd.n2804 dvdd.t700 26.5955
R6600 dvdd.n2804 dvdd.t684 26.5955
R6601 dvdd.n2812 dvdd.t303 26.5955
R6602 dvdd.n2812 dvdd.t299 26.5955
R6603 dvdd.n2813 dvdd.t279 26.5955
R6604 dvdd.n2813 dvdd.t275 26.5955
R6605 dvdd.n2816 dvdd.t289 26.5955
R6606 dvdd.n2816 dvdd.t301 26.5955
R6607 dvdd.n2833 dvdd.t285 26.5955
R6608 dvdd.n2833 dvdd.t297 26.5955
R6609 dvdd.n2819 dvdd.t295 26.5955
R6610 dvdd.n2819 dvdd.t273 26.5955
R6611 dvdd.n2824 dvdd.t293 26.5955
R6612 dvdd.n2824 dvdd.t283 26.5955
R6613 dvdd.n2822 dvdd.t287 26.5955
R6614 dvdd.n2822 dvdd.t281 26.5955
R6615 dvdd.n288 dvdd.n85 26.3534
R6616 dvdd.n788 dvdd.n761 26.3534
R6617 dvdd.n1272 dvdd.n1255 26.3534
R6618 dvdd.n2036 dvdd.n2014 26.3534
R6619 dvdd.n2163 dvdd.n2162 26.3341
R6620 dvdd.n197 dvdd.n77 25.977
R6621 dvdd.n493 dvdd.n475 25.977
R6622 dvdd.n772 dvdd.n771 25.977
R6623 dvdd.n984 dvdd.n983 25.977
R6624 dvdd.n1083 dvdd.n1057 25.977
R6625 dvdd.n1172 dvdd.n1171 25.977
R6626 dvdd.n1273 dvdd.n1272 25.977
R6627 dvdd.n1758 dvdd.n1687 25.977
R6628 dvdd.n387 dvdd.n386 25.8177
R6629 dvdd.n2246 dvdd.n2245 25.8177
R6630 dvdd.n763 dvdd.t759 25.6105
R6631 dvdd.n967 dvdd.t1119 25.6105
R6632 dvdd.n1831 dvdd.t1306 25.6105
R6633 dvdd.n2013 dvdd.t800 25.6105
R6634 dvdd.n2016 dvdd.t798 25.6105
R6635 dvdd.n109 dvdd.n87 25.6005
R6636 dvdd.n1424 dvdd.n1413 25.6005
R6637 dvdd.n1567 dvdd.n1566 25.6005
R6638 dvdd.n1553 dvdd.n1552 25.6005
R6639 dvdd.n2031 dvdd.n2030 25.6005
R6640 dvdd.n2197 dvdd.n2196 25.6005
R6641 dvdd.n2500 dvdd.n2386 25.6005
R6642 dvdd.n2495 dvdd.n2490 25.6005
R6643 dvdd.n2640 dvdd.n2639 25.6005
R6644 dvdd.n1653 dvdd.n1652 25.224
R6645 dvdd.n1602 dvdd.n1599 25.1912
R6646 dvdd.n1981 dvdd.n1980 25.1912
R6647 dvdd.n293 dvdd.n292 25.1912
R6648 dvdd.n171 dvdd.n163 25.1912
R6649 dvdd.n784 dvdd.n765 25.1912
R6650 dvdd.n974 dvdd.n952 25.1912
R6651 dvdd.n1144 dvdd.n1143 25.1912
R6652 dvdd.n1615 dvdd.n1510 25.1912
R6653 dvdd.n1592 dvdd.n1523 25.1912
R6654 dvdd.n1917 dvdd.n1811 25.1912
R6655 dvdd.n2331 dvdd.n2121 25.1912
R6656 dvdd.n2612 dvdd.n2567 25.1912
R6657 dvdd.t350 dvdd 25.1772
R6658 dvdd.t170 dvdd 25.1772
R6659 dvdd.n738 dvdd.n737 24.8691
R6660 dvdd.n1950 dvdd.n1794 24.8691
R6661 dvdd.n113 dvdd.n107 24.8476
R6662 dvdd.n906 dvdd.n619 24.8476
R6663 dvdd.n994 dvdd.n991 24.8476
R6664 dvdd.n1079 dvdd.n1061 24.8476
R6665 dvdd.n1290 dvdd.n1289 24.8476
R6666 dvdd.n1617 dvdd.n1616 24.8476
R6667 dvdd.n1873 dvdd.n1824 24.8476
R6668 dvdd.n2201 dvdd.n2186 24.8476
R6669 dvdd.n2620 dvdd.n2565 24.8476
R6670 dvdd.n66 dvdd.t1062 24.6255
R6671 dvdd.n66 dvdd.t1060 24.6255
R6672 dvdd.n2653 dvdd.t900 24.6255
R6673 dvdd.n2653 dvdd.t898 24.6255
R6674 dvdd.n737 dvdd.n632 24.5034
R6675 dvdd.n322 dvdd.n77 24.4711
R6676 dvdd.n983 dvdd.n950 24.4711
R6677 dvdd.n1280 dvdd.n1249 24.4711
R6678 dvdd.n1479 dvdd.n1478 24.4711
R6679 dvdd.n1767 dvdd.n1766 24.4711
R6680 dvdd.n507 dvdd.n471 24.4382
R6681 dvdd.n487 dvdd.n486 24.0946
R6682 dvdd.n1075 dvdd.n1074 24.0946
R6683 dvdd.n1268 dvdd.n1267 24.0946
R6684 dvdd.n1568 dvdd.n1567 24.0946
R6685 dvdd.n1754 dvdd.n1753 24.0946
R6686 dvdd.n2032 dvdd.n2014 24.0946
R6687 dvdd.n2528 dvdd.n2367 24.0946
R6688 dvdd.n2639 dvdd.n2638 24.0946
R6689 dvdd.n2613 dvdd.n2612 24.0946
R6690 dvdd.n1369 dvdd.n1368 23.7719
R6691 dvdd.n1577 dvdd.n1531 23.7181
R6692 dvdd.n2067 dvdd.n1998 23.7181
R6693 dvdd.n280 dvdd.n194 23.7181
R6694 dvdd.n283 dvdd.n86 23.7181
R6695 dvdd.n386 dvdd.n383 23.7181
R6696 dvdd.n1099 dvdd.n1098 23.7181
R6697 dvdd.n1069 dvdd.n1068 23.7181
R6698 dvdd.n1132 dvdd.n1129 23.7181
R6699 dvdd.n1385 dvdd.n1221 23.7181
R6700 dvdd.n1287 dvdd.n1245 23.7181
R6701 dvdd.n1283 dvdd.n1245 23.7181
R6702 dvdd.n1263 dvdd.n1256 23.7181
R6703 dvdd.n1461 dvdd.n1460 23.7181
R6704 dvdd.n1460 dvdd.n1459 23.7181
R6705 dvdd.n1761 dvdd.n1760 23.7181
R6706 dvdd.n1644 dvdd.n1492 23.7181
R6707 dvdd.n1673 dvdd.n1630 23.7181
R6708 dvdd.n1715 dvdd.n1714 23.7181
R6709 dvdd.n1842 dvdd.n1839 23.7181
R6710 dvdd.n2026 dvdd.n2025 23.7181
R6711 dvdd.n2245 dvdd.n2242 23.7181
R6712 dvdd.n2351 dvdd.n2350 23.7181
R6713 dvdd.n2554 dvdd.n2386 23.7181
R6714 dvdd.n2554 dvdd.n2387 23.7181
R6715 dvdd.n2536 dvdd.n2535 23.7181
R6716 dvdd.n2421 dvdd.n2418 23.7181
R6717 dvdd.n2633 dvdd.n2632 23.7181
R6718 dvdd dvdd.t1195 23.4987
R6719 dvdd.t1274 dvdd 23.4987
R6720 dvdd.t352 dvdd 23.4987
R6721 dvdd.t1073 dvdd.t230 23.4987
R6722 dvdd.t385 dvdd.t1259 23.4987
R6723 dvdd dvdd.t1221 23.4987
R6724 dvdd.t122 dvdd.t32 23.4987
R6725 dvdd.t744 dvdd.t1440 23.4987
R6726 dvdd.n460 dvdd.n354 23.3417
R6727 dvdd.n593 dvdd.n349 23.3417
R6728 dvdd.n987 dvdd.n986 23.3417
R6729 dvdd.n1646 dvdd.n1644 23.3417
R6730 dvdd.n1679 dvdd.n1502 23.3417
R6731 dvdd.n3115 dvdd.n3102 23.252
R6732 dvdd.n512 dvdd.n511 22.9652
R6733 dvdd.n601 dvdd.n348 22.9652
R6734 dvdd.n581 dvdd.n532 22.9652
R6735 dvdd.n1028 dvdd.n1027 22.9652
R6736 dvdd.n1045 dvdd.n930 22.9652
R6737 dvdd.n1056 dvdd.n1055 22.9652
R6738 dvdd.n1068 dvdd.n920 22.9652
R6739 dvdd.n1194 dvdd.n923 22.9652
R6740 dvdd.n1165 dvdd.n1164 22.9652
R6741 dvdd.n1428 dvdd.n1406 22.9652
R6742 dvdd.n1652 dvdd.n1640 22.9652
R6743 dvdd.n1593 dvdd.n1592 22.9652
R6744 dvdd.n1749 dvdd.n1748 22.9652
R6745 dvdd.n1719 dvdd.n1706 22.9652
R6746 dvdd.n1913 dvdd.n1911 22.9652
R6747 dvdd.n1160 dvdd.n1159 22.9323
R6748 dvdd.n410 dvdd.n409 22.8981
R6749 dvdd.n1660 dvdd.n1659 22.8837
R6750 dvdd.n804 dvdd.n755 22.6748
R6751 dvdd.n1969 dvdd.n1968 22.6748
R6752 dvdd.n1966 dvdd.n1965 22.6748
R6753 dvdd.n796 dvdd.n758 22.5887
R6754 dvdd.n1074 dvdd.n1063 22.5887
R6755 dvdd.n1173 dvdd.n1172 22.5887
R6756 dvdd.n1288 dvdd.n1287 22.5887
R6757 dvdd.n2032 dvdd.n2031 22.5887
R6758 dvdd.n2550 dvdd.n2387 22.5887
R6759 dvdd.n3091 dvdd 22.5644
R6760 dvdd.n2799 dvdd.n2798 22.5272
R6761 dvdd.n2795 dvdd.n2794 22.5272
R6762 dvdd.n2791 dvdd.n2790 22.5272
R6763 dvdd.n2787 dvdd.n2786 22.5272
R6764 dvdd.n2783 dvdd.n2782 22.5272
R6765 dvdd.n2779 dvdd.n2778 22.5272
R6766 dvdd.n2775 dvdd.n2774 22.5272
R6767 dvdd.n2771 dvdd.n2770 22.5272
R6768 dvdd.n2767 dvdd.n2766 22.5272
R6769 dvdd.n2720 dvdd.n2719 22.5272
R6770 dvdd.n2724 dvdd.n2723 22.5272
R6771 dvdd.n2728 dvdd.n2727 22.5272
R6772 dvdd.n2732 dvdd.n2731 22.5272
R6773 dvdd.n2736 dvdd.n2735 22.5272
R6774 dvdd.n2740 dvdd.n2739 22.5272
R6775 dvdd.n2744 dvdd.n2743 22.5272
R6776 dvdd.n2748 dvdd.n2747 22.5272
R6777 dvdd.n2752 dvdd.n2751 22.5272
R6778 dvdd.n2542 dvdd.n2517 22.4557
R6779 dvdd.n1047 dvdd.n1045 22.2123
R6780 dvdd.n1321 dvdd.n1320 22.2123
R6781 dvdd.n1320 dvdd.n1319 22.2123
R6782 dvdd.n1426 dvdd.n1425 22.2123
R6783 dvdd.n2041 dvdd.n2012 22.2123
R6784 dvdd.n2037 dvdd.n2012 22.2123
R6785 dvdd.n1391 dvdd.n1390 21.8358
R6786 dvdd.t572 dvdd.t875 21.8203
R6787 dvdd.t921 dvdd.t826 21.8203
R6788 dvdd.t516 dvdd.t886 21.8203
R6789 dvdd.t116 dvdd 21.8203
R6790 dvdd.n1387 dvdd.t859 21.8203
R6791 dvdd.n1992 dvdd.t1377 21.8203
R6792 dvdd.n1993 dvdd.t908 21.8203
R6793 dvdd.n586 dvdd.n530 21.4593
R6794 dvdd.n577 dvdd.n576 21.4593
R6795 dvdd.n576 dvdd.n575 21.4593
R6796 dvdd.n772 dvdd.n619 21.4593
R6797 dvdd.n1001 dvdd.n1000 21.4593
R6798 dvdd.n1027 dvdd.n933 21.4593
R6799 dvdd.n1184 dvdd.n923 21.4593
R6800 dvdd.n1164 dvdd.n1111 21.4593
R6801 dvdd.n1316 dvdd.n1226 21.4593
R6802 dvdd.n1478 dvdd.n1209 21.4593
R6803 dvdd.n1467 dvdd.n1466 21.4593
R6804 dvdd.n1428 dvdd.n1427 21.4593
R6805 dvdd.n1663 dvdd.n1660 21.4593
R6806 dvdd.n1616 dvdd.n1615 21.4593
R6807 dvdd.n1594 dvdd.n1593 21.4593
R6808 dvdd.n1749 dvdd.n1688 21.4593
R6809 dvdd.n1715 dvdd.n1706 21.4593
R6810 dvdd.n1876 dvdd.n1875 21.4593
R6811 dvdd.n1913 dvdd.n1811 21.4593
R6812 dvdd.n1977 dvdd.n1933 21.4593
R6813 dvdd.n2042 dvdd.n2041 21.4593
R6814 dvdd.n1759 dvdd.n1758 21.0829
R6815 dvdd.n1168 dvdd.n1105 20.7064
R6816 dvdd.n2162 dvdd.n2150 20.4852
R6817 dvdd.n731 dvdd.n632 20.4805
R6818 dvdd.n1380 dvdd.n1326 20.4805
R6819 dvdd.n1668 dvdd.n1667 20.3532
R6820 dvdd.n602 dvdd.n601 20.3299
R6821 dvdd.n905 dvdd.n904 20.3299
R6822 dvdd.n1003 dvdd.n940 20.3299
R6823 dvdd.n1139 dvdd.n1118 20.3299
R6824 dvdd.n1447 dvdd.n1394 20.3299
R6825 dvdd.n1622 dvdd.n1621 20.3299
R6826 dvdd.n2525 dvdd.n2522 20.3299
R6827 dvdd.n2638 dvdd.n2370 20.3299
R6828 dvdd dvdd.t612 20.1418
R6829 dvdd.t500 dvdd 20.1418
R6830 dvdd.t606 dvdd.t389 20.1418
R6831 dvdd.t1487 dvdd.t987 20.1418
R6832 dvdd.t433 dvdd.t752 20.1418
R6833 dvdd.t110 dvdd.t1255 20.1418
R6834 dvdd.t1327 dvdd.t585 20.1418
R6835 dvdd.n1683 dvdd.t1093 20.1418
R6836 dvdd.t311 dvdd.t74 20.1418
R6837 dvdd.n1372 dvdd.n1371 20.1148
R6838 dvdd.n1371 dvdd.n1370 20.1148
R6839 dvdd.n582 dvdd.n530 19.9534
R6840 dvdd.n993 dvdd.n992 19.9534
R6841 dvdd.n1177 dvdd.n1102 19.9534
R6842 dvdd.n1322 dvdd.n1321 19.9534
R6843 dvdd.n1275 dvdd.n1274 19.9534
R6844 dvdd.n1575 dvdd.n1574 19.9534
R6845 dvdd.n885 dvdd.n884 19.6971
R6846 dvdd.n109 dvdd.n107 19.577
R6847 dvdd.n1082 dvdd.n1081 19.577
R6848 dvdd.n1213 dvdd.n1209 19.577
R6849 dvdd.n1425 dvdd.n1424 19.577
R6850 dvdd.n1570 dvdd.n1569 19.577
R6851 dvdd.n2197 dvdd.n2186 19.577
R6852 dvdd.n2494 dvdd.n2493 19.577
R6853 dvdd.n2634 dvdd.n2633 19.577
R6854 dvdd.n2080 dvdd.n1798 19.2314
R6855 dvdd.n258 dvdd.n257 19.2067
R6856 dvdd.n488 dvdd.n480 19.2005
R6857 dvdd.n1195 dvdd.n920 19.2005
R6858 dvdd.n1291 dvdd.n1290 19.2005
R6859 dvdd.n749 dvdd.n748 19.0176
R6860 dvdd.n2540 dvdd.n2539 18.9384
R6861 dvdd.n2068 dvdd.n2067 18.8301
R6862 dvdd.n488 dvdd.n487 18.824
R6863 dvdd.n1179 dvdd.n1178 18.824
R6864 dvdd.n1573 dvdd.n1534 18.824
R6865 dvdd.n1669 dvdd.n1630 18.824
R6866 dvdd.n2601 dvdd.n2600 18.7912
R6867 dvdd.t1309 dvdd 18.4634
R6868 dvdd.t789 dvdd.t168 18.4634
R6869 dvdd.t148 dvdd 18.4634
R6870 dvdd.n523 dvdd.n351 18.4476
R6871 dvdd.n603 dvdd.n602 18.4476
R6872 dvdd.n589 dvdd.n527 18.4476
R6873 dvdd.n728 dvdd.n727 18.4476
R6874 dvdd.n1013 dvdd.n938 18.4476
R6875 dvdd.n1095 dvdd.n1094 18.4476
R6876 dvdd.n1381 dvdd.n1219 18.4476
R6877 dvdd.n1452 dvdd.n1451 18.4476
R6878 dvdd.n1439 dvdd.n1402 18.4476
R6879 dvdd.n1766 dvdd.n1765 18.4476
R6880 dvdd.n1675 dvdd.n1629 18.4476
R6881 dvdd.n809 dvdd.n627 18.2862
R6882 dvdd.n1362 dvdd.n1361 18.2862
R6883 dvdd.n2830 dvdd.n2820 18.1174
R6884 dvdd.n2835 dvdd.n2832 18.1174
R6885 dvdd.n2839 dvdd.n2817 18.1174
R6886 dvdd.n2842 dvdd.n2841 18.1174
R6887 dvdd.n2850 dvdd.n2849 18.1174
R6888 dvdd.n2854 dvdd.n2853 18.1174
R6889 dvdd.n2858 dvdd.n2857 18.1174
R6890 dvdd.n2859 dvdd.n2858 18.1174
R6891 dvdd.n2864 dvdd.n2862 18.1174
R6892 dvdd.n2868 dvdd.n2805 18.1174
R6893 dvdd.n2869 dvdd.n2868 18.1174
R6894 dvdd.n582 dvdd.n581 18.0711
R6895 dvdd.n801 dvdd.n800 18.0711
R6896 dvdd.n1022 dvdd.n1021 18.0711
R6897 dvdd.n1669 dvdd.n1668 18.0711
R6898 dvdd.n1903 dvdd.n1815 18.0711
R6899 dvdd.n1973 dvdd.n1937 18.0711
R6900 dvdd.n2546 dvdd.n2545 18.0711
R6901 dvdd.n2826 dvdd.n2823 17.9205
R6902 dvdd.n1048 dvdd.n928 17.6946
R6903 dvdd.n1887 dvdd.n1820 17.6946
R6904 dvdd.n301 dvdd.n299 17.612
R6905 dvdd.n134 dvdd.n98 17.612
R6906 dvdd.n682 dvdd.n681 17.612
R6907 dvdd.n1355 dvdd.n1354 17.5548
R6908 dvdd.n3092 dvdd.n3091 17.4938
R6909 dvdd.n2800 dvdd.n2799 17.4938
R6910 dvdd.n2796 dvdd.n2795 17.4938
R6911 dvdd.n2792 dvdd.n2791 17.4938
R6912 dvdd.n2788 dvdd.n2787 17.4938
R6913 dvdd.n2784 dvdd.n2783 17.4938
R6914 dvdd.n2780 dvdd.n2779 17.4938
R6915 dvdd.n2776 dvdd.n2775 17.4938
R6916 dvdd.n2772 dvdd.n2771 17.4938
R6917 dvdd.n2768 dvdd.n2767 17.4938
R6918 dvdd.n2719 dvdd.n2718 17.4938
R6919 dvdd.n2723 dvdd.n2722 17.4938
R6920 dvdd.n2727 dvdd.n2726 17.4938
R6921 dvdd.n2731 dvdd.n2730 17.4938
R6922 dvdd.n2735 dvdd.n2734 17.4938
R6923 dvdd.n2739 dvdd.n2738 17.4938
R6924 dvdd.n2743 dvdd.n2742 17.4938
R6925 dvdd.n2747 dvdd.n2746 17.4938
R6926 dvdd.n2751 dvdd.n2750 17.4938
R6927 dvdd.n238 dvdd.n237 17.3413
R6928 dvdd.n796 dvdd.n795 17.3181
R6929 dvdd.n3155 dvdd.n3154 17.1481
R6930 dvdd.n1427 dvdd.n1426 16.9417
R6931 dvdd.n2859 dvdd.n2806 16.9359
R6932 dvdd.n2870 dvdd.n2869 16.9359
R6933 dvdd.t1750 dvdd.t532 16.785
R6934 dvdd.t1307 dvdd.t1001 16.785
R6935 dvdd.t1389 dvdd.t830 16.785
R6936 dvdd.t1092 dvdd.t98 16.785
R6937 dvdd.t1481 dvdd.t979 16.785
R6938 dvdd.n1315 dvdd.n1314 16.6212
R6939 dvdd.n795 dvdd.n794 16.5652
R6940 dvdd.n1385 dvdd.n1219 16.5652
R6941 dvdd.n3116 dvdd.n3100 16.3333
R6942 dvdd.n456 dvdd.n354 16.2447
R6943 dvdd.n463 dvdd.n351 16.1887
R6944 dvdd.n592 dvdd.n527 16.1887
R6945 dvdd.n1094 dvdd.n1093 16.1887
R6946 dvdd.n1734 dvdd.n1733 16.1887
R6947 dvdd.n1732 dvdd.n1698 16.1887
R6948 dvdd.n2640 dvdd.n2367 16.1887
R6949 dvdd.n2063 dvdd.n1998 16.139
R6950 dvdd.n2468 dvdd.n2464 16.139
R6951 dvdd.n2896 dvdd.n2886 16.132
R6952 dvdd.n2901 dvdd.n2898 16.132
R6953 dvdd.n2905 dvdd.n2883 16.132
R6954 dvdd.n2916 dvdd.n2915 16.132
R6955 dvdd.n2921 dvdd.n2919 16.132
R6956 dvdd.n2925 dvdd.n2875 16.132
R6957 dvdd.n2926 dvdd.n2925 16.132
R6958 dvdd.n1356 dvdd.n1355 16.0919
R6959 dvdd.n2892 dvdd.n2889 15.9567
R6960 dvdd.n3050 dvdd.n3040 15.914
R6961 dvdd.n3055 dvdd.n3052 15.914
R6962 dvdd.n3059 dvdd.n3037 15.914
R6963 dvdd.n3070 dvdd.n3069 15.914
R6964 dvdd.n3075 dvdd.n3073 15.914
R6965 dvdd.n3079 dvdd.n3029 15.914
R6966 dvdd.n3080 dvdd.n3079 15.914
R6967 dvdd.n2993 dvdd.n2983 15.914
R6968 dvdd.n2998 dvdd.n2995 15.914
R6969 dvdd.n3002 dvdd.n2980 15.914
R6970 dvdd.n3013 dvdd.n3012 15.914
R6971 dvdd.n3018 dvdd.n3016 15.914
R6972 dvdd.n3022 dvdd.n2972 15.914
R6973 dvdd.n3023 dvdd.n3022 15.914
R6974 dvdd.n322 dvdd.n321 15.8683
R6975 dvdd.n192 dvdd.n191 15.8683
R6976 dvdd.n2318 dvdd.n2124 15.8683
R6977 dvdd.n1180 dvdd.n1179 15.8123
R6978 dvdd.n1570 dvdd.n1534 15.8123
R6979 dvdd.n2600 dvdd.n2599 15.7794
R6980 dvdd.n2857 dvdd.n2809 15.7543
R6981 dvdd.n2863 dvdd.n2805 15.7543
R6982 dvdd.n3046 dvdd.n3043 15.741
R6983 dvdd.n2989 dvdd.n2986 15.741
R6984 dvdd.n745 dvdd.n743 15.7262
R6985 dvdd.n1954 dvdd.n1946 15.7262
R6986 dvdd.n1662 dvdd.n1635 15.6103
R6987 dvdd.n2914 dvdd.n2913 15.606
R6988 dvdd.n2845 dvdd.n2814 15.5574
R6989 dvdd.n2763 dvdd.n2762 15.5123
R6990 dvdd.n2756 dvdd.n2755 15.5123
R6991 dvdd.n1445 dvdd.n1444 15.4358
R6992 dvdd.n1402 dvdd.n1401 15.4358
R6993 dvdd.n1754 dvdd.n1687 15.4358
R6994 dvdd.n3068 dvdd.n3067 15.3951
R6995 dvdd.n3011 dvdd.n3010 15.3951
R6996 dvdd.n812 dvdd.n627 15.3605
R6997 dvdd.n1363 dvdd.n1362 15.3605
R6998 dvdd.n150 dvdd.n149 15.3162
R6999 dvdd.n2826 dvdd.n2825 15.1636
R7000 dvdd.n2850 dvdd.n2810 15.1636
R7001 dvdd.t766 dvdd.t470 15.1065
R7002 dvdd.t1025 dvdd.t758 15.1065
R7003 dvdd.t457 dvdd.t1209 15.1065
R7004 dvdd.t453 dvdd.t100 15.1065
R7005 dvdd.t18 dvdd.t1007 15.1065
R7006 dvdd dvdd.t1142 15.1065
R7007 dvdd.n2927 dvdd.n2926 15.08
R7008 dvdd.n978 dvdd.n950 15.0593
R7009 dvdd.n1168 dvdd.n1167 15.0593
R7010 dvdd.n1569 dvdd.n1568 15.0593
R7011 dvdd.n1653 dvdd.n1638 14.9121
R7012 dvdd.n2910 dvdd.n2909 14.9046
R7013 dvdd.n575 dvdd.n574 14.9
R7014 dvdd.n864 dvdd.n863 14.9
R7015 dvdd.n3064 dvdd.n3063 14.8762
R7016 dvdd.n3081 dvdd.n3080 14.8762
R7017 dvdd.n3007 dvdd.n3006 14.8762
R7018 dvdd.n3024 dvdd.n3023 14.8762
R7019 dvdd.n1174 dvdd.n1102 14.6829
R7020 dvdd.n1268 dvdd.n1255 14.6829
R7021 dvdd.n1778 dvdd.n1777 14.6829
R7022 dvdd.n1629 dvdd.n1626 14.6829
R7023 dvdd.n2547 dvdd.n2546 14.6829
R7024 dvdd.n2334 dvdd.n2333 14.65
R7025 dvdd.n407 dvdd.n406 14.5851
R7026 dvdd.n555 dvdd.n554 14.5851
R7027 dvdd.n844 dvdd.n843 14.5851
R7028 dvdd.n2267 dvdd.n2144 14.5851
R7029 dvdd.n1289 dvdd.n1288 14.3064
R7030 dvdd.n2531 dvdd.n2525 14.3064
R7031 dvdd.n280 dvdd.n195 14.2735
R7032 dvdd.n208 dvdd.n197 14.2735
R7033 dvdd.n192 dvdd.n88 14.2735
R7034 dvdd.n664 dvdd.n663 14.2735
R7035 dvdd.n776 dvdd.n771 14.2735
R7036 dvdd.n963 dvdd.n960 14.2735
R7037 dvdd.n1991 dvdd.n1808 14.2735
R7038 dvdd.n2321 dvdd.n2124 14.2735
R7039 dvdd.n2589 dvdd.n2588 14.2735
R7040 dvdd.n2909 dvdd.n2908 14.2313
R7041 dvdd.n3145 dvdd.n3144 14.2313
R7042 dvdd.n3142 dvdd.n3138 14.2313
R7043 dvdd.n2920 dvdd.n2875 14.0279
R7044 dvdd.n2615 dvdd.n2613 13.9837
R7045 dvdd.n1433 dvdd.n1432 13.9299
R7046 dvdd.n748 dvdd.n625 13.8976
R7047 dvdd.n2913 dvdd.n2880 13.8526
R7048 dvdd.n3074 dvdd.n3029 13.8383
R7049 dvdd.n3017 dvdd.n2972 13.8383
R7050 dvdd.n3063 dvdd.n3062 13.7042
R7051 dvdd.n3006 dvdd.n3005 13.7042
R7052 dvdd.n3067 dvdd.n3034 13.6654
R7053 dvdd.n3010 dvdd.n2977 13.6654
R7054 dvdd.n1274 dvdd.n1273 13.5534
R7055 dvdd.n2379 dvdd.n2370 13.5534
R7056 dvdd.n2892 dvdd.n2891 13.5019
R7057 dvdd.n2916 dvdd.n2876 13.5019
R7058 dvdd.t441 dvdd.t1159 13.4281
R7059 dvdd.t490 dvdd.t534 13.4281
R7060 dvdd.t1071 dvdd.t1269 13.4281
R7061 dvdd.t520 dvdd.t717 13.4281
R7062 dvdd.t845 dvdd.t915 13.4281
R7063 dvdd.n1101 dvdd.t88 13.4281
R7064 dvdd.t1254 dvdd.t1402 13.4281
R7065 dvdd dvdd.t863 13.4281
R7066 dvdd.t249 dvdd.t1053 13.4281
R7067 dvdd.t1083 dvdd.t172 13.4281
R7068 dvdd.t1733 dvdd.t818 13.4281
R7069 dvdd.t1449 dvdd.t740 13.4281
R7070 dvdd.t731 dvdd.t675 13.4281
R7071 dvdd.t2 dvdd.t1515 13.4281
R7072 dvdd.n3046 dvdd.n3045 13.3194
R7073 dvdd.n3070 dvdd.n3030 13.3194
R7074 dvdd.n2989 dvdd.n2988 13.3194
R7075 dvdd.n3013 dvdd.n2973 13.3194
R7076 dvdd.n283 dvdd.n87 13.177
R7077 dvdd.n906 dvdd.n905 13.177
R7078 dvdd.n994 dvdd.n993 13.177
R7079 dvdd.n1099 dvdd.n928 13.177
R7080 dvdd.n1322 dvdd.n1221 13.177
R7081 dvdd.n1479 dvdd.n1208 13.177
R7082 dvdd.n1468 dvdd.n1467 13.177
R7083 dvdd.n1454 dvdd.n1453 13.177
R7084 dvdd.n1420 dvdd.n1413 13.177
R7085 dvdd.n1552 dvdd.n1551 13.177
R7086 dvdd.n1647 dvdd.n1646 13.177
R7087 dvdd.n1760 dvdd.n1759 13.177
R7088 dvdd.n2196 dvdd.n2195 13.177
R7089 dvdd.n2490 dvdd.n2489 13.177
R7090 dvdd.n1357 dvdd.n1356 13.1662
R7091 dvdd.n2082 dvdd.n1794 13.1662
R7092 dvdd.n2489 dvdd.n2391 12.9693
R7093 dvdd.n1868 dvdd.n1825 12.9273
R7094 dvdd.n987 dvdd.n945 12.8005
R7095 dvdd.n985 dvdd.n984 12.8005
R7096 dvdd.n1869 dvdd.n1868 12.8005
R7097 dvdd.n1869 dvdd.n1824 12.8005
R7098 dvdd.n1875 dvdd.n1874 12.8005
R7099 dvdd.n2352 dvdd.n2351 12.8005
R7100 dvdd.n2548 dvdd.n2547 12.8005
R7101 dvdd.n1292 dvdd.n1291 12.7507
R7102 dvdd.n2758 dvdd.n2757 12.5617
R7103 dvdd.n2166 dvdd.n2165 12.4487
R7104 dvdd.n1576 dvdd.n1575 12.424
R7105 dvdd.n2495 dvdd.n2494 12.424
R7106 dvdd.n2841 dvdd.n2840 12.4067
R7107 dvdd dvdd.n0 12.3787
R7108 dvdd.n3102 dvdd.n3101 12.2424
R7109 dvdd.n2760 dvdd.n2759 12.1783
R7110 dvdd.n3154 dvdd.n3153 12.1678
R7111 dvdd.n1167 dvdd.n1166 12.0476
R7112 dvdd.n1933 dvdd.n1931 12.0476
R7113 dvdd.n2831 dvdd.n2830 12.0128
R7114 dvdd.n2848 dvdd.n2847 12.0128
R7115 dvdd.t664 dvdd.t372 11.7496
R7116 dvdd.t651 dvdd.t781 11.7496
R7117 dvdd.t1111 dvdd.t1384 11.7496
R7118 dvdd.t106 dvdd.t756 11.7496
R7119 dvdd.t226 dvdd.t1200 11.7496
R7120 dvdd.t152 dvdd.t1121 11.7496
R7121 dvdd.t857 dvdd.t888 11.7496
R7122 dvdd.t673 dvdd.t1130 11.7496
R7123 dvdd.n2536 dvdd.n2521 11.7249
R7124 dvdd.n511 dvdd.n510 11.6711
R7125 dvdd.n596 dvdd.n349 11.2946
R7126 dvdd.n1010 dvdd.n1009 11.2946
R7127 dvdd.n1089 dvdd.n1056 11.2946
R7128 dvdd.n1390 dvdd.n1388 11.2946
R7129 dvdd.n1779 dvdd.n1778 11.2946
R7130 dvdd.n1682 dvdd.n1502 11.2946
R7131 dvdd.n1736 dvdd.n1735 11.2946
R7132 dvdd.n1729 dvdd.n1700 11.2946
R7133 dvdd.n2847 dvdd.n2846 11.2126
R7134 dvdd.n3095 dvdd.n3094 11.1517
R7135 dvdd.n2907 dvdd.n2906 11.0471
R7136 dvdd.n807 dvdd.n755 10.9719
R7137 dvdd.n1968 dvdd.n1967 10.9719
R7138 dvdd.n1967 dvdd.n1966 10.9719
R7139 dvdd.n3061 dvdd.n3060 10.8978
R7140 dvdd.n3004 dvdd.n3003 10.8978
R7141 dvdd.n893 dvdd.n621 10.8853
R7142 dvdd.n2897 dvdd.n2896 10.6964
R7143 dvdd.n2010 dvdd.n2008 10.6672
R7144 dvdd.n3051 dvdd.n3050 10.5519
R7145 dvdd.n2994 dvdd.n2993 10.5519
R7146 dvdd.n991 dvdd.n945 10.5417
R7147 dvdd.n1623 dvdd.n1622 10.5417
R7148 dvdd.n2871 dvdd.n2870 10.482
R7149 dvdd.n2928 dvdd.n2927 10.3526
R7150 dvdd.n3082 dvdd.n3081 10.3383
R7151 dvdd.n3025 dvdd.n3024 10.3383
R7152 dvdd.n1959 dvdd.n1958 10.2405
R7153 dvdd.n2616 dvdd.n2565 10.1652
R7154 dvdd.t1323 dvdd.n524 10.0712
R7155 dvdd.t725 dvdd.t594 10.0712
R7156 dvdd.t494 dvdd.t871 10.0712
R7157 dvdd dvdd.t1319 10.0712
R7158 dvdd.t366 dvdd 10.0712
R7159 dvdd.t1189 dvdd.t1187 10.0712
R7160 dvdd.t1509 dvdd.t1087 10.0712
R7161 dvdd.t1511 dvdd.t180 10.0712
R7162 dvdd.t427 dvdd.t156 10.0712
R7163 dvdd.t1444 dvdd.t1338 10.0712
R7164 dvdd.n2765 dvdd.n2764 10.0534
R7165 dvdd.n2754 dvdd.n2753 10.0534
R7166 dvdd.n1033 dvdd.n1030 10.0005
R7167 dvdd.n1042 dvdd.n1041 10.0005
R7168 dvdd.n577 dvdd.n532 9.78874
R7169 dvdd.n1083 dvdd.n1082 9.78874
R7170 dvdd.n1143 dvdd.n1118 9.78874
R7171 dvdd.n2872 dvdd.n2802 9.76224
R7172 dvdd dvdd.t325 9.73577
R7173 dvdd.n254 dvdd.n253 9.73273
R7174 dvdd.n253 dvdd.n252 9.73273
R7175 dvdd.n249 dvdd.n248 9.73273
R7176 dvdd.n248 dvdd.n247 9.73273
R7177 dvdd.n247 dvdd.n227 9.73273
R7178 dvdd.n243 dvdd.n227 9.73273
R7179 dvdd.n243 dvdd.n242 9.73273
R7180 dvdd.n242 dvdd.n241 9.73273
R7181 dvdd.n274 dvdd.n273 9.73273
R7182 dvdd.n273 dvdd.n217 9.73273
R7183 dvdd.n269 dvdd.n268 9.73273
R7184 dvdd.n268 dvdd.n267 9.73273
R7185 dvdd.n267 dvdd.n220 9.73273
R7186 dvdd.n263 dvdd.n220 9.73273
R7187 dvdd.n263 dvdd.n262 9.73273
R7188 dvdd.n262 dvdd.n261 9.73273
R7189 dvdd.n305 dvdd.n82 9.73273
R7190 dvdd.n306 dvdd.n305 9.73273
R7191 dvdd.n308 dvdd.n80 9.73273
R7192 dvdd.n312 dvdd.n80 9.73273
R7193 dvdd.n313 dvdd.n312 9.73273
R7194 dvdd.n314 dvdd.n313 9.73273
R7195 dvdd.n314 dvdd.n78 9.73273
R7196 dvdd.n318 dvdd.n78 9.73273
R7197 dvdd.n130 dvdd.n129 9.73273
R7198 dvdd.n129 dvdd.n128 9.73273
R7199 dvdd.n125 dvdd.n124 9.73273
R7200 dvdd.n124 dvdd.n123 9.73273
R7201 dvdd.n123 dvdd.n103 9.73273
R7202 dvdd.n119 dvdd.n103 9.73273
R7203 dvdd.n119 dvdd.n118 9.73273
R7204 dvdd.n118 dvdd.n117 9.73273
R7205 dvdd.n176 dvdd.n175 9.73273
R7206 dvdd.n177 dvdd.n176 9.73273
R7207 dvdd.n181 dvdd.n180 9.73273
R7208 dvdd.n182 dvdd.n181 9.73273
R7209 dvdd.n182 dvdd.n158 9.73273
R7210 dvdd.n186 dvdd.n158 9.73273
R7211 dvdd.n187 dvdd.n186 9.73273
R7212 dvdd.n188 dvdd.n187 9.73273
R7213 dvdd.n445 dvdd.n444 9.73273
R7214 dvdd.n452 dvdd.n357 9.73273
R7215 dvdd.n714 dvdd.n641 9.73273
R7216 dvdd.n717 dvdd.n716 9.73273
R7217 dvdd.n721 dvdd.n720 9.73273
R7218 dvdd.n722 dvdd.n721 9.73273
R7219 dvdd.n686 dvdd.n685 9.73273
R7220 dvdd.n693 dvdd.n647 9.73273
R7221 dvdd.n878 dvdd.n877 9.73273
R7222 dvdd.n877 dvdd.n819 9.73273
R7223 dvdd.n871 dvdd.n870 9.73273
R7224 dvdd.n870 dvdd.n822 9.73273
R7225 dvdd.n1296 dvdd.n1295 9.73273
R7226 dvdd.n1298 dvdd.n1296 9.73273
R7227 dvdd.n1302 dvdd.n1301 9.73273
R7228 dvdd.n1304 dvdd.n1231 9.73273
R7229 dvdd.n1308 dvdd.n1231 9.73273
R7230 dvdd.n1309 dvdd.n1308 9.73273
R7231 dvdd.n1311 dvdd.n1309 9.73273
R7232 dvdd.n1848 dvdd.n1832 9.73273
R7233 dvdd.n1852 dvdd.n1829 9.73273
R7234 dvdd.n1856 dvdd.n1829 9.73273
R7235 dvdd.n2059 dvdd.n2000 9.73273
R7236 dvdd.n2055 dvdd.n2054 9.73273
R7237 dvdd.n2054 dvdd.n2053 9.73273
R7238 dvdd.n2053 dvdd.n2005 9.73273
R7239 dvdd.n2049 dvdd.n2005 9.73273
R7240 dvdd.n2047 dvdd.n2046 9.73273
R7241 dvdd.n2316 dvdd.n2315 9.73273
R7242 dvdd.n2269 dvdd.n2143 9.73273
R7243 dvdd.n2273 dvdd.n2143 9.73273
R7244 dvdd.n2206 dvdd.n2182 9.73273
R7245 dvdd.n2481 dvdd.n2398 9.73273
R7246 dvdd.n2485 dvdd.n2483 9.73273
R7247 dvdd.n2472 dvdd.n2400 9.73273
R7248 dvdd.n2453 dvdd.n2404 9.73273
R7249 dvdd.n2456 dvdd.n2455 9.73273
R7250 dvdd.n164 dvdd 9.6274
R7251 dvdd.n233 dvdd.n231 9.60526
R7252 dvdd.n737 dvdd.n735 9.56172
R7253 dvdd.n745 dvdd.n628 9.56172
R7254 dvdd.n866 dvdd.n824 9.52116
R7255 dvdd.n461 dvdd.n460 9.41227
R7256 dvdd.n1008 dvdd.n1007 9.41227
R7257 dvdd.n1350 dvdd.n1208 9.41227
R7258 dvdd.n1444 dvdd.n1443 9.41227
R7259 dvdd.n1888 dvdd.n1887 9.41227
R7260 dvdd.n1895 dvdd.n1817 9.41227
R7261 dvdd.n2342 dvdd.n2113 9.41227
R7262 dvdd.n2561 dvdd.n2558 9.41227
R7263 dvdd.n2626 dvdd.n2625 9.41227
R7264 dvdd.n168 dvdd.n167 9.3005
R7265 dvdd.n169 dvdd.n163 9.3005
R7266 dvdd.n171 dvdd.n170 9.3005
R7267 dvdd.n173 dvdd.n172 9.3005
R7268 dvdd.n175 dvdd.n174 9.3005
R7269 dvdd.n176 dvdd.n161 9.3005
R7270 dvdd.n178 dvdd.n177 9.3005
R7271 dvdd.n180 dvdd.n179 9.3005
R7272 dvdd.n181 dvdd.n159 9.3005
R7273 dvdd.n183 dvdd.n182 9.3005
R7274 dvdd.n184 dvdd.n158 9.3005
R7275 dvdd.n186 dvdd.n185 9.3005
R7276 dvdd.n187 dvdd.n157 9.3005
R7277 dvdd.n189 dvdd.n188 9.3005
R7278 dvdd.n191 dvdd.n190 9.3005
R7279 dvdd.n192 dvdd.n155 9.3005
R7280 dvdd.n154 dvdd.n88 9.3005
R7281 dvdd.n153 dvdd.n152 9.3005
R7282 dvdd.n150 dvdd.n89 9.3005
R7283 dvdd.n149 dvdd.n148 9.3005
R7284 dvdd.n147 dvdd.n146 9.3005
R7285 dvdd.n95 dvdd.n93 9.3005
R7286 dvdd.n141 dvdd.n140 9.3005
R7287 dvdd.n139 dvdd.n96 9.3005
R7288 dvdd.n138 dvdd.n137 9.3005
R7289 dvdd.n136 dvdd.n97 9.3005
R7290 dvdd.n134 dvdd.n133 9.3005
R7291 dvdd.n132 dvdd.n98 9.3005
R7292 dvdd.n131 dvdd.n130 9.3005
R7293 dvdd.n129 dvdd.n99 9.3005
R7294 dvdd.n128 dvdd.n127 9.3005
R7295 dvdd.n126 dvdd.n125 9.3005
R7296 dvdd.n124 dvdd.n102 9.3005
R7297 dvdd.n123 dvdd.n122 9.3005
R7298 dvdd.n121 dvdd.n103 9.3005
R7299 dvdd.n120 dvdd.n119 9.3005
R7300 dvdd.n118 dvdd.n104 9.3005
R7301 dvdd.n117 dvdd.n116 9.3005
R7302 dvdd.n115 dvdd.n114 9.3005
R7303 dvdd.n113 dvdd.n112 9.3005
R7304 dvdd.n111 dvdd.n107 9.3005
R7305 dvdd.n110 dvdd.n109 9.3005
R7306 dvdd.n108 dvdd.n87 9.3005
R7307 dvdd.n284 dvdd.n283 9.3005
R7308 dvdd.n285 dvdd.n86 9.3005
R7309 dvdd.n287 dvdd.n286 9.3005
R7310 dvdd.n289 dvdd.n288 9.3005
R7311 dvdd.n290 dvdd.n85 9.3005
R7312 dvdd.n292 dvdd.n291 9.3005
R7313 dvdd.n293 dvdd 9.3005
R7314 dvdd.n297 dvdd.n296 9.3005
R7315 dvdd.n299 dvdd.n298 9.3005
R7316 dvdd.n302 dvdd.n301 9.3005
R7317 dvdd.n303 dvdd.n82 9.3005
R7318 dvdd.n305 dvdd.n304 9.3005
R7319 dvdd.n306 dvdd.n81 9.3005
R7320 dvdd.n309 dvdd.n308 9.3005
R7321 dvdd.n310 dvdd.n80 9.3005
R7322 dvdd.n312 dvdd.n311 9.3005
R7323 dvdd.n313 dvdd.n79 9.3005
R7324 dvdd.n315 dvdd.n314 9.3005
R7325 dvdd.n316 dvdd.n78 9.3005
R7326 dvdd.n318 dvdd.n317 9.3005
R7327 dvdd.n321 dvdd.n320 9.3005
R7328 dvdd.n323 dvdd.n322 9.3005
R7329 dvdd.n198 dvdd.n77 9.3005
R7330 dvdd.n206 dvdd.n197 9.3005
R7331 dvdd.n208 dvdd.n207 9.3005
R7332 dvdd.n211 dvdd.n196 9.3005
R7333 dvdd.n214 dvdd.n213 9.3005
R7334 dvdd.n215 dvdd.n195 9.3005
R7335 dvdd.n280 dvdd.n279 9.3005
R7336 dvdd.n278 dvdd.n194 9.3005
R7337 dvdd.n277 dvdd.n276 9.3005
R7338 dvdd.n274 dvdd.n216 9.3005
R7339 dvdd.n273 dvdd.n272 9.3005
R7340 dvdd.n271 dvdd.n217 9.3005
R7341 dvdd.n270 dvdd.n269 9.3005
R7342 dvdd.n268 dvdd.n218 9.3005
R7343 dvdd.n267 dvdd.n266 9.3005
R7344 dvdd.n265 dvdd.n220 9.3005
R7345 dvdd.n264 dvdd.n263 9.3005
R7346 dvdd.n262 dvdd.n221 9.3005
R7347 dvdd.n261 dvdd.n260 9.3005
R7348 dvdd.n259 dvdd.n258 9.3005
R7349 dvdd.n257 dvdd.n256 9.3005
R7350 dvdd.n255 dvdd.n254 9.3005
R7351 dvdd.n253 dvdd.n224 9.3005
R7352 dvdd.n252 dvdd.n251 9.3005
R7353 dvdd.n250 dvdd.n249 9.3005
R7354 dvdd.n248 dvdd.n226 9.3005
R7355 dvdd.n247 dvdd.n246 9.3005
R7356 dvdd.n245 dvdd.n227 9.3005
R7357 dvdd.n244 dvdd.n243 9.3005
R7358 dvdd.n242 dvdd.n228 9.3005
R7359 dvdd.n241 dvdd.n240 9.3005
R7360 dvdd.n239 dvdd.n238 9.3005
R7361 dvdd.n237 dvdd.n236 9.3005
R7362 dvdd.n235 dvdd.n234 9.3005
R7363 dvdd.n386 dvdd.n385 9.3005
R7364 dvdd.n388 dvdd.n387 9.3005
R7365 dvdd.n390 dvdd.n389 9.3005
R7366 dvdd.n391 dvdd.n375 9.3005
R7367 dvdd.n393 dvdd.n392 9.3005
R7368 dvdd.n395 dvdd.n394 9.3005
R7369 dvdd.n396 dvdd.n373 9.3005
R7370 dvdd.n398 dvdd.n397 9.3005
R7371 dvdd.n399 dvdd.n372 9.3005
R7372 dvdd.n401 dvdd.n400 9.3005
R7373 dvdd.n402 dvdd.n371 9.3005
R7374 dvdd.n404 dvdd.n403 9.3005
R7375 dvdd.n406 dvdd.n405 9.3005
R7376 dvdd.n412 dvdd.n411 9.3005
R7377 dvdd.n414 dvdd.n413 9.3005
R7378 dvdd.n415 dvdd.n368 9.3005
R7379 dvdd.n419 dvdd.n418 9.3005
R7380 dvdd.n420 dvdd.n367 9.3005
R7381 dvdd.n422 dvdd.n421 9.3005
R7382 dvdd.n424 dvdd.n366 9.3005
R7383 dvdd.n426 dvdd.n425 9.3005
R7384 dvdd.n427 dvdd.n365 9.3005
R7385 dvdd.n429 dvdd.n428 9.3005
R7386 dvdd.n430 dvdd.n364 9.3005
R7387 dvdd.n434 dvdd.n433 9.3005
R7388 dvdd.n437 dvdd.n436 9.3005
R7389 dvdd.n439 dvdd.n361 9.3005
R7390 dvdd.n442 dvdd.n441 9.3005
R7391 dvdd.n444 dvdd.n443 9.3005
R7392 dvdd.n445 dvdd.n358 9.3005
R7393 dvdd.n449 dvdd.n448 9.3005
R7394 dvdd.n450 dvdd.n357 9.3005
R7395 dvdd.n452 dvdd.n451 9.3005
R7396 dvdd.n454 dvdd.n355 9.3005
R7397 dvdd.n457 dvdd.n456 9.3005
R7398 dvdd.n458 dvdd.n354 9.3005
R7399 dvdd.n460 dvdd.n459 9.3005
R7400 dvdd.n461 dvdd.n353 9.3005
R7401 dvdd.n464 dvdd.n463 9.3005
R7402 dvdd.n523 dvdd.n522 9.3005
R7403 dvdd.n521 dvdd.n352 9.3005
R7404 dvdd.n520 dvdd.n519 9.3005
R7405 dvdd.n518 dvdd.n517 9.3005
R7406 dvdd.n516 dvdd.n515 9.3005
R7407 dvdd.n513 dvdd.n467 9.3005
R7408 dvdd.n512 dvdd.n468 9.3005
R7409 dvdd.n510 dvdd.n509 9.3005
R7410 dvdd.n508 dvdd.n507 9.3005
R7411 dvdd.n504 dvdd.n503 9.3005
R7412 dvdd.n502 dvdd.n501 9.3005
R7413 dvdd.n499 dvdd.n473 9.3005
R7414 dvdd.n497 dvdd.n496 9.3005
R7415 dvdd.n495 dvdd.n475 9.3005
R7416 dvdd.n494 dvdd.n493 9.3005
R7417 dvdd.n492 dvdd.n476 9.3005
R7418 dvdd.n491 dvdd.n490 9.3005
R7419 dvdd.n489 dvdd.n488 9.3005
R7420 dvdd.n487 dvdd.n481 9.3005
R7421 dvdd.n486 dvdd.n485 9.3005
R7422 dvdd.n483 dvdd.n333 9.3005
R7423 dvdd.n606 dvdd.n605 9.3005
R7424 dvdd.n603 dvdd.n337 9.3005
R7425 dvdd.n602 dvdd.n347 9.3005
R7426 dvdd.n601 dvdd.n600 9.3005
R7427 dvdd.n599 dvdd.n348 9.3005
R7428 dvdd.n598 dvdd.n597 9.3005
R7429 dvdd.n596 dvdd.n595 9.3005
R7430 dvdd.n594 dvdd.n593 9.3005
R7431 dvdd.n592 dvdd.n591 9.3005
R7432 dvdd.n590 dvdd.n589 9.3005
R7433 dvdd.n587 dvdd.n528 9.3005
R7434 dvdd.n586 dvdd.n585 9.3005
R7435 dvdd.n584 dvdd.n530 9.3005
R7436 dvdd.n583 dvdd.n582 9.3005
R7437 dvdd.n581 dvdd.n580 9.3005
R7438 dvdd.n579 dvdd.n532 9.3005
R7439 dvdd.n578 dvdd.n577 9.3005
R7440 dvdd.n576 dvdd.n533 9.3005
R7441 dvdd.n575 dvdd.n538 9.3005
R7442 dvdd.n574 dvdd.n573 9.3005
R7443 dvdd.n572 dvdd.n571 9.3005
R7444 dvdd.n570 dvdd.n541 9.3005
R7445 dvdd.n569 dvdd.n568 9.3005
R7446 dvdd.n567 dvdd.n566 9.3005
R7447 dvdd.n565 dvdd.n543 9.3005
R7448 dvdd.n564 dvdd.n563 9.3005
R7449 dvdd.n562 dvdd.n544 9.3005
R7450 dvdd.n561 dvdd.n560 9.3005
R7451 dvdd.n559 dvdd.n545 9.3005
R7452 dvdd.n558 dvdd.n557 9.3005
R7453 dvdd.n556 dvdd.n555 9.3005
R7454 dvdd.n665 dvdd.n664 9.3005
R7455 dvdd.n667 dvdd.n666 9.3005
R7456 dvdd.n669 dvdd.n653 9.3005
R7457 dvdd.n672 dvdd.n671 9.3005
R7458 dvdd.n673 dvdd.n652 9.3005
R7459 dvdd.n675 dvdd.n674 9.3005
R7460 dvdd.n679 dvdd.n678 9.3005
R7461 dvdd.n681 dvdd.n680 9.3005
R7462 dvdd.n683 dvdd.n682 9.3005
R7463 dvdd.n685 dvdd.n684 9.3005
R7464 dvdd.n686 dvdd.n648 9.3005
R7465 dvdd.n690 dvdd.n689 9.3005
R7466 dvdd.n691 dvdd.n647 9.3005
R7467 dvdd.n693 dvdd.n692 9.3005
R7468 dvdd.n696 dvdd.n695 9.3005
R7469 dvdd.n698 dvdd.n697 9.3005
R7470 dvdd.n699 dvdd.n644 9.3005
R7471 dvdd.n702 dvdd.n701 9.3005
R7472 dvdd.n706 dvdd.n642 9.3005
R7473 dvdd.n711 dvdd.n710 9.3005
R7474 dvdd.n712 dvdd.n641 9.3005
R7475 dvdd.n714 dvdd.n713 9.3005
R7476 dvdd.n716 dvdd.n640 9.3005
R7477 dvdd.n718 dvdd.n717 9.3005
R7478 dvdd.n720 dvdd.n719 9.3005
R7479 dvdd.n721 dvdd.n637 9.3005
R7480 dvdd.n723 dvdd.n722 9.3005
R7481 dvdd.n725 dvdd.n724 9.3005
R7482 dvdd.n727 dvdd.n635 9.3005
R7483 dvdd.n728 dvdd.n633 9.3005
R7484 dvdd.n733 dvdd.n732 9.3005
R7485 dvdd.n734 dvdd.n632 9.3005
R7486 dvdd.n738 dvdd.n630 9.3005
R7487 dvdd.n741 dvdd.n740 9.3005
R7488 dvdd.n743 dvdd.n742 9.3005
R7489 dvdd.n751 dvdd.n750 9.3005
R7490 dvdd.n752 dvdd.n625 9.3005
R7491 dvdd.n812 dvdd.n811 9.3005
R7492 dvdd.n810 dvdd.n809 9.3005
R7493 dvdd.n807 dvdd.n806 9.3005
R7494 dvdd.n805 dvdd.n804 9.3005
R7495 dvdd.n801 dvdd.n756 9.3005
R7496 dvdd.n800 dvdd.n799 9.3005
R7497 dvdd.n798 dvdd.n758 9.3005
R7498 dvdd.n797 dvdd.n796 9.3005
R7499 dvdd.n793 dvdd.n759 9.3005
R7500 dvdd.n792 dvdd.n791 9.3005
R7501 dvdd.n790 dvdd.n761 9.3005
R7502 dvdd.n789 dvdd.n788 9.3005
R7503 dvdd.n786 dvdd.n762 9.3005
R7504 dvdd.n784 dvdd.n783 9.3005
R7505 dvdd.n782 dvdd.n765 9.3005
R7506 dvdd.n781 dvdd.n780 9.3005
R7507 dvdd.n779 dvdd.n766 9.3005
R7508 dvdd.n776 dvdd.n775 9.3005
R7509 dvdd.n774 dvdd.n771 9.3005
R7510 dvdd.n773 dvdd.n772 9.3005
R7511 dvdd.n619 dvdd.n616 9.3005
R7512 dvdd.n907 dvdd.n906 9.3005
R7513 dvdd.n903 dvdd.n902 9.3005
R7514 dvdd.n895 dvdd.n621 9.3005
R7515 dvdd.n894 dvdd.n893 9.3005
R7516 dvdd.n890 dvdd.n623 9.3005
R7517 dvdd.n889 dvdd.n888 9.3005
R7518 dvdd.n887 dvdd.n886 9.3005
R7519 dvdd.n884 dvdd.n883 9.3005
R7520 dvdd.n882 dvdd.n815 9.3005
R7521 dvdd.n881 dvdd.n880 9.3005
R7522 dvdd.n878 dvdd.n816 9.3005
R7523 dvdd.n877 dvdd.n876 9.3005
R7524 dvdd.n875 dvdd.n819 9.3005
R7525 dvdd.n874 dvdd.n873 9.3005
R7526 dvdd.n871 dvdd.n820 9.3005
R7527 dvdd.n870 dvdd.n869 9.3005
R7528 dvdd.n868 dvdd.n822 9.3005
R7529 dvdd.n867 dvdd.n866 9.3005
R7530 dvdd.n863 dvdd.n862 9.3005
R7531 dvdd.n861 dvdd.n860 9.3005
R7532 dvdd.n859 dvdd.n830 9.3005
R7533 dvdd.n858 dvdd.n857 9.3005
R7534 dvdd.n856 dvdd.n855 9.3005
R7535 dvdd.n854 dvdd.n832 9.3005
R7536 dvdd.n853 dvdd.n852 9.3005
R7537 dvdd.n851 dvdd.n833 9.3005
R7538 dvdd.n850 dvdd.n849 9.3005
R7539 dvdd.n848 dvdd.n834 9.3005
R7540 dvdd.n847 dvdd.n846 9.3005
R7541 dvdd.n845 dvdd.n844 9.3005
R7542 dvdd.n963 dvdd.n962 9.3005
R7543 dvdd.n966 dvdd.n953 9.3005
R7544 dvdd.n971 dvdd.n970 9.3005
R7545 dvdd.n972 dvdd.n952 9.3005
R7546 dvdd.n974 dvdd.n973 9.3005
R7547 dvdd.n975 dvdd.n951 9.3005
R7548 dvdd.n980 dvdd.n979 9.3005
R7549 dvdd.n981 dvdd.n950 9.3005
R7550 dvdd.n983 dvdd.n982 9.3005
R7551 dvdd.n984 dvdd.n949 9.3005
R7552 dvdd.n985 dvdd.n948 9.3005
R7553 dvdd.n986 dvdd.n946 9.3005
R7554 dvdd.n988 dvdd.n987 9.3005
R7555 dvdd.n989 dvdd.n945 9.3005
R7556 dvdd.n991 dvdd.n990 9.3005
R7557 dvdd.n995 dvdd.n994 9.3005
R7558 dvdd.n996 dvdd.n943 9.3005
R7559 dvdd.n998 dvdd.n997 9.3005
R7560 dvdd.n1001 dvdd.n941 9.3005
R7561 dvdd.n1004 dvdd.n1003 9.3005
R7562 dvdd.n1005 dvdd.n940 9.3005
R7563 dvdd.n1007 dvdd.n1006 9.3005
R7564 dvdd.n1008 dvdd.n939 9.3005
R7565 dvdd.n1011 dvdd.n1010 9.3005
R7566 dvdd.n1013 dvdd.n1012 9.3005
R7567 dvdd.n1014 dvdd.n936 9.3005
R7568 dvdd.n1018 dvdd.n1017 9.3005
R7569 dvdd.n1019 dvdd.n935 9.3005
R7570 dvdd.n1021 dvdd.n1020 9.3005
R7571 dvdd.n1022 dvdd.n934 9.3005
R7572 dvdd.n1024 dvdd.n1023 9.3005
R7573 dvdd.n1025 dvdd.n933 9.3005
R7574 dvdd.n1027 dvdd.n1026 9.3005
R7575 dvdd.n1035 dvdd.n1034 9.3005
R7576 dvdd.n1036 dvdd.n931 9.3005
R7577 dvdd.n1038 dvdd.n1037 9.3005
R7578 dvdd.n1044 dvdd.n1043 9.3005
R7579 dvdd.n1045 dvdd 9.3005
R7580 dvdd.n1047 dvdd.n929 9.3005
R7581 dvdd.n1049 dvdd.n1048 9.3005
R7582 dvdd.n1050 dvdd.n928 9.3005
R7583 dvdd.n1099 dvdd.n1051 9.3005
R7584 dvdd.n1098 dvdd.n1097 9.3005
R7585 dvdd.n1096 dvdd.n1095 9.3005
R7586 dvdd.n1093 dvdd.n1053 9.3005
R7587 dvdd.n1092 dvdd.n1091 9.3005
R7588 dvdd.n1090 dvdd.n1089 9.3005
R7589 dvdd.n1087 dvdd.n1086 9.3005
R7590 dvdd.n1085 dvdd.n1057 9.3005
R7591 dvdd.n1084 dvdd.n1083 9.3005
R7592 dvdd.n1082 dvdd.n1058 9.3005
R7593 dvdd.n1081 dvdd.n1060 9.3005
R7594 dvdd.n1079 dvdd.n1078 9.3005
R7595 dvdd.n1077 dvdd.n1061 9.3005
R7596 dvdd.n1076 dvdd.n1075 9.3005
R7597 dvdd.n1074 dvdd.n1073 9.3005
R7598 dvdd.n1072 dvdd.n1063 9.3005
R7599 dvdd.n1071 dvdd.n1070 9.3005
R7600 dvdd.n1068 dvdd.n1067 9.3005
R7601 dvdd.n920 dvdd.n917 9.3005
R7602 dvdd.n1196 dvdd.n1195 9.3005
R7603 dvdd.n1194 dvdd.n1193 9.3005
R7604 dvdd.n1186 dvdd.n923 9.3005
R7605 dvdd.n1185 dvdd.n1184 9.3005
R7606 dvdd.n1183 dvdd.n1182 9.3005
R7607 dvdd.n1181 dvdd.n1180 9.3005
R7608 dvdd.n1178 dvdd.n926 9.3005
R7609 dvdd.n1177 dvdd.n1176 9.3005
R7610 dvdd.n1175 dvdd.n1174 9.3005
R7611 dvdd.n1172 dvdd.n1103 9.3005
R7612 dvdd.n1171 dvdd.n1170 9.3005
R7613 dvdd.n1169 dvdd.n1168 9.3005
R7614 dvdd.n1167 dvdd.n1106 9.3005
R7615 dvdd.n1166 dvdd.n1108 9.3005
R7616 dvdd.n1165 dvdd.n1109 9.3005
R7617 dvdd.n1164 dvdd.n1163 9.3005
R7618 dvdd.n1162 dvdd.n1111 9.3005
R7619 dvdd.n1161 dvdd.n1160 9.3005
R7620 dvdd.n1159 dvdd.n1158 9.3005
R7621 dvdd.n1157 dvdd.n1156 9.3005
R7622 dvdd.n1154 dvdd.n1113 9.3005
R7623 dvdd.n1153 dvdd.n1152 9.3005
R7624 dvdd.n1151 dvdd.n1150 9.3005
R7625 dvdd.n1149 dvdd.n1116 9.3005
R7626 dvdd.n1147 dvdd.n1146 9.3005
R7627 dvdd.n1145 dvdd.n1144 9.3005
R7628 dvdd.n1143 dvdd.n1142 9.3005
R7629 dvdd.n1141 dvdd.n1118 9.3005
R7630 dvdd.n1140 dvdd.n1139 9.3005
R7631 dvdd.n1138 dvdd.n1137 9.3005
R7632 dvdd.n1136 dvdd.n1135 9.3005
R7633 dvdd.n1134 dvdd.n1121 9.3005
R7634 dvdd.n1132 dvdd.n1131 9.3005
R7635 dvdd.n1265 dvdd.n1256 9.3005
R7636 dvdd.n1267 dvdd.n1266 9.3005
R7637 dvdd.n1269 dvdd.n1268 9.3005
R7638 dvdd.n1270 dvdd.n1255 9.3005
R7639 dvdd.n1272 dvdd.n1271 9.3005
R7640 dvdd.n1273 dvdd.n1253 9.3005
R7641 dvdd.n1274 dvdd.n1252 9.3005
R7642 dvdd.n1275 dvdd.n1250 9.3005
R7643 dvdd.n1277 dvdd.n1276 9.3005
R7644 dvdd.n1278 dvdd.n1249 9.3005
R7645 dvdd.n1280 dvdd.n1279 9.3005
R7646 dvdd.n1282 dvdd.n1246 9.3005
R7647 dvdd.n1284 dvdd.n1283 9.3005
R7648 dvdd.n1285 dvdd.n1245 9.3005
R7649 dvdd.n1287 dvdd.n1286 9.3005
R7650 dvdd.n1288 dvdd.n1242 9.3005
R7651 dvdd.n1289 dvdd.n1241 9.3005
R7652 dvdd.n1291 dvdd.n1238 9.3005
R7653 dvdd.n1293 dvdd.n1292 9.3005
R7654 dvdd.n1295 dvdd.n1294 9.3005
R7655 dvdd.n1296 dvdd.n1235 9.3005
R7656 dvdd.n1299 dvdd.n1298 9.3005
R7657 dvdd.n1301 dvdd.n1300 9.3005
R7658 dvdd.n1302 dvdd.n1232 9.3005
R7659 dvdd.n1305 dvdd.n1304 9.3005
R7660 dvdd.n1306 dvdd.n1231 9.3005
R7661 dvdd.n1308 dvdd.n1307 9.3005
R7662 dvdd.n1309 dvdd.n1230 9.3005
R7663 dvdd.n1312 dvdd.n1311 9.3005
R7664 dvdd.n1314 dvdd.n1313 9.3005
R7665 dvdd.n1315 dvdd.n1227 9.3005
R7666 dvdd.n1317 dvdd.n1316 9.3005
R7667 dvdd.n1318 dvdd.n1226 9.3005
R7668 dvdd.n1319 dvdd 9.3005
R7669 dvdd.n1320 dvdd.n1224 9.3005
R7670 dvdd.n1321 dvdd.n1222 9.3005
R7671 dvdd.n1323 dvdd.n1322 9.3005
R7672 dvdd.n1324 dvdd.n1221 9.3005
R7673 dvdd.n1325 dvdd.n1221 9.3005
R7674 dvdd.n1385 dvdd.n1384 9.3005
R7675 dvdd.n1383 dvdd.n1219 9.3005
R7676 dvdd.n1382 dvdd.n1381 9.3005
R7677 dvdd.n1380 dvdd.n1379 9.3005
R7678 dvdd.n1380 dvdd.n1377 9.3005
R7679 dvdd.n1376 dvdd.n1326 9.3005
R7680 dvdd.n1375 dvdd.n1374 9.3005
R7681 dvdd.n1372 dvdd.n1328 9.3005
R7682 dvdd.n1371 dvdd.n1332 9.3005
R7683 dvdd.n1370 dvdd.n1333 9.3005
R7684 dvdd.n1369 dvdd.n1336 9.3005
R7685 dvdd.n1368 dvdd.n1337 9.3005
R7686 dvdd.n1366 dvdd.n1365 9.3005
R7687 dvdd.n1364 dvdd.n1363 9.3005
R7688 dvdd.n1361 dvdd.n1360 9.3005
R7689 dvdd.n1359 dvdd.n1358 9.3005
R7690 dvdd.n1356 dvdd.n1343 9.3005
R7691 dvdd.n1354 dvdd.n1353 9.3005
R7692 dvdd.n1352 dvdd.n1351 9.3005
R7693 dvdd.n1350 dvdd.n1348 9.3005
R7694 dvdd.n1208 dvdd.n1206 9.3005
R7695 dvdd.n1480 dvdd.n1479 9.3005
R7696 dvdd.n1478 dvdd.n1477 9.3005
R7697 dvdd.n1470 dvdd.n1209 9.3005
R7698 dvdd.n1469 dvdd.n1468 9.3005
R7699 dvdd.n1466 dvdd.n1211 9.3005
R7700 dvdd.n1464 dvdd.n1463 9.3005
R7701 dvdd.n1462 dvdd.n1461 9.3005
R7702 dvdd.n1460 dvdd.n1217 9.3005
R7703 dvdd.n1459 dvdd.n1458 9.3005
R7704 dvdd.n1457 dvdd.n1388 9.3005
R7705 dvdd.n1456 dvdd.n1455 9.3005
R7706 dvdd.n1454 dvdd.n1389 9.3005
R7707 dvdd.n1451 dvdd.n1450 9.3005
R7708 dvdd.n1449 dvdd.n1394 9.3005
R7709 dvdd.n1448 dvdd.n1447 9.3005
R7710 dvdd.n1446 dvdd.n1395 9.3005
R7711 dvdd.n1445 dvdd.n1396 9.3005
R7712 dvdd.n1444 dvdd.n1397 9.3005
R7713 dvdd.n1443 dvdd.n1442 9.3005
R7714 dvdd.n1441 dvdd.n1398 9.3005
R7715 dvdd.n1440 dvdd.n1439 9.3005
R7716 dvdd.n1438 dvdd.n1437 9.3005
R7717 dvdd.n1436 dvdd.n1403 9.3005
R7718 dvdd.n1435 dvdd.n1434 9.3005
R7719 dvdd.n1433 dvdd.n1404 9.3005
R7720 dvdd.n1432 dvdd.n1431 9.3005
R7721 dvdd.n1430 dvdd.n1406 9.3005
R7722 dvdd.n1429 dvdd.n1428 9.3005
R7723 dvdd.n1427 dvdd.n1407 9.3005
R7724 dvdd.n1426 dvdd.n1410 9.3005
R7725 dvdd.n1425 dvdd.n1411 9.3005
R7726 dvdd.n1424 dvdd.n1423 9.3005
R7727 dvdd.n1422 dvdd.n1413 9.3005
R7728 dvdd.n1552 dvdd.n1543 9.3005
R7729 dvdd.n1553 dvdd.n1541 9.3005
R7730 dvdd.n1558 dvdd.n1557 9.3005
R7731 dvdd.n1559 dvdd.n1540 9.3005
R7732 dvdd.n1561 dvdd.n1560 9.3005
R7733 dvdd.n1564 dvdd.n1563 9.3005
R7734 dvdd.n1566 dvdd.n1565 9.3005
R7735 dvdd.n1567 dvdd.n1537 9.3005
R7736 dvdd.n1568 dvdd.n1535 9.3005
R7737 dvdd.n1571 dvdd.n1570 9.3005
R7738 dvdd.n1573 dvdd.n1572 9.3005
R7739 dvdd.n1574 dvdd.n1532 9.3005
R7740 dvdd.n1578 dvdd.n1577 9.3005
R7741 dvdd.n1579 dvdd.n1531 9.3005
R7742 dvdd.n1580 dvdd.n1531 9.3005
R7743 dvdd.n1583 dvdd.n1582 9.3005
R7744 dvdd.n1584 dvdd.n1524 9.3005
R7745 dvdd.n1589 dvdd.n1588 9.3005
R7746 dvdd.n1590 dvdd.n1523 9.3005
R7747 dvdd.n1592 dvdd.n1591 9.3005
R7748 dvdd.n1593 dvdd.n1522 9.3005
R7749 dvdd.n1593 dvdd.n1521 9.3005
R7750 dvdd.n1594 dvdd.n1515 9.3005
R7751 dvdd.n1597 dvdd.n1596 9.3005
R7752 dvdd.n1599 dvdd.n1598 9.3005
R7753 dvdd.n1603 dvdd.n1602 9.3005
R7754 dvdd.n1604 dvdd.n1512 9.3005
R7755 dvdd.n1606 dvdd.n1605 9.3005
R7756 dvdd.n1607 dvdd.n1511 9.3005
R7757 dvdd.n1612 dvdd.n1611 9.3005
R7758 dvdd.n1613 dvdd.n1510 9.3005
R7759 dvdd.n1615 dvdd.n1614 9.3005
R7760 dvdd.n1616 dvdd.n1508 9.3005
R7761 dvdd.n1618 dvdd.n1617 9.3005
R7762 dvdd.n1620 dvdd.n1619 9.3005
R7763 dvdd.n1621 dvdd.n1505 9.3005
R7764 dvdd.n1622 dvdd.n1503 9.3005
R7765 dvdd.n1624 dvdd.n1623 9.3005
R7766 dvdd.n1625 dvdd.n1501 9.3005
R7767 dvdd.n1682 dvdd.n1681 9.3005
R7768 dvdd.n1680 dvdd.n1679 9.3005
R7769 dvdd.n1678 dvdd.n1677 9.3005
R7770 dvdd.n1676 dvdd.n1675 9.3005
R7771 dvdd.n1674 dvdd.n1627 9.3005
R7772 dvdd.n1673 dvdd.n1672 9.3005
R7773 dvdd.n1671 dvdd.n1630 9.3005
R7774 dvdd.n1670 dvdd.n1669 9.3005
R7775 dvdd.n1668 dvdd.n1631 9.3005
R7776 dvdd.n1667 dvdd.n1666 9.3005
R7777 dvdd.n1665 dvdd.n1664 9.3005
R7778 dvdd.n1660 dvdd.n1634 9.3005
R7779 dvdd.n1639 dvdd.n1636 9.3005
R7780 dvdd.n1656 dvdd.n1655 9.3005
R7781 dvdd.n1654 dvdd.n1653 9.3005
R7782 dvdd.n1652 dvdd.n1651 9.3005
R7783 dvdd.n1650 dvdd.n1640 9.3005
R7784 dvdd.n1649 dvdd.n1648 9.3005
R7785 dvdd.n1646 dvdd.n1641 9.3005
R7786 dvdd.n1644 dvdd.n1643 9.3005
R7787 dvdd.n1492 dvdd.n1490 9.3005
R7788 dvdd.n1781 dvdd.n1780 9.3005
R7789 dvdd.n1777 dvdd.n1776 9.3005
R7790 dvdd.n1769 dvdd.n1495 9.3005
R7791 dvdd.n1768 dvdd.n1767 9.3005
R7792 dvdd.n1766 dvdd.n1497 9.3005
R7793 dvdd.n1764 dvdd.n1763 9.3005
R7794 dvdd.n1762 dvdd.n1761 9.3005
R7795 dvdd.n1760 dvdd.n1500 9.3005
R7796 dvdd.n1759 dvdd.n1686 9.3005
R7797 dvdd.n1758 dvdd.n1757 9.3005
R7798 dvdd.n1756 dvdd.n1687 9.3005
R7799 dvdd.n1755 dvdd.n1754 9.3005
R7800 dvdd.n1753 dvdd.n1752 9.3005
R7801 dvdd.n1751 dvdd.n1688 9.3005
R7802 dvdd.n1750 dvdd.n1749 9.3005
R7803 dvdd.n1748 dvdd.n1689 9.3005
R7804 dvdd.n1746 dvdd.n1745 9.3005
R7805 dvdd.n1744 dvdd.n1743 9.3005
R7806 dvdd.n1741 dvdd.n1692 9.3005
R7807 dvdd.n1740 dvdd.n1739 9.3005
R7808 dvdd.n1738 dvdd.n1694 9.3005
R7809 dvdd.n1737 dvdd.n1736 9.3005
R7810 dvdd.n1733 dvdd.n1695 9.3005
R7811 dvdd.n1732 dvdd.n1731 9.3005
R7812 dvdd.n1730 dvdd.n1729 9.3005
R7813 dvdd.n1728 dvdd.n1699 9.3005
R7814 dvdd.n1727 dvdd.n1726 9.3005
R7815 dvdd.n1725 dvdd.n1701 9.3005
R7816 dvdd.n1724 dvdd.n1723 9.3005
R7817 dvdd.n1721 dvdd.n1702 9.3005
R7818 dvdd.n1719 dvdd.n1718 9.3005
R7819 dvdd.n1717 dvdd.n1706 9.3005
R7820 dvdd.n1716 dvdd.n1715 9.3005
R7821 dvdd.n1842 dvdd.n1841 9.3005
R7822 dvdd.n1845 dvdd.n1844 9.3005
R7823 dvdd.n1846 dvdd.n1832 9.3005
R7824 dvdd.n1848 dvdd.n1847 9.3005
R7825 dvdd.n1850 dvdd.n1830 9.3005
R7826 dvdd.n1853 dvdd.n1852 9.3005
R7827 dvdd.n1854 dvdd.n1829 9.3005
R7828 dvdd.n1856 dvdd.n1855 9.3005
R7829 dvdd.n1859 dvdd.n1858 9.3005
R7830 dvdd.n1860 dvdd.n1828 9.3005
R7831 dvdd.n1862 dvdd.n1861 9.3005
R7832 dvdd.n1863 dvdd.n1827 9.3005
R7833 dvdd.n1866 dvdd.n1865 9.3005
R7834 dvdd.n1868 dvdd.n1867 9.3005
R7835 dvdd.n1870 dvdd.n1869 9.3005
R7836 dvdd.n1871 dvdd.n1824 9.3005
R7837 dvdd.n1873 dvdd.n1872 9.3005
R7838 dvdd.n1877 dvdd.n1876 9.3005
R7839 dvdd.n1879 dvdd.n1878 9.3005
R7840 dvdd.n1881 dvdd.n1821 9.3005
R7841 dvdd.n1884 dvdd.n1883 9.3005
R7842 dvdd.n1885 dvdd.n1820 9.3005
R7843 dvdd.n1887 dvdd.n1886 9.3005
R7844 dvdd.n1888 dvdd.n1818 9.3005
R7845 dvdd.n1892 dvdd.n1891 9.3005
R7846 dvdd.n1893 dvdd.n1817 9.3005
R7847 dvdd.n1895 dvdd.n1894 9.3005
R7848 dvdd.n1896 dvdd.n1816 9.3005
R7849 dvdd.n1900 dvdd.n1899 9.3005
R7850 dvdd.n1901 dvdd.n1815 9.3005
R7851 dvdd.n1903 dvdd.n1902 9.3005
R7852 dvdd.n1904 dvdd.n1814 9.3005
R7853 dvdd.n1908 dvdd.n1907 9.3005
R7854 dvdd.n1910 dvdd.n1909 9.3005
R7855 dvdd.n1911 dvdd.n1812 9.3005
R7856 dvdd.n1914 dvdd.n1913 9.3005
R7857 dvdd.n1915 dvdd.n1811 9.3005
R7858 dvdd.n1917 dvdd.n1916 9.3005
R7859 dvdd.n1921 dvdd.n1809 9.3005
R7860 dvdd.n1924 dvdd.n1923 9.3005
R7861 dvdd.n1925 dvdd.n1808 9.3005
R7862 dvdd.n1991 dvdd.n1926 9.3005
R7863 dvdd.n1988 dvdd.n1987 9.3005
R7864 dvdd.n1986 dvdd.n1985 9.3005
R7865 dvdd.n1984 dvdd.n1983 9.3005
R7866 dvdd.n1982 dvdd.n1981 9.3005
R7867 dvdd.n1980 dvdd.n1979 9.3005
R7868 dvdd.n1978 dvdd.n1977 9.3005
R7869 dvdd.n1975 dvdd.n1932 9.3005
R7870 dvdd.n1973 dvdd.n1972 9.3005
R7871 dvdd.n1971 dvdd.n1937 9.3005
R7872 dvdd.n1970 dvdd.n1969 9.3005
R7873 dvdd.n1967 dvdd.n1938 9.3005
R7874 dvdd.n1965 dvdd.n1964 9.3005
R7875 dvdd.n1963 dvdd.n1962 9.3005
R7876 dvdd.n1960 dvdd.n1942 9.3005
R7877 dvdd.n1958 dvdd.n1957 9.3005
R7878 dvdd.n1956 dvdd.n1946 9.3005
R7879 dvdd.n1955 dvdd.n1954 9.3005
R7880 dvdd.n1953 dvdd.n1947 9.3005
R7881 dvdd.n1950 dvdd.n1949 9.3005
R7882 dvdd.n1794 dvdd.n1791 9.3005
R7883 dvdd.n2083 dvdd.n2082 9.3005
R7884 dvdd.n2081 dvdd.n1797 9.3005
R7885 dvdd.n2080 dvdd.n2079 9.3005
R7886 dvdd.n2078 dvdd.n2077 9.3005
R7887 dvdd.n2074 dvdd.n2073 9.3005
R7888 dvdd.n2072 dvdd.n2071 9.3005
R7889 dvdd.n2069 dvdd.n1807 9.3005
R7890 dvdd.n2067 dvdd.n2066 9.3005
R7891 dvdd.n2064 dvdd.n2063 9.3005
R7892 dvdd.n2061 dvdd.n1999 9.3005
R7893 dvdd.n2059 dvdd.n2058 9.3005
R7894 dvdd.n2057 dvdd.n2000 9.3005
R7895 dvdd.n2056 dvdd.n2055 9.3005
R7896 dvdd.n2054 dvdd.n2001 9.3005
R7897 dvdd.n2053 dvdd.n2052 9.3005
R7898 dvdd.n2051 dvdd.n2005 9.3005
R7899 dvdd.n2050 dvdd.n2049 9.3005
R7900 dvdd.n2047 dvdd.n2006 9.3005
R7901 dvdd.n2046 dvdd.n2045 9.3005
R7902 dvdd.n2044 dvdd.n2043 9.3005
R7903 dvdd.n2041 dvdd.n2040 9.3005
R7904 dvdd.n2039 dvdd.n2012 9.3005
R7905 dvdd.n2038 dvdd.n2037 9.3005
R7906 dvdd.n2036 dvdd.n2035 9.3005
R7907 dvdd.n2034 dvdd.n2014 9.3005
R7908 dvdd.n2033 dvdd.n2032 9.3005
R7909 dvdd.n2031 dvdd.n2015 9.3005
R7910 dvdd.n2030 dvdd.n2029 9.3005
R7911 dvdd.n2028 dvdd.n2017 9.3005
R7912 dvdd.n2027 dvdd.n2026 9.3005
R7913 dvdd.n2245 dvdd.n2244 9.3005
R7914 dvdd.n2247 dvdd.n2246 9.3005
R7915 dvdd.n2249 dvdd.n2248 9.3005
R7916 dvdd.n2250 dvdd.n2234 9.3005
R7917 dvdd.n2252 dvdd.n2251 9.3005
R7918 dvdd.n2254 dvdd.n2253 9.3005
R7919 dvdd.n2255 dvdd.n2232 9.3005
R7920 dvdd.n2257 dvdd.n2256 9.3005
R7921 dvdd.n2258 dvdd.n2231 9.3005
R7922 dvdd.n2260 dvdd.n2259 9.3005
R7923 dvdd.n2261 dvdd.n2230 9.3005
R7924 dvdd.n2264 dvdd.n2263 9.3005
R7925 dvdd.n2265 dvdd.n2144 9.3005
R7926 dvdd.n2267 dvdd.n2266 9.3005
R7927 dvdd.n2270 dvdd.n2269 9.3005
R7928 dvdd.n2271 dvdd.n2143 9.3005
R7929 dvdd.n2273 dvdd.n2272 9.3005
R7930 dvdd.n2276 dvdd.n2275 9.3005
R7931 dvdd.n2278 dvdd.n2277 9.3005
R7932 dvdd.n2279 dvdd.n2138 9.3005
R7933 dvdd.n2281 dvdd.n2280 9.3005
R7934 dvdd.n2283 dvdd.n2282 9.3005
R7935 dvdd.n2284 dvdd.n2136 9.3005
R7936 dvdd.n2287 dvdd.n2286 9.3005
R7937 dvdd.n2288 dvdd.n2135 9.3005
R7938 dvdd.n2290 dvdd.n2289 9.3005
R7939 dvdd.n2292 dvdd.n2134 9.3005
R7940 dvdd.n2294 dvdd.n2293 9.3005
R7941 dvdd.n2296 dvdd.n2295 9.3005
R7942 dvdd.n2299 dvdd.n2298 9.3005
R7943 dvdd.n2301 dvdd.n2300 9.3005
R7944 dvdd.n2302 dvdd.n2131 9.3005
R7945 dvdd.n2304 dvdd.n2303 9.3005
R7946 dvdd.n2306 dvdd.n2305 9.3005
R7947 dvdd.n2307 dvdd.n2129 9.3005
R7948 dvdd.n2309 dvdd.n2308 9.3005
R7949 dvdd.n2311 dvdd.n2310 9.3005
R7950 dvdd.n2313 dvdd.n2312 9.3005
R7951 dvdd.n2315 dvdd.n2314 9.3005
R7952 dvdd.n2316 dvdd.n2125 9.3005
R7953 dvdd dvdd.n2318 9.3005
R7954 dvdd.n2319 dvdd.n2124 9.3005
R7955 dvdd.n2321 dvdd.n2320 9.3005
R7956 dvdd.n2325 dvdd.n2122 9.3005
R7957 dvdd.n2328 dvdd.n2327 9.3005
R7958 dvdd.n2329 dvdd.n2121 9.3005
R7959 dvdd.n2331 dvdd.n2330 9.3005
R7960 dvdd.n2332 dvdd.n2120 9.3005
R7961 dvdd.n2333 dvdd.n2118 9.3005
R7962 dvdd.n2334 dvdd.n2117 9.3005
R7963 dvdd.n2338 dvdd.n2337 9.3005
R7964 dvdd.n2340 dvdd.n2339 9.3005
R7965 dvdd.n2341 dvdd.n2114 9.3005
R7966 dvdd.n2343 dvdd.n2342 9.3005
R7967 dvdd.n2345 dvdd.n2344 9.3005
R7968 dvdd.n2346 dvdd.n2111 9.3005
R7969 dvdd.n2348 dvdd.n2347 9.3005
R7970 dvdd.n2350 dvdd.n2349 9.3005
R7971 dvdd.n2352 dvdd.n2093 9.3005
R7972 dvdd.n2353 dvdd.n2352 9.3005
R7973 dvdd.n2352 dvdd.n2103 9.3005
R7974 dvdd.n2352 dvdd.n2095 9.3005
R7975 dvdd.n2156 dvdd.n2155 9.3005
R7976 dvdd.n2158 dvdd.n2151 9.3005
R7977 dvdd.n2160 dvdd.n2159 9.3005
R7978 dvdd.n2162 dvdd.n2161 9.3005
R7979 dvdd.n2226 dvdd.n2149 9.3005
R7980 dvdd.n2226 dvdd.n2225 9.3005
R7981 dvdd.n2222 dvdd.n2221 9.3005
R7982 dvdd.n2218 dvdd.n2174 9.3005
R7983 dvdd.n2217 dvdd.n2216 9.3005
R7984 dvdd.n2215 dvdd.n2176 9.3005
R7985 dvdd.n2214 dvdd.n2213 9.3005
R7986 dvdd.n2212 dvdd.n2177 9.3005
R7987 dvdd.n2211 dvdd.n2210 9.3005
R7988 dvdd.n2209 dvdd.n2179 9.3005
R7989 dvdd.n2208 dvdd.n2207 9.3005
R7990 dvdd.n2206 dvdd.n2205 9.3005
R7991 dvdd.n2204 dvdd.n2182 9.3005
R7992 dvdd.n2203 dvdd.n2202 9.3005
R7993 dvdd.n2201 dvdd.n2200 9.3005
R7994 dvdd.n2199 dvdd.n2186 9.3005
R7995 dvdd.n2198 dvdd.n2197 9.3005
R7996 dvdd.n2196 dvdd.n2187 9.3005
R7997 dvdd.n2421 dvdd.n2420 9.3005
R7998 dvdd.n2423 dvdd.n2422 9.3005
R7999 dvdd.n2425 dvdd.n2424 9.3005
R8000 dvdd.n2427 dvdd.n2410 9.3005
R8001 dvdd.n2431 dvdd.n2430 9.3005
R8002 dvdd.n2432 dvdd.n2409 9.3005
R8003 dvdd.n2434 dvdd.n2433 9.3005
R8004 dvdd.n2435 dvdd.n2408 9.3005
R8005 dvdd.n2437 dvdd.n2436 9.3005
R8006 dvdd.n2439 dvdd.n2438 9.3005
R8007 dvdd.n2440 dvdd.n2406 9.3005
R8008 dvdd.n2443 dvdd.n2442 9.3005
R8009 dvdd.n2445 dvdd.n2444 9.3005
R8010 dvdd.n2450 dvdd.n2449 9.3005
R8011 dvdd.n2451 dvdd.n2404 9.3005
R8012 dvdd.n2453 dvdd.n2452 9.3005
R8013 dvdd.n2455 dvdd.n2402 9.3005
R8014 dvdd.n2457 dvdd.n2456 9.3005
R8015 dvdd.n2464 dvdd.n2463 9.3005
R8016 dvdd.n2469 dvdd.n2468 9.3005
R8017 dvdd.n2470 dvdd.n2400 9.3005
R8018 dvdd.n2472 dvdd.n2471 9.3005
R8019 dvdd.n2479 dvdd.n2398 9.3005
R8020 dvdd.n2481 dvdd.n2480 9.3005
R8021 dvdd.n2483 dvdd.n2396 9.3005
R8022 dvdd.n2486 dvdd.n2485 9.3005
R8023 dvdd.n2489 dvdd.n2488 9.3005
R8024 dvdd.n2490 dvdd.n2390 9.3005
R8025 dvdd.n2496 dvdd.n2495 9.3005
R8026 dvdd.n2497 dvdd.n2389 9.3005
R8027 dvdd.n2499 dvdd.n2498 9.3005
R8028 dvdd.n2501 dvdd.n2500 9.3005
R8029 dvdd.n2502 dvdd.n2386 9.3005
R8030 dvdd.n2554 dvdd.n2553 9.3005
R8031 dvdd.n2552 dvdd.n2387 9.3005
R8032 dvdd.n2551 dvdd.n2550 9.3005
R8033 dvdd.n2549 dvdd.n2503 9.3005
R8034 dvdd.n2547 dvdd.n2509 9.3005
R8035 dvdd.n2546 dvdd.n2515 9.3005
R8036 dvdd.n2545 dvdd.n2544 9.3005
R8037 dvdd.n2543 dvdd.n2542 9.3005
R8038 dvdd.n2540 dvdd.n2518 9.3005
R8039 dvdd.n2539 dvdd.n2538 9.3005
R8040 dvdd.n2537 dvdd.n2536 9.3005
R8041 dvdd.n2535 dvdd.n2534 9.3005
R8042 dvdd.n2533 dvdd.n2522 9.3005
R8043 dvdd.n2532 dvdd.n2531 9.3005
R8044 dvdd.n2529 dvdd.n2523 9.3005
R8045 dvdd.n2528 dvdd.n2527 9.3005
R8046 dvdd.n2367 dvdd.n2363 9.3005
R8047 dvdd.n2641 dvdd.n2640 9.3005
R8048 dvdd.n2639 dvdd.n2368 9.3005
R8049 dvdd.n2638 dvdd.n2637 9.3005
R8050 dvdd.n2636 dvdd.n2635 9.3005
R8051 dvdd.n2634 dvdd.n2378 9.3005
R8052 dvdd.n2633 dvdd.n2383 9.3005
R8053 dvdd.n2632 dvdd.n2631 9.3005
R8054 dvdd.n2630 dvdd.n2558 9.3005
R8055 dvdd.n2629 dvdd.n2628 9.3005
R8056 dvdd.n2627 dvdd.n2559 9.3005
R8057 dvdd.n2625 dvdd.n2624 9.3005
R8058 dvdd.n2623 dvdd.n2563 9.3005
R8059 dvdd.n2622 dvdd.n2621 9.3005
R8060 dvdd.n2620 dvdd.n2619 9.3005
R8061 dvdd.n2618 dvdd.n2565 9.3005
R8062 dvdd.n2617 dvdd.n2616 9.3005
R8063 dvdd.n2613 dvdd.n2566 9.3005
R8064 dvdd.n2612 dvdd.n2611 9.3005
R8065 dvdd.n2610 dvdd.n2567 9.3005
R8066 dvdd.n2609 dvdd.n2608 9.3005
R8067 dvdd.n2607 dvdd.n2568 9.3005
R8068 dvdd.n2606 dvdd.n2605 9.3005
R8069 dvdd.n2604 dvdd.n2603 9.3005
R8070 dvdd.n2601 dvdd.n2574 9.3005
R8071 dvdd.n2600 dvdd.n2575 9.3005
R8072 dvdd.n2599 dvdd.n2598 9.3005
R8073 dvdd.n2597 dvdd.n2596 9.3005
R8074 dvdd.n2595 dvdd.n2594 9.3005
R8075 dvdd.n2593 dvdd.n2578 9.3005
R8076 dvdd.n2592 dvdd.n2591 9.3005
R8077 dvdd.n2589 dvdd.n2579 9.3005
R8078 dvdd.n3093 dvdd.n3092 9.3005
R8079 dvdd.n2893 dvdd.n2892 9.3005
R8080 dvdd.n2894 dvdd.n2886 9.3005
R8081 dvdd.n2896 dvdd.n2895 9.3005
R8082 dvdd.n2898 dvdd.n2884 9.3005
R8083 dvdd.n2902 dvdd.n2901 9.3005
R8084 dvdd.n2903 dvdd.n2883 9.3005
R8085 dvdd.n2905 dvdd.n2904 9.3005
R8086 dvdd.n2907 dvdd.n2881 9.3005
R8087 dvdd.n2911 dvdd.n2910 9.3005
R8088 dvdd.n2913 dvdd.n2912 9.3005
R8089 dvdd.n2915 dvdd.n2877 9.3005
R8090 dvdd.n2917 dvdd.n2916 9.3005
R8091 dvdd.n2919 dvdd.n2918 9.3005
R8092 dvdd.n2922 dvdd.n2921 9.3005
R8093 dvdd.n2923 dvdd.n2875 9.3005
R8094 dvdd.n2925 dvdd.n2924 9.3005
R8095 dvdd.n2926 dvdd.n2873 9.3005
R8096 dvdd.n3080 dvdd.n3027 9.3005
R8097 dvdd.n3079 dvdd.n3078 9.3005
R8098 dvdd.n3077 dvdd.n3029 9.3005
R8099 dvdd.n3076 dvdd.n3075 9.3005
R8100 dvdd.n3073 dvdd.n3072 9.3005
R8101 dvdd.n3071 dvdd.n3070 9.3005
R8102 dvdd.n3069 dvdd.n3031 9.3005
R8103 dvdd.n3067 dvdd.n3066 9.3005
R8104 dvdd.n3065 dvdd.n3064 9.3005
R8105 dvdd.n3061 dvdd.n3035 9.3005
R8106 dvdd.n3059 dvdd.n3058 9.3005
R8107 dvdd.n3057 dvdd.n3037 9.3005
R8108 dvdd.n3056 dvdd.n3055 9.3005
R8109 dvdd.n3052 dvdd.n3038 9.3005
R8110 dvdd.n3050 dvdd.n3049 9.3005
R8111 dvdd.n3048 dvdd.n3040 9.3005
R8112 dvdd.n3047 dvdd.n3046 9.3005
R8113 dvdd.n3023 dvdd.n2970 9.3005
R8114 dvdd.n3022 dvdd.n3021 9.3005
R8115 dvdd.n3020 dvdd.n2972 9.3005
R8116 dvdd.n3019 dvdd.n3018 9.3005
R8117 dvdd.n3016 dvdd.n3015 9.3005
R8118 dvdd.n3014 dvdd.n3013 9.3005
R8119 dvdd.n3012 dvdd.n2974 9.3005
R8120 dvdd.n3010 dvdd.n3009 9.3005
R8121 dvdd.n3008 dvdd.n3007 9.3005
R8122 dvdd.n3004 dvdd.n2978 9.3005
R8123 dvdd.n3002 dvdd.n3001 9.3005
R8124 dvdd.n3000 dvdd.n2980 9.3005
R8125 dvdd.n2999 dvdd.n2998 9.3005
R8126 dvdd.n2995 dvdd.n2981 9.3005
R8127 dvdd.n2993 dvdd.n2992 9.3005
R8128 dvdd.n2991 dvdd.n2983 9.3005
R8129 dvdd.n2990 dvdd.n2989 9.3005
R8130 dvdd.n2862 dvdd.n2861 9.3005
R8131 dvdd.n2869 dvdd.n2803 9.3005
R8132 dvdd.n2868 dvdd.n2867 9.3005
R8133 dvdd.n2866 dvdd.n2805 9.3005
R8134 dvdd.n2865 dvdd.n2864 9.3005
R8135 dvdd.n2860 dvdd.n2859 9.3005
R8136 dvdd.n2858 dvdd.n2807 9.3005
R8137 dvdd.n2857 dvdd.n2856 9.3005
R8138 dvdd.n2855 dvdd.n2854 9.3005
R8139 dvdd.n2853 dvdd.n2852 9.3005
R8140 dvdd.n2851 dvdd.n2850 9.3005
R8141 dvdd.n2849 dvdd.n2811 9.3005
R8142 dvdd.n2845 dvdd.n2844 9.3005
R8143 dvdd.n2843 dvdd.n2842 9.3005
R8144 dvdd.n2841 dvdd.n2815 9.3005
R8145 dvdd.n2839 dvdd.n2838 9.3005
R8146 dvdd.n2837 dvdd.n2817 9.3005
R8147 dvdd.n2836 dvdd.n2835 9.3005
R8148 dvdd.n2832 dvdd.n2818 9.3005
R8149 dvdd.n2830 dvdd.n2829 9.3005
R8150 dvdd.n2828 dvdd.n2820 9.3005
R8151 dvdd.n2827 dvdd.n2826 9.3005
R8152 dvdd.n2769 dvdd.n2768 9.3005
R8153 dvdd.n2773 dvdd.n2772 9.3005
R8154 dvdd.n2777 dvdd.n2776 9.3005
R8155 dvdd.n2781 dvdd.n2780 9.3005
R8156 dvdd.n2785 dvdd.n2784 9.3005
R8157 dvdd.n2789 dvdd.n2788 9.3005
R8158 dvdd.n2793 dvdd.n2792 9.3005
R8159 dvdd.n2797 dvdd.n2796 9.3005
R8160 dvdd.n2801 dvdd.n2800 9.3005
R8161 dvdd.n2750 dvdd.n2749 9.3005
R8162 dvdd.n2746 dvdd.n2745 9.3005
R8163 dvdd.n2742 dvdd.n2741 9.3005
R8164 dvdd.n2738 dvdd.n2737 9.3005
R8165 dvdd.n2734 dvdd.n2733 9.3005
R8166 dvdd.n2730 dvdd.n2729 9.3005
R8167 dvdd.n2726 dvdd.n2725 9.3005
R8168 dvdd.n2722 dvdd.n2721 9.3005
R8169 dvdd.n2718 dvdd.n2717 9.3005
R8170 dvdd.n3146 dvdd.n3137 9.3005
R8171 dvdd.n2834 dvdd.n2817 9.25588
R8172 dvdd.n254 dvdd.n223 9.09802
R8173 dvdd.n241 dvdd.n229 9.09802
R8174 dvdd.n275 dvdd.n274 9.09802
R8175 dvdd.n261 dvdd.n222 9.09802
R8176 dvdd.n300 dvdd.n82 9.09802
R8177 dvdd.n319 dvdd.n318 9.09802
R8178 dvdd.n130 dvdd.n100 9.09802
R8179 dvdd.n117 dvdd.n105 9.09802
R8180 dvdd.n175 dvdd.n162 9.09802
R8181 dvdd.n188 dvdd.n156 9.09802
R8182 dvdd.n414 dvdd.n369 9.09802
R8183 dvdd.n455 dvdd.n454 9.09802
R8184 dvdd.n710 dvdd.n707 9.09802
R8185 dvdd.n722 dvdd.n636 9.09802
R8186 dvdd.n685 dvdd.n650 9.09802
R8187 dvdd.n879 dvdd.n878 9.09802
R8188 dvdd.n1295 dvdd.n1236 9.09802
R8189 dvdd.n1843 dvdd.n1832 9.09802
R8190 dvdd.n2062 dvdd.n2061 9.09802
R8191 dvdd.n2046 dvdd.n2007 9.09802
R8192 dvdd.n2315 dvdd.n2127 9.09802
R8193 dvdd.n2317 dvdd.n2316 9.09802
R8194 dvdd.n2183 dvdd.n2182 9.09802
R8195 dvdd.n1138 dvdd.n1120 9.03579
R8196 dvdd.n1620 dvdd.n1507 9.03579
R8197 dvdd.n1747 dvdd.n1746 9.03579
R8198 dvdd.n1721 dvdd.n1720 9.03579
R8199 dvdd.n1883 dvdd.n1882 9.03579
R8200 dvdd.n2482 dvdd.n2481 8.99224
R8201 dvdd.n2454 dvdd.n2453 8.99224
R8202 dvdd.n2164 dvdd.n2163 8.9761
R8203 dvdd.n2147 dvdd 8.9245
R8204 dvdd.n3154 dvdd.n3096 8.89596
R8205 dvdd.n2835 dvdd.n2834 8.86204
R8206 dvdd.n1965 dvdd.n1941 8.77764
R8207 dvdd dvdd.n3095 8.72508
R8208 dvdd.n979 dvdd.n978 8.65932
R8209 dvdd.n1780 dvdd.n1779 8.65932
R8210 dvdd.n415 dvdd.n414 8.49383
R8211 dvdd.n2312 dvdd.n2311 8.44958
R8212 dvdd.n2207 dvdd.n2206 8.44958
R8213 dvdd.n2449 dvdd.n2445 8.44958
R8214 dvdd.t580 dvdd.t762 8.39273
R8215 dvdd dvdd.t1343 8.39273
R8216 dvdd.t313 dvdd.t1652 8.39273
R8217 dvdd.t1315 dvdd.t1661 8.39273
R8218 dvdd.t1407 dvdd.t1391 8.39273
R8219 dvdd.t1447 dvdd.t1197 8.39273
R8220 dvdd.t944 dvdd.t669 8.39273
R8221 dvdd.n454 dvdd.n453 8.35752
R8222 dvdd.n720 dvdd.n639 8.35752
R8223 dvdd.n2467 dvdd.n2466 8.35752
R8224 dvdd.n1000 dvdd.n999 8.28285
R8225 dvdd.n1166 dvdd.n1165 8.28285
R8226 dvdd.n1316 dvdd.n1315 8.28285
R8227 dvdd.n2900 dvdd.n2883 8.2416
R8228 dvdd.n2941 dvdd.n2940 8.2025
R8229 dvdd.n3054 dvdd.n3037 8.13023
R8230 dvdd.n2997 dvdd.n2980 8.13023
R8231 dvdd.n1075 dvdd.n1061 7.90638
R8232 dvdd.n2901 dvdd.n2900 7.89091
R8233 dvdd.n448 dvdd.n446 7.8286
R8234 dvdd.n3055 dvdd.n3054 7.78428
R8235 dvdd.n2998 dvdd.n2997 7.78428
R8236 dvdd.n695 dvdd.n693 7.75995
R8237 dvdd.n1858 dvdd.n1856 7.75995
R8238 dvdd.n872 dvdd.n871 7.72281
R8239 dvdd.n2048 dvdd.n2047 7.72281
R8240 dvdd.n2082 dvdd.n2081 7.6805
R8241 dvdd.n1381 dvdd.n1380 7.52991
R8242 dvdd.n1765 dvdd.n1764 7.52991
R8243 dvdd.n687 dvdd.n686 7.40546
R8244 dvdd.n2165 dvdd.n2164 7.39867
R8245 dvdd.n2290 dvdd.n2135 7.21067
R8246 dvdd.n515 dvdd.n514 7.15344
R8247 dvdd.n1743 dvdd.n1691 7.15344
R8248 dvdd.n1735 dvdd.n1734 7.15344
R8249 dvdd.n1700 dvdd.n1698 7.15344
R8250 dvdd.n1723 dvdd.n1722 7.15344
R8251 dvdd.n2425 dvdd.n2411 7.12524
R8252 dvdd.n144 dvdd.n143 7.11866
R8253 dvdd.n1310 dvdd.n1229 7.0881
R8254 dvdd.n2541 dvdd.n2540 7.0168
R8255 dvdd.n740 dvdd.n629 6.94907
R8256 dvdd.n1593 dvdd.n1520 6.8512
R8257 dvdd.n986 dvdd.n985 6.77697
R8258 dvdd.n2347 dvdd.n2110 6.77697
R8259 dvdd.n2159 dvdd.n2150 6.73838
R8260 dvdd.t409 dvdd 6.71428
R8261 dvdd.t1297 dvdd.t903 6.71428
R8262 dvdd dvdd.t136 6.71428
R8263 dvdd.t78 dvdd.t260 6.71428
R8264 dvdd.t530 dvdd.t1181 6.71428
R8265 dvdd.t146 dvdd.t1009 6.71428
R8266 dvdd.n437 dvdd.n362 6.66496
R8267 dvdd.n706 dvdd.n705 6.66496
R8268 dvdd.n866 dvdd.n865 6.66496
R8269 dvdd.n2485 dvdd.n2484 6.66496
R8270 dvdd.n2473 dvdd.n2472 6.66496
R8271 dvdd.n2456 dvdd.n2401 6.66496
R8272 dvdd.n2764 dvdd.n2763 6.58874
R8273 dvdd.n2755 dvdd.n2754 6.58874
R8274 dvdd.n1354 dvdd.n1347 6.58336
R8275 dvdd.n2060 dvdd.n2059 6.55918
R8276 dvdd.n2440 dvdd.n2439 6.52104
R8277 dvdd.n2395 dvdd.n2394 6.48583
R8278 dvdd.n2473 dvdd.n2399 6.45339
R8279 dvdd.n1023 dvdd.n933 6.4005
R8280 dvdd.n1906 dvdd.n1813 6.4005
R8281 dvdd.n2226 dvdd.n2148 6.4005
R8282 dvdd.n1849 dvdd.n1848 6.34761
R8283 dvdd.n727 dvdd.n726 6.29507
R8284 dvdd.n2823 dvdd.n2821 6.14225
R8285 dvdd.n444 dvdd.n360 6.13604
R8286 dvdd.n1520 dvdd.n1516 6.13008
R8287 dvdd.n2832 dvdd.n2831 6.10512
R8288 dvdd.n1656 dvdd.n1636 6.0706
R8289 dvdd.n3143 dvdd.t1352 6.06249
R8290 dvdd.n2268 dvdd.n2267 6.04885
R8291 dvdd.n447 dvdd.n357 6.03025
R8292 dvdd.n716 dvdd.n715 6.03025
R8293 dvdd.n1017 dvdd.n1016 6.02403
R8294 dvdd.n1899 dvdd.n1898 6.02403
R8295 dvdd.n2464 dvdd.n2401 5.98311
R8296 dvdd.n2966 dvdd.n2947 5.96824
R8297 dvdd.t701 dvdd.n2947 5.96824
R8298 dvdd.n2962 dvdd.n2961 5.96824
R8299 dvdd.t701 dvdd.n2962 5.96824
R8300 dvdd.n3150 dvdd.n3099 5.9447
R8301 dvdd.n3136 dvdd.n3099 5.94023
R8302 dvdd.n2889 dvdd.n2887 5.87299
R8303 dvdd.n1962 dvdd.n1941 5.85193
R8304 dvdd.n1961 dvdd.n1960 5.85193
R8305 dvdd.n3043 dvdd.n3041 5.84114
R8306 dvdd.n2986 dvdd.n2984 5.84114
R8307 dvdd.n3094 dvdd 5.83822
R8308 dvdd.n2840 dvdd.n2839 5.71127
R8309 dvdd.n391 dvdd.n390 5.66204
R8310 dvdd.n392 dvdd.n391 5.66204
R8311 dvdd.n396 dvdd.n395 5.66204
R8312 dvdd.n397 dvdd.n396 5.66204
R8313 dvdd.n397 dvdd.n372 5.66204
R8314 dvdd.n401 dvdd.n372 5.66204
R8315 dvdd.n402 dvdd.n401 5.66204
R8316 dvdd.n403 dvdd.n402 5.66204
R8317 dvdd.n422 dvdd.n367 5.66204
R8318 dvdd.n425 dvdd.n424 5.66204
R8319 dvdd.n425 dvdd.n365 5.66204
R8320 dvdd.n429 dvdd.n365 5.66204
R8321 dvdd.n430 dvdd.n429 5.66204
R8322 dvdd.n571 dvdd.n570 5.66204
R8323 dvdd.n570 dvdd.n569 5.66204
R8324 dvdd.n566 dvdd.n565 5.66204
R8325 dvdd.n565 dvdd.n564 5.66204
R8326 dvdd.n564 dvdd.n544 5.66204
R8327 dvdd.n560 dvdd.n544 5.66204
R8328 dvdd.n560 dvdd.n559 5.66204
R8329 dvdd.n559 dvdd.n558 5.66204
R8330 dvdd.n860 dvdd.n859 5.66204
R8331 dvdd.n859 dvdd.n858 5.66204
R8332 dvdd.n855 dvdd.n854 5.66204
R8333 dvdd.n854 dvdd.n853 5.66204
R8334 dvdd.n853 dvdd.n833 5.66204
R8335 dvdd.n849 dvdd.n833 5.66204
R8336 dvdd.n849 dvdd.n848 5.66204
R8337 dvdd.n848 dvdd.n847 5.66204
R8338 dvdd.n2250 dvdd.n2249 5.66204
R8339 dvdd.n2251 dvdd.n2250 5.66204
R8340 dvdd.n2255 dvdd.n2254 5.66204
R8341 dvdd.n2256 dvdd.n2255 5.66204
R8342 dvdd.n2256 dvdd.n2231 5.66204
R8343 dvdd.n2260 dvdd.n2231 5.66204
R8344 dvdd.n2261 dvdd.n2260 5.66204
R8345 dvdd.n2263 dvdd.n2261 5.66204
R8346 dvdd.n2302 dvdd.n2301 5.66204
R8347 dvdd.n2303 dvdd.n2302 5.66204
R8348 dvdd.n2307 dvdd.n2306 5.66204
R8349 dvdd.n2308 dvdd.n2307 5.66204
R8350 dvdd.n2293 dvdd.n2292 5.66204
R8351 dvdd.n2279 dvdd.n2278 5.66204
R8352 dvdd.n2280 dvdd.n2279 5.66204
R8353 dvdd.n2284 dvdd.n2283 5.66204
R8354 dvdd.n2286 dvdd.n2284 5.66204
R8355 dvdd.n2218 dvdd.n2217 5.66204
R8356 dvdd.n2217 dvdd.n2176 5.66204
R8357 dvdd.n2213 dvdd.n2212 5.66204
R8358 dvdd.n2212 dvdd.n2211 5.66204
R8359 dvdd.n2211 dvdd.n2179 5.66204
R8360 dvdd.n1048 dvdd.n1047 5.64756
R8361 dvdd.n1160 dvdd.n1111 5.64756
R8362 dvdd.n2847 dvdd.n2845 5.51435
R8363 dvdd.n433 dvdd.n432 5.48759
R8364 dvdd.n2898 dvdd.n2897 5.43612
R8365 dvdd.n2221 dvdd.n2175 5.42606
R8366 dvdd.n670 dvdd.n654 5.40233
R8367 dvdd.n3052 dvdd.n3051 5.36266
R8368 dvdd.n2995 dvdd.n2994 5.36266
R8369 dvdd.n390 dvdd.n376 5.29281
R8370 dvdd.n403 dvdd.n370 5.29281
R8371 dvdd.n418 dvdd.n416 5.29281
R8372 dvdd.n431 dvdd.n430 5.29281
R8373 dvdd.n571 dvdd.n540 5.29281
R8374 dvdd.n558 dvdd.n546 5.29281
R8375 dvdd.n860 dvdd.n829 5.29281
R8376 dvdd.n847 dvdd.n835 5.29281
R8377 dvdd.n2249 dvdd.n2235 5.29281
R8378 dvdd.n2263 dvdd.n2262 5.29281
R8379 dvdd.n2301 dvdd.n2132 5.29281
R8380 dvdd.n2308 dvdd.n2128 5.29281
R8381 dvdd.n2292 dvdd.n2291 5.29281
R8382 dvdd.n2293 dvdd.n2133 5.29281
R8383 dvdd.n2278 dvdd.n2139 5.29281
R8384 dvdd.n2286 dvdd.n2285 5.29281
R8385 dvdd.n2180 dvdd.n2179 5.29281
R8386 dvdd.n2442 dvdd.n2441 5.29281
R8387 dvdd.n2442 dvdd.n2405 5.29281
R8388 dvdd.n2393 dvdd.n2392 5.29117
R8389 dvdd.n438 dvdd.n437 5.28976
R8390 dvdd.n786 dvdd.n785 5.27109
R8391 dvdd.n1282 dvdd.n1281 5.27109
R8392 dvdd.n1468 dvdd.n1213 5.27109
R8393 dvdd.n252 dvdd.n225 5.18397
R8394 dvdd.n219 dvdd.n217 5.18397
R8395 dvdd.n307 dvdd.n306 5.18397
R8396 dvdd.n128 dvdd.n101 5.18397
R8397 dvdd.n177 dvdd.n160 5.18397
R8398 dvdd.n440 dvdd.n439 5.18397
R8399 dvdd.n710 dvdd.n709 5.18397
R8400 dvdd.n689 dvdd.n688 5.18397
R8401 dvdd.n821 dvdd.n819 5.18397
R8402 dvdd.n1304 dvdd.n1303 5.18397
R8403 dvdd.n1851 dvdd.n1850 5.18397
R8404 dvdd.n2449 dvdd.n2447 5.18397
R8405 dvdd.n2872 dvdd 5.14764
R8406 dvdd.n3026 dvdd 5.14243
R8407 dvdd.n3083 dvdd 5.13722
R8408 dvdd.n2906 dvdd.n2905 5.08543
R8409 dvdd dvdd.t270 5.03584
R8410 dvdd.t604 dvdd.t1405 5.03584
R8411 dvdd.t901 dvdd.t1233 5.03584
R8412 dvdd.t1051 dvdd.t1372 5.03584
R8413 dvdd.t735 dvdd.t437 5.03584
R8414 dvdd.t677 dvdd.t894 5.03584
R8415 dvdd.t824 dvdd.t4 5.03584
R8416 dvdd.n2274 dvdd.n2273 5.03171
R8417 dvdd.n3060 dvdd.n3059 5.01672
R8418 dvdd.n3003 dvdd.n3002 5.01672
R8419 dvdd.n2173 dvdd.n2172 4.94058
R8420 dvdd.n999 dvdd.n998 4.89462
R8421 dvdd.n1009 dvdd.n938 4.89462
R8422 dvdd.n1464 dvdd.n1216 4.89462
R8423 dvdd.n1743 dvdd.n1742 4.89462
R8424 dvdd.n1723 dvdd.n1704 4.89462
R8425 dvdd.n1880 dvdd.n1879 4.89462
R8426 dvdd.n1975 dvdd.n1974 4.89462
R8427 dvdd.n701 dvdd.n643 4.79796
R8428 dvdd.n1953 dvdd.n1952 4.75479
R8429 dvdd.n213 dvdd.n211 4.67352
R8430 dvdd.n137 dvdd.n96 4.67352
R8431 dvdd.n137 dvdd.n136 4.67352
R8432 dvdd.n678 dvdd.n675 4.67352
R8433 dvdd.n671 dvdd.n652 4.67352
R8434 dvdd.n780 dvdd.n779 4.67352
R8435 dvdd.n890 dvdd.n889 4.67352
R8436 dvdd.n970 dvdd.n966 4.67352
R8437 dvdd.n1038 dvdd.n931 4.67352
R8438 dvdd.n1154 dvdd.n1153 4.67352
R8439 dvdd.n1150 dvdd.n1149 4.67352
R8440 dvdd.n1606 dvdd.n1512 4.67352
R8441 dvdd.n1607 dvdd.n1606 4.67352
R8442 dvdd.n1584 dvdd.n1583 4.67352
R8443 dvdd.n1588 dvdd.n1584 4.67352
R8444 dvdd.n1923 dvdd.n1921 4.67352
R8445 dvdd.n1985 dvdd.n1984 4.67352
R8446 dvdd.n2159 dvdd.n2158 4.67352
R8447 dvdd.n2327 dvdd.n2325 4.67352
R8448 dvdd.n2608 dvdd.n2607 4.67352
R8449 dvdd.n2607 dvdd.n2606 4.67352
R8450 dvdd.n2596 dvdd.n2595 4.67352
R8451 dvdd.n2595 dvdd.n2578 4.67352
R8452 dvdd.n2591 dvdd.n2578 4.67352
R8453 dvdd.n675 dvdd.n652 4.67352
R8454 dvdd.n2069 dvdd.n2068 4.62834
R8455 dvdd.n575 dvdd.n539 4.62124
R8456 dvdd.n1069 dvdd.n1064 4.62124
R8457 dvdd.n1290 dvdd.n1239 4.62124
R8458 dvdd.n2548 dvdd.n2507 4.62124
R8459 dvdd.n2547 dvdd.n2510 4.62124
R8460 dvdd.n2633 dvdd.n2384 4.62124
R8461 dvdd.n435 dvdd.n363 4.62124
R8462 dvdd.n704 dvdd.n703 4.62124
R8463 dvdd.n1581 dvdd.n1531 4.62124
R8464 dvdd.n2487 dvdd.n2395 4.62124
R8465 dvdd.n2158 dvdd.n2157 4.57193
R8466 dvdd.n249 dvdd.n225 4.54926
R8467 dvdd.n269 dvdd.n219 4.54926
R8468 dvdd.n308 dvdd.n307 4.54926
R8469 dvdd.n125 dvdd.n101 4.54926
R8470 dvdd.n180 dvdd.n160 4.54926
R8471 dvdd.n441 dvdd.n440 4.54926
R8472 dvdd.n688 dvdd.n647 4.54926
R8473 dvdd.n873 dvdd.n821 4.54926
R8474 dvdd.n1301 dvdd.n1234 4.54926
R8475 dvdd.n1303 dvdd.n1302 4.54926
R8476 dvdd.n1852 dvdd.n1851 4.54926
R8477 dvdd.n2003 dvdd.n2000 4.54926
R8478 dvdd.n2055 dvdd.n2004 4.54926
R8479 dvdd.n326 dvdd.n74 4.51401
R8480 dvdd.n205 dvdd.n204 4.51401
R8481 dvdd.n609 dvdd.n331 4.51401
R8482 dvdd.n346 dvdd.n345 4.51401
R8483 dvdd.n910 dvdd.n614 4.51401
R8484 dvdd.n901 dvdd.n900 4.51401
R8485 dvdd.n1199 dvdd.n915 4.51401
R8486 dvdd.n1192 dvdd.n1191 4.51401
R8487 dvdd.n1483 dvdd.n1204 4.51401
R8488 dvdd.n1476 dvdd.n1475 4.51401
R8489 dvdd.n1784 dvdd.n1488 4.51401
R8490 dvdd.n1775 dvdd.n1774 4.51401
R8491 dvdd.n2086 dvdd.n1789 4.51401
R8492 dvdd.n1805 dvdd.n1804 4.51401
R8493 dvdd.n2356 dvdd.n2091 4.51401
R8494 dvdd.n2102 dvdd.n2101 4.51401
R8495 dvdd.n2644 dvdd.n2361 4.51401
R8496 dvdd.n2377 dvdd.n2376 4.51401
R8497 dvdd.n325 dvdd.n324 4.5005
R8498 dvdd.n199 dvdd.n76 4.5005
R8499 dvdd.n203 dvdd.n202 4.5005
R8500 dvdd.n608 dvdd.n607 4.5005
R8501 dvdd.n340 dvdd.n334 4.5005
R8502 dvdd.n344 dvdd.n343 4.5005
R8503 dvdd.n909 dvdd.n908 4.5005
R8504 dvdd.n896 dvdd.n617 4.5005
R8505 dvdd.n899 dvdd.n622 4.5005
R8506 dvdd.n1198 dvdd.n1197 4.5005
R8507 dvdd.n1187 dvdd.n918 4.5005
R8508 dvdd.n1190 dvdd.n924 4.5005
R8509 dvdd.n1482 dvdd.n1481 4.5005
R8510 dvdd.n1471 dvdd.n1207 4.5005
R8511 dvdd.n1474 dvdd.n1210 4.5005
R8512 dvdd.n1783 dvdd.n1782 4.5005
R8513 dvdd.n1770 dvdd.n1491 4.5005
R8514 dvdd.n1773 dvdd.n1496 4.5005
R8515 dvdd.n2085 dvdd.n2084 4.5005
R8516 dvdd.n1799 dvdd.n1792 4.5005
R8517 dvdd.n1803 dvdd.n1802 4.5005
R8518 dvdd.n2355 dvdd.n2354 4.5005
R8519 dvdd.n2097 dvdd.n2094 4.5005
R8520 dvdd.n2100 dvdd.n2096 4.5005
R8521 dvdd.n2643 dvdd.n2642 4.5005
R8522 dvdd.n2371 dvdd.n2364 4.5005
R8523 dvdd.n2375 dvdd.n2374 4.5005
R8524 dvdd.n2943 dvdd.n2942 4.5005
R8525 dvdd.n2341 dvdd.n2340 4.48528
R8526 dvdd.n1611 dvdd.n1608 4.47034
R8527 dvdd.n2074 dvdd.n1806 4.47034
R8528 dvdd.n439 dvdd.n438 4.44348
R8529 dvdd.n740 dvdd.n739 4.38907
R8530 dvdd.n1367 dvdd.n1366 4.38907
R8531 dvdd.n1960 dvdd.n1959 4.38907
R8532 dvdd.n234 dvdd.n233 4.36875
R8533 dvdd.n213 dvdd.n212 4.36875
R8534 dvdd.n296 dvdd.n83 4.36875
R8535 dvdd.n136 dvdd.n135 4.36875
R8536 dvdd.n152 dvdd.n151 4.36875
R8537 dvdd.n167 dvdd.n164 4.36875
R8538 dvdd.n501 dvdd.n500 4.36875
R8539 dvdd.n667 dvdd.n655 4.36875
R8540 dvdd.n779 dvdd.n778 4.36875
R8541 dvdd.n889 dvdd.n624 4.36875
R8542 dvdd.n1039 dvdd.n1038 4.36875
R8543 dvdd.n1156 dvdd.n1112 4.36875
R8544 dvdd.n1147 dvdd.n1117 4.36875
R8545 dvdd.n1611 dvdd.n1610 4.36875
R8546 dvdd.n1923 dvdd.n1922 4.36875
R8547 dvdd.n1984 dvdd.n1929 4.36875
R8548 dvdd.n2071 dvdd.n2070 4.36875
R8549 dvdd.n2337 dvdd.n2116 4.36875
R8550 dvdd.n2327 dvdd.n2326 4.36875
R8551 dvdd.n2603 dvdd.n2602 4.36875
R8552 dvdd.n2591 dvdd.n2590 4.36875
R8553 dvdd.n2447 dvdd.n2446 4.33769
R8554 dvdd.n3091 dvdd.n3090 4.32258
R8555 dvdd.n2799 dvdd.n9 4.32258
R8556 dvdd.n2795 dvdd.n16 4.32258
R8557 dvdd.n2791 dvdd.n23 4.32258
R8558 dvdd.n2787 dvdd.n30 4.32258
R8559 dvdd.n2783 dvdd.n37 4.32258
R8560 dvdd.n2779 dvdd.n44 4.32258
R8561 dvdd.n2775 dvdd.n51 4.32258
R8562 dvdd.n2771 dvdd.n58 4.32258
R8563 dvdd.n2767 dvdd.n65 4.32258
R8564 dvdd.n2719 dvdd.n2715 4.32258
R8565 dvdd.n2723 dvdd.n2708 4.32258
R8566 dvdd.n2727 dvdd.n2701 4.32258
R8567 dvdd.n2731 dvdd.n2694 4.32258
R8568 dvdd.n2735 dvdd.n2687 4.32258
R8569 dvdd.n2739 dvdd.n2680 4.32258
R8570 dvdd.n2743 dvdd.n2673 4.32258
R8571 dvdd.n2747 dvdd.n2666 4.32258
R8572 dvdd.n2751 dvdd.n2659 4.32258
R8573 dvdd.n3149 dvdd.n3148 4.29291
R8574 dvdd.n3137 dvdd.n3136 4.26836
R8575 dvdd.n2577 dvdd.n2576 4.26717
R8576 dvdd.n141 dvdd.n96 4.18384
R8577 dvdd.n1601 dvdd.n1600 4.16558
R8578 dvdd.n709 dvdd.n708 4.12612
R8579 dvdd.n2608 dvdd.n2571 4.11479
R8580 dvdd dvdd.n3155 4.0955
R8581 dvdd.n383 dvdd.n379 4.02033
R8582 dvdd.n383 dvdd.n382 4.02033
R8583 dvdd.n575 dvdd.n537 4.02033
R8584 dvdd.n554 dvdd.n549 4.02033
R8585 dvdd.n554 dvdd.n552 4.02033
R8586 dvdd.n663 dvdd.n658 4.02033
R8587 dvdd.n663 dvdd.n662 4.02033
R8588 dvdd.n864 dvdd.n827 4.02033
R8589 dvdd.n843 dvdd.n838 4.02033
R8590 dvdd.n843 dvdd.n841 4.02033
R8591 dvdd.n960 dvdd.n956 4.02033
R8592 dvdd.n960 dvdd.n959 4.02033
R8593 dvdd.n1129 dvdd.n1125 4.02033
R8594 dvdd.n1129 dvdd.n1128 4.02033
R8595 dvdd.n1263 dvdd.n1259 4.02033
R8596 dvdd.n1263 dvdd.n1262 4.02033
R8597 dvdd.n1420 dvdd.n1416 4.02033
R8598 dvdd.n1420 dvdd.n1419 4.02033
R8599 dvdd.n1551 dvdd.n1546 4.02033
R8600 dvdd.n1551 dvdd.n1550 4.02033
R8601 dvdd.n1714 dvdd.n1709 4.02033
R8602 dvdd.n1714 dvdd.n1712 4.02033
R8603 dvdd.n1839 dvdd.n1835 4.02033
R8604 dvdd.n1839 dvdd.n1838 4.02033
R8605 dvdd.n1998 dvdd.n1997 4.02033
R8606 dvdd.n2025 dvdd.n2020 4.02033
R8607 dvdd.n2025 dvdd.n2023 4.02033
R8608 dvdd.n2242 dvdd.n2238 4.02033
R8609 dvdd.n2242 dvdd.n2241 4.02033
R8610 dvdd.n2351 dvdd.n2109 4.02033
R8611 dvdd.n2195 dvdd.n2190 4.02033
R8612 dvdd.n2195 dvdd.n2193 4.02033
R8613 dvdd.n2477 dvdd.n2476 4.02033
R8614 dvdd.n2547 dvdd.n2513 4.02033
R8615 dvdd.n2461 dvdd.n2460 4.02033
R8616 dvdd.n2418 dvdd.n2414 4.02033
R8617 dvdd.n2418 dvdd.n2417 4.02033
R8618 dvdd.n2633 dvdd.n2382 4.02033
R8619 dvdd.n2588 dvdd.n2583 4.02033
R8620 dvdd.n2588 dvdd.n2586 4.02033
R8621 dvdd.n818 dvdd.n815 3.91436
R8622 dvdd.n886 dvdd.n885 3.86515
R8623 dvdd.n2760 dvdd 3.85769
R8624 dvdd.n432 dvdd.n363 3.78037
R8625 dvdd.n705 dvdd.n704 3.78037
R8626 dvdd.n491 dvdd.n480 3.76521
R8627 dvdd.n729 dvdd.n728 3.76521
R8628 dvdd.n1016 dvdd.n1014 3.76521
R8629 dvdd.n1171 dvdd.n1105 3.76521
R8630 dvdd.n1648 dvdd.n1647 3.76521
R8631 dvdd.n1891 dvdd.n1890 3.76521
R8632 dvdd.n1898 dvdd.n1896 3.76521
R8633 dvdd.n2333 dvdd.n2332 3.76521
R8634 dvdd.n2802 dvdd 3.73954
R8635 dvdd dvdd.n1 3.73954
R8636 dvdd.n448 dvdd.n447 3.70298
R8637 dvdd.n715 dvdd.n714 3.70298
R8638 dvdd.n363 dvdd.n362 3.69446
R8639 dvdd.n704 dvdd.n643 3.69446
R8640 dvdd.n1991 dvdd.n1990 3.68131
R8641 dvdd.n2484 dvdd.n2395 3.66983
R8642 dvdd.n1363 dvdd.n1340 3.65764
R8643 dvdd.n1962 dvdd.n1961 3.65764
R8644 dvdd.n441 dvdd.n360 3.59719
R8645 dvdd.n501 dvdd.n472 3.55606
R8646 dvdd.n1588 dvdd.n1587 3.55606
R8647 dvdd.n234 dvdd.n232 3.50526
R8648 dvdd.n296 dvdd.n295 3.50526
R8649 dvdd.n152 dvdd.n91 3.50526
R8650 dvdd.n167 dvdd.n166 3.50526
R8651 dvdd.n2337 dvdd.n2336 3.50526
R8652 dvdd.n699 dvdd.n698 3.47425
R8653 dvdd.n1862 dvdd.n1828 3.47425
R8654 dvdd.n1863 dvdd.n1862 3.47425
R8655 dvdd.n2434 dvdd.n2409 3.47425
R8656 dvdd.n2435 dvdd.n2434 3.47425
R8657 dvdd.n2436 dvdd.n2435 3.47425
R8658 dvdd.n204 dvdd.n72 3.43925
R8659 dvdd.n327 dvdd.n326 3.43925
R8660 dvdd.n345 dvdd.n329 3.43925
R8661 dvdd.n610 dvdd.n609 3.43925
R8662 dvdd.n900 dvdd.n612 3.43925
R8663 dvdd.n911 dvdd.n910 3.43925
R8664 dvdd.n1191 dvdd.n913 3.43925
R8665 dvdd.n1200 dvdd.n1199 3.43925
R8666 dvdd.n1475 dvdd.n1202 3.43925
R8667 dvdd.n1484 dvdd.n1483 3.43925
R8668 dvdd.n1774 dvdd.n1486 3.43925
R8669 dvdd.n1785 dvdd.n1784 3.43925
R8670 dvdd.n1804 dvdd.n1787 3.43925
R8671 dvdd.n2087 dvdd.n2086 3.43925
R8672 dvdd.n2101 dvdd.n2089 3.43925
R8673 dvdd.n2357 dvdd.n2356 3.43925
R8674 dvdd.n2376 dvdd.n2359 3.43925
R8675 dvdd.n2645 dvdd.n2644 3.43925
R8676 dvdd.n75 dvdd.n73 3.4105
R8677 dvdd.n201 dvdd.n200 3.4105
R8678 dvdd.n332 dvdd.n330 3.4105
R8679 dvdd.n342 dvdd.n341 3.4105
R8680 dvdd.n615 dvdd.n613 3.4105
R8681 dvdd.n898 dvdd.n897 3.4105
R8682 dvdd.n916 dvdd.n914 3.4105
R8683 dvdd.n1189 dvdd.n1188 3.4105
R8684 dvdd.n1205 dvdd.n1203 3.4105
R8685 dvdd.n1473 dvdd.n1472 3.4105
R8686 dvdd.n1489 dvdd.n1487 3.4105
R8687 dvdd.n1772 dvdd.n1771 3.4105
R8688 dvdd.n1790 dvdd.n1788 3.4105
R8689 dvdd.n1801 dvdd.n1800 3.4105
R8690 dvdd.n2092 dvdd.n2090 3.4105
R8691 dvdd.n2099 dvdd.n2098 3.4105
R8692 dvdd.n2362 dvdd.n2360 3.4105
R8693 dvdd.n2373 dvdd.n2372 3.4105
R8694 dvdd.n1890 dvdd.n1817 3.38874
R8695 dvdd.n1850 dvdd.n1849 3.38562
R8696 dvdd.n2275 dvdd.n2274 3.37141
R8697 dvdd.n3141 dvdd.n3140 3.36414
R8698 dvdd.n3143 dvdd.n3141 3.36414
R8699 dvdd.n3147 dvdd.n3139 3.36414
R8700 dvdd.n3143 dvdd.n3139 3.36414
R8701 dvdd.n2968 dvdd.n2967 3.36211
R8702 dvdd dvdd.t536 3.35739
R8703 dvdd.t728 dvdd.t1413 3.35739
R8704 dvdd dvdd.t1415 3.35739
R8705 dvdd.t719 dvdd 3.35739
R8706 dvdd.t1263 dvdd.t120 3.35739
R8707 dvdd.t927 dvdd.t981 3.35739
R8708 dvdd.t847 dvdd.t17 3.35739
R8709 dvdd.t315 dvdd.t1643 3.35739
R8710 dvdd.t671 dvdd.t681 3.35739
R8711 dvdd.t628 dvdd.t733 3.35739
R8712 dvdd.n677 dvdd.n651 3.35288
R8713 dvdd.n2763 dvdd.n71 3.34378
R8714 dvdd.n2755 dvdd.n2652 3.34378
R8715 dvdd.n1865 dvdd.n1825 3.32144
R8716 dvdd.n700 dvdd.n699 3.2477
R8717 dvdd.n1857 dvdd.n1828 3.2477
R8718 dvdd.n1864 dvdd.n1863 3.2477
R8719 dvdd.n2427 dvdd.n2426 3.2477
R8720 dvdd.n2436 dvdd.n2407 3.2477
R8721 dvdd.n1298 dvdd.n1297 3.17405
R8722 dvdd.n2061 dvdd.n2060 3.17405
R8723 dvdd.n142 dvdd.n95 3.16454
R8724 dvdd.n1149 dvdd.n1148 3.14971
R8725 dvdd.n2934 dvdd.n2930 3.13609
R8726 dvdd.n2935 dvdd.n2934 3.13609
R8727 dvdd.n2939 dvdd.n2938 3.13609
R8728 dvdd.n2938 dvdd.n2937 3.13609
R8729 dvdd.n2143 dvdd.n2142 3.12116
R8730 dvdd.n2647 dvdd.n2 3.09532
R8731 dvdd.n2043 dvdd.n2042 3.06827
R8732 dvdd.n2269 dvdd.n2268 3.06827
R8733 dvdd.n384 dvdd.n383 3.05586
R8734 dvdd.n663 dvdd.n659 3.05586
R8735 dvdd.n961 dvdd.n960 3.05586
R8736 dvdd.n1264 dvdd.n1263 3.05586
R8737 dvdd.n1551 dvdd.n1547 3.05586
R8738 dvdd.n1840 dvdd.n1839 3.05586
R8739 dvdd.n2243 dvdd.n2242 3.05586
R8740 dvdd.n2419 dvdd.n2418 3.05586
R8741 dvdd.n2164 dvdd.n2148 3.05371
R8742 dvdd.n554 dvdd.n553 3.04861
R8743 dvdd.n843 dvdd.n842 3.04861
R8744 dvdd.n864 dvdd.n828 3.04861
R8745 dvdd.n1130 dvdd.n1129 3.04861
R8746 dvdd.n1421 dvdd.n1420 3.04861
R8747 dvdd.n1714 dvdd.n1713 3.04861
R8748 dvdd.n2025 dvdd.n2024 3.04861
R8749 dvdd.n2065 dvdd.n1998 3.04861
R8750 dvdd.n2195 dvdd.n2194 3.04861
R8751 dvdd.n2351 dvdd.n2106 3.04861
R8752 dvdd.n2588 dvdd.n2587 3.04861
R8753 dvdd.n2223 dvdd.n2173 3.04861
R8754 dvdd.n2462 dvdd.n2461 3.04861
R8755 dvdd.n2478 dvdd.n2477 3.04861
R8756 dvdd.n3101 dvdd.n3096 3.04784
R8757 dvdd.n1635 dvdd.n1633 3.03555
R8758 dvdd.n392 dvdd.n374 3.01588
R8759 dvdd.n418 dvdd.n417 3.01588
R8760 dvdd.n423 dvdd.n422 3.01588
R8761 dvdd.n569 dvdd.n542 3.01588
R8762 dvdd.n858 dvdd.n831 3.01588
R8763 dvdd.n2251 dvdd.n2233 3.01588
R8764 dvdd.n2303 dvdd.n2130 3.01588
R8765 dvdd.n2280 dvdd.n2137 3.01588
R8766 dvdd.n2178 dvdd.n2176 3.01588
R8767 dvdd.n1453 dvdd.n1452 3.01226
R8768 dvdd.n1583 dvdd.n1525 2.99733
R8769 dvdd.n2156 dvdd.n2154 2.99733
R8770 dvdd.n411 dvdd.n407 2.96248
R8771 dvdd.n2825 dvdd.n2820 2.95435
R8772 dvdd.n2853 dvdd.n2810 2.95435
R8773 dvdd.n2766 dvdd 2.9391
R8774 dvdd.n2770 dvdd 2.9391
R8775 dvdd.n2774 dvdd 2.9391
R8776 dvdd.n2778 dvdd 2.9391
R8777 dvdd.n2782 dvdd 2.9391
R8778 dvdd.n2786 dvdd 2.9391
R8779 dvdd.n2790 dvdd 2.9391
R8780 dvdd.n2794 dvdd 2.9391
R8781 dvdd.n2798 dvdd 2.9391
R8782 dvdd dvdd.n2748 2.9391
R8783 dvdd dvdd.n2744 2.9391
R8784 dvdd dvdd.n2740 2.9391
R8785 dvdd dvdd.n2736 2.9391
R8786 dvdd dvdd.n2732 2.9391
R8787 dvdd dvdd.n2728 2.9391
R8788 dvdd dvdd.n2724 2.9391
R8789 dvdd dvdd.n2720 2.9391
R8790 dvdd dvdd.n2752 2.9369
R8791 dvdd.n2951 dvdd.n2945 2.90005
R8792 dvdd.n1531 dvdd.n1527 2.87861
R8793 dvdd.n2352 dvdd.n2104 2.87861
R8794 dvdd.n2394 dvdd.n2392 2.8165
R8795 dvdd.n880 dvdd.n818 2.80769
R8796 dvdd.n3108 dvdd.n3103 2.80353
R8797 dvdd.n3109 dvdd.n3108 2.80353
R8798 dvdd.n3113 dvdd.n3112 2.80353
R8799 dvdd.n3112 dvdd.n3111 2.80353
R8800 dvdd.n146 dvdd.n145 2.76904
R8801 dvdd.n969 dvdd.n968 2.74336
R8802 dvdd.n2606 dvdd.n2573 2.74336
R8803 dvdd.n395 dvdd.n374 2.64665
R8804 dvdd.n417 dvdd.n367 2.64665
R8805 dvdd.n424 dvdd.n423 2.64665
R8806 dvdd.n566 dvdd.n542 2.64665
R8807 dvdd.n855 dvdd.n831 2.64665
R8808 dvdd.n2254 dvdd.n2233 2.64665
R8809 dvdd.n2306 dvdd.n2130 2.64665
R8810 dvdd.n2283 dvdd.n2137 2.64665
R8811 dvdd.n2220 dvdd.n2219 2.64665
R8812 dvdd.n2219 dvdd.n2218 2.64665
R8813 dvdd.n2213 dvdd.n2178 2.64665
R8814 dvdd.n2228 dvdd.t737 2.63714
R8815 dvdd.n1563 dvdd.n1539 2.63579
R8816 dvdd.n1557 dvdd.n1554 2.63579
R8817 dvdd.n2493 dvdd.n2389 2.63579
R8818 dvdd.n379 dvdd.n377 2.63539
R8819 dvdd.n382 dvdd.n380 2.63539
R8820 dvdd.n537 dvdd.n535 2.63539
R8821 dvdd.n549 dvdd.n547 2.63539
R8822 dvdd.n552 dvdd.n550 2.63539
R8823 dvdd.n658 dvdd.n656 2.63539
R8824 dvdd.n662 dvdd.n660 2.63539
R8825 dvdd.n827 dvdd.n825 2.63539
R8826 dvdd.n838 dvdd.n836 2.63539
R8827 dvdd.n841 dvdd.n839 2.63539
R8828 dvdd.n956 dvdd.n954 2.63539
R8829 dvdd.n959 dvdd.n957 2.63539
R8830 dvdd.n1125 dvdd.n1123 2.63539
R8831 dvdd.n1128 dvdd.n1126 2.63539
R8832 dvdd.n1259 dvdd.n1257 2.63539
R8833 dvdd.n1262 dvdd.n1260 2.63539
R8834 dvdd.n1416 dvdd.n1414 2.63539
R8835 dvdd.n1419 dvdd.n1417 2.63539
R8836 dvdd.n1546 dvdd.n1544 2.63539
R8837 dvdd.n1550 dvdd.n1548 2.63539
R8838 dvdd.n1709 dvdd.n1707 2.63539
R8839 dvdd.n1712 dvdd.n1710 2.63539
R8840 dvdd.n1835 dvdd.n1833 2.63539
R8841 dvdd.n1838 dvdd.n1836 2.63539
R8842 dvdd.n1997 dvdd.n1995 2.63539
R8843 dvdd.n2020 dvdd.n2018 2.63539
R8844 dvdd.n2023 dvdd.n2021 2.63539
R8845 dvdd.n2142 dvdd.n2140 2.63539
R8846 dvdd.n2238 dvdd.n2236 2.63539
R8847 dvdd.n2241 dvdd.n2239 2.63539
R8848 dvdd.n2109 dvdd.n2107 2.63539
R8849 dvdd.n2190 dvdd.n2188 2.63539
R8850 dvdd.n2193 dvdd.n2191 2.63539
R8851 dvdd.n2476 dvdd.n2474 2.63539
R8852 dvdd.n2513 dvdd.n2511 2.63539
R8853 dvdd.n2382 dvdd.n2380 2.63539
R8854 dvdd.n2460 dvdd.n2458 2.63539
R8855 dvdd.n2414 dvdd.n2412 2.63539
R8856 dvdd.n2417 dvdd.n2415 2.63539
R8857 dvdd.n2583 dvdd.n2581 2.63539
R8858 dvdd.n2586 dvdd.n2584 2.63539
R8859 dvdd.n2891 dvdd.n2886 2.63064
R8860 dvdd.n2919 dvdd.n2876 2.63064
R8861 dvdd.n2172 dvdd.n2171 2.62644
R8862 dvdd.n1526 dvdd.n1525 2.61352
R8863 dvdd.n2154 dvdd.n2153 2.61352
R8864 dvdd.n3045 dvdd.n3040 2.59509
R8865 dvdd.n3073 dvdd.n3030 2.59509
R8866 dvdd.n2988 dvdd.n2983 2.59509
R8867 dvdd.n3016 dvdd.n2973 2.59509
R8868 dvdd.n1374 dvdd.n1373 2.5605
R8869 dvdd.n2842 dvdd.n2814 2.5605
R8870 dvdd.t737 dvdd.t668 2.53573
R8871 dvdd.n2969 dvdd.n2968 2.52884
R8872 dvdd.n3101 dvdd.n0 2.49068
R8873 dvdd.n1153 dvdd.n1115 2.48939
R8874 dvdd.n668 dvdd.n667 2.4386
R8875 dvdd.n1156 dvdd.n1155 2.4386
R8876 dvdd.n1667 dvdd.n1633 2.37576
R8877 dvdd.n381 dvdd.n380 2.37495
R8878 dvdd.n378 dvdd.n377 2.37495
R8879 dvdd.n536 dvdd.n535 2.37495
R8880 dvdd.n551 dvdd.n550 2.37495
R8881 dvdd.n548 dvdd.n547 2.37495
R8882 dvdd.n661 dvdd.n660 2.37495
R8883 dvdd.n657 dvdd.n656 2.37495
R8884 dvdd.n826 dvdd.n825 2.37495
R8885 dvdd.n840 dvdd.n839 2.37495
R8886 dvdd.n837 dvdd.n836 2.37495
R8887 dvdd.n958 dvdd.n957 2.37495
R8888 dvdd.n955 dvdd.n954 2.37495
R8889 dvdd.n1127 dvdd.n1126 2.37495
R8890 dvdd.n1124 dvdd.n1123 2.37495
R8891 dvdd.n1261 dvdd.n1260 2.37495
R8892 dvdd.n1258 dvdd.n1257 2.37495
R8893 dvdd.n1418 dvdd.n1417 2.37495
R8894 dvdd.n1415 dvdd.n1414 2.37495
R8895 dvdd.n1549 dvdd.n1548 2.37495
R8896 dvdd.n1545 dvdd.n1544 2.37495
R8897 dvdd.n1711 dvdd.n1710 2.37495
R8898 dvdd.n1708 dvdd.n1707 2.37495
R8899 dvdd.n1837 dvdd.n1836 2.37495
R8900 dvdd.n1834 dvdd.n1833 2.37495
R8901 dvdd.n1996 dvdd.n1995 2.37495
R8902 dvdd.n2022 dvdd.n2021 2.37495
R8903 dvdd.n2019 dvdd.n2018 2.37495
R8904 dvdd.n2141 dvdd.n2140 2.37495
R8905 dvdd.n2240 dvdd.n2239 2.37495
R8906 dvdd.n2237 dvdd.n2236 2.37495
R8907 dvdd.n2108 dvdd.n2107 2.37495
R8908 dvdd.n2192 dvdd.n2191 2.37495
R8909 dvdd.n2189 dvdd.n2188 2.37495
R8910 dvdd.n2475 dvdd.n2474 2.37495
R8911 dvdd.n2512 dvdd.n2511 2.37495
R8912 dvdd.n2459 dvdd.n2458 2.37495
R8913 dvdd.n2416 dvdd.n2415 2.37495
R8914 dvdd.n2413 dvdd.n2412 2.37495
R8915 dvdd.n2381 dvdd.n2380 2.37495
R8916 dvdd.n2585 dvdd.n2584 2.37495
R8917 dvdd.n2582 dvdd.n2581 2.37495
R8918 dvdd.n2854 dvdd.n2809 2.36358
R8919 dvdd.n2864 dvdd.n2863 2.36358
R8920 dvdd.n211 dvdd.n210 2.33701
R8921 dvdd.n505 dvdd.n504 2.33701
R8922 dvdd.n670 dvdd.n669 2.33701
R8923 dvdd.n671 dvdd.n670 2.33701
R8924 dvdd.n891 dvdd.n890 2.33701
R8925 dvdd.n966 dvdd.n965 2.33701
R8926 dvdd.n1031 dvdd.n931 2.33701
R8927 dvdd.n1921 dvdd.n1920 2.33701
R8928 dvdd.n1985 dvdd.n1928 2.33701
R8929 dvdd.n2075 dvdd.n2074 2.33701
R8930 dvdd.n689 dvdd.n687 2.32777
R8931 dvdd.n865 dvdd.n864 2.32777
R8932 dvdd.n2175 dvdd.n2173 2.28432
R8933 dvdd.n2168 dvdd.n2167 2.28407
R8934 dvdd.n2169 dvdd.n2168 2.28407
R8935 dvdd.n2910 dvdd.n2880 2.27995
R8936 dvdd.n2477 dvdd.n2473 2.27488
R8937 dvdd.n2461 dvdd.n2401 2.27488
R8938 dvdd.n515 dvdd.n466 2.25932
R8939 dvdd.n979 dvdd.n976 2.25932
R8940 dvdd.n1465 dvdd.n1464 2.25932
R8941 dvdd.n1577 dvdd.n1576 2.25932
R8942 dvdd.n1976 dvdd.n1975 2.25932
R8943 dvdd.n3064 dvdd.n3034 2.24915
R8944 dvdd.n3007 dvdd.n2977 2.24915
R8945 dvdd.n669 dvdd.n668 2.23542
R8946 dvdd.n1155 dvdd.n1154 2.23542
R8947 dvdd.n1370 dvdd.n1369 2.19479
R8948 dvdd.n1952 dvdd.n1951 2.19479
R8949 dvdd.n2647 dvdd 2.19219
R8950 dvdd.n1150 dvdd.n1115 2.18463
R8951 dvdd.n2392 dvdd.n2391 2.1843
R8952 dvdd.n3096 dvdd 2.16978
R8953 dvdd.n94 dvdd.n92 2.1578
R8954 dvdd.n2921 dvdd.n2920 2.10461
R8955 dvdd.n2932 dvdd.n2929 2.10277
R8956 dvdd.n2936 dvdd.n2932 2.10277
R8957 dvdd.n2940 dvdd.n2931 2.10277
R8958 dvdd.n2933 dvdd.n2931 2.10277
R8959 dvdd.n3075 dvdd.n3074 2.07618
R8960 dvdd.n3018 dvdd.n3017 2.07618
R8961 dvdd.n2166 dvdd.n2148 2.07374
R8962 dvdd.n2171 dvdd.n2170 2.07374
R8963 dvdd.n210 dvdd.n209 2.03225
R8964 dvdd.n506 dvdd.n505 2.03225
R8965 dvdd.n769 dvdd.n768 2.03225
R8966 dvdd.n892 dvdd.n891 2.03225
R8967 dvdd.n965 dvdd.n964 2.03225
R8968 dvdd.n1032 dvdd.n1031 2.03225
R8969 dvdd.n1928 dvdd.n1927 2.03225
R8970 dvdd.n2076 dvdd.n2075 2.03225
R8971 dvdd.n2323 dvdd.n2322 2.03225
R8972 dvdd.n873 dvdd.n872 2.01042
R8973 dvdd.n1297 dvdd.n1234 2.01042
R8974 dvdd.n1311 dvdd.n1310 2.01042
R8975 dvdd.n2049 dvdd.n2048 2.01042
R8976 dvdd.n2324 dvdd.n2323 1.98145
R8977 dvdd.n726 dvdd.n725 1.95345
R8978 dvdd.n2603 dvdd.n2573 1.93066
R8979 dvdd.n3094 dvdd.n3083 1.92238
R8980 dvdd.n446 dvdd.n445 1.90463
R8981 dvdd.n2297 dvdd.n2296 1.88325
R8982 dvdd.n604 dvdd.n603 1.88285
R8983 dvdd.n1134 dvdd.n1133 1.88285
R8984 dvdd.n2430 dvdd.n2429 1.85065
R8985 dvdd.n2428 dvdd.n2427 1.81289
R8986 dvdd.n2224 dvdd.n2168 1.76897
R8987 dvdd.n698 dvdd.n645 1.73737
R8988 dvdd.n2542 dvdd.n2541 1.70717
R8989 dvdd.n2802 dvdd.n1 1.69386
R8990 dvdd.n2646 dvdd.n2359 1.69188
R8991 dvdd.n2646 dvdd.n2645 1.69188
R8992 dvdd.n2358 dvdd.n2089 1.69188
R8993 dvdd.n2358 dvdd.n2357 1.69188
R8994 dvdd.n2088 dvdd.n1787 1.69188
R8995 dvdd.n2088 dvdd.n2087 1.69188
R8996 dvdd.n1786 dvdd.n1486 1.69188
R8997 dvdd.n1786 dvdd.n1785 1.69188
R8998 dvdd.n1485 dvdd.n1202 1.69188
R8999 dvdd.n1485 dvdd.n1484 1.69188
R9000 dvdd.n1201 dvdd.n913 1.69188
R9001 dvdd.n1201 dvdd.n1200 1.69188
R9002 dvdd.n912 dvdd.n612 1.69188
R9003 dvdd.n912 dvdd.n911 1.69188
R9004 dvdd.n611 dvdd.n329 1.69188
R9005 dvdd.n611 dvdd.n610 1.69188
R9006 dvdd.n328 dvdd.n72 1.69188
R9007 dvdd.n328 dvdd.n327 1.69188
R9008 dvdd.t1278 dvdd.t803 1.67895
R9009 dvdd.n813 dvdd.t482 1.67895
R9010 dvdd.t8 dvdd.t1077 1.67895
R9011 dvdd dvdd.t1239 1.67895
R9012 dvdd.t1107 dvdd.t1505 1.67895
R9013 dvdd.t76 dvdd.t504 1.67895
R9014 dvdd.t1056 dvdd.t1387 1.67895
R9015 dvdd.t250 dvdd.t1382 1.67895
R9016 dvdd.t1245 dvdd.t867 1.67895
R9017 dvdd.t164 dvdd.t1485 1.67895
R9018 dvdd.n2430 dvdd.n2428 1.66186
R9019 dvdd.n2757 dvdd 1.653
R9020 dvdd.n2761 dvdd 1.64081
R9021 dvdd.n970 dvdd.n969 1.6259
R9022 dvdd.n2429 dvdd.n2409 1.6241
R9023 dvdd.t325 dvdd.n2146 1.62304
R9024 dvdd.n2298 dvdd.n2297 1.62136
R9025 dvdd.n770 dvdd.n769 1.52431
R9026 dvdd.n1148 dvdd.n1147 1.52431
R9027 dvdd.t1522 dvdd.t618 1.52164
R9028 dvdd.n694 dvdd.n645 1.51082
R9029 dvdd.n463 dvdd.n462 1.50638
R9030 dvdd.n484 dvdd.n483 1.50638
R9031 dvdd.n483 dvdd.n336 1.50638
R9032 dvdd.n992 dvdd.n943 1.50638
R9033 dvdd.n1089 dvdd.n1088 1.50638
R9034 dvdd.n1276 dvdd.n1249 1.50638
R9035 dvdd.n1455 dvdd.n1391 1.50638
R9036 dvdd.n1678 dvdd.n1626 1.50638
R9037 dvdd.n1599 dvdd.n1514 1.50638
R9038 dvdd.n1879 dvdd.n1823 1.50638
R9039 dvdd.n2531 dvdd.n2530 1.50638
R9040 dvdd.n1034 dvdd.n1028 1.47352
R9041 dvdd.n1043 dvdd.n930 1.47352
R9042 dvdd.n499 dvdd.n498 1.46742
R9043 dvdd.n1368 dvdd.n1367 1.46336
R9044 dvdd.n1358 dvdd.n1357 1.46336
R9045 dvdd.n2146 dvdd.t522 1.42023
R9046 dvdd.t618 dvdd.n2147 1.42023
R9047 dvdd.n453 dvdd.n452 1.37571
R9048 dvdd.n717 dvdd.n639 1.37571
R9049 dvdd.n1920 dvdd.n1919 1.32113
R9050 dvdd.t70 dvdd.t1556 1.31882
R9051 dvdd.t668 dvdd.t1522 1.31882
R9052 dvdd.n2969 dvdd.n2943 1.26417
R9053 dvdd.n1527 dvdd.n1525 1.2502
R9054 dvdd.n2154 dvdd.n2104 1.2502
R9055 dvdd.n2909 dvdd.n2907 1.2279
R9056 dvdd.n2862 dvdd.n2806 1.18204
R9057 dvdd.n1656 dvdd.n1638 1.15949
R9058 dvdd.n3095 dvdd.n2 1.15094
R9059 dvdd.n787 dvdd.n786 1.12991
R9060 dvdd.n904 dvdd.n903 1.12991
R9061 dvdd.n1095 dvdd.n1052 1.12991
R9062 dvdd.n1174 dvdd.n1173 1.12991
R9063 dvdd.n1980 dvdd.n1931 1.12991
R9064 dvdd.n504 dvdd.n472 1.11796
R9065 dvdd.n2539 dvdd.n2521 1.07613
R9066 dvdd.n3047 dvdd.n3041 1.06234
R9067 dvdd.n2990 dvdd.n2984 1.06234
R9068 dvdd.n2893 dvdd.n2887 1.05227
R9069 dvdd.n3149 dvdd.n3116 1.04961
R9070 dvdd.n3063 dvdd.n3061 1.03834
R9071 dvdd.n3006 dvdd.n3004 1.03834
R9072 dvdd.n678 dvdd.n677 1.01637
R9073 dvdd.n2167 dvdd.n2148 0.992049
R9074 dvdd.n2171 dvdd.n2169 0.992049
R9075 dvdd.n2827 dvdd.n2821 0.968765
R9076 dvdd.n2967 dvdd.n2945 0.955857
R9077 dvdd.n3155 dvdd.n1 0.951672
R9078 dvdd.n146 dvdd.n94 0.935332
R9079 dvdd.n2757 dvdd.n2756 0.910588
R9080 dvdd.n232 dvdd.n230 0.863992
R9081 dvdd.n295 dvdd.n294 0.863992
R9082 dvdd.n91 dvdd.n90 0.863992
R9083 dvdd.n166 dvdd.n165 0.863992
R9084 dvdd.n2336 dvdd.n2335 0.863992
R9085 dvdd.n3026 dvdd.n2969 0.836438
R9086 dvdd.n2762 dvdd.n2761 0.83164
R9087 dvdd.n780 dvdd.n770 0.813198
R9088 dvdd.n1587 dvdd.n1586 0.813198
R9089 dvdd.t1556 dvdd.t1027 0.811772
R9090 dvdd.n3083 dvdd.n3026 0.808117
R9091 dvdd.n3123 dvdd.n3122 0.787085
R9092 dvdd.n1990 dvdd.n1988 0.783573
R9093 dvdd.n328 dvdd.n2 0.782766
R9094 dvdd.n2633 dvdd.n2557 0.775896
R9095 dvdd.n510 dvdd.n471 0.753441
R9096 dvdd.n493 dvdd.n492 0.753441
R9097 dvdd.n605 dvdd.n604 0.753441
R9098 dvdd.n589 dvdd.n588 0.753441
R9099 dvdd.n794 dvdd.n793 0.753441
R9100 dvdd.n1080 dvdd.n1079 0.753441
R9101 dvdd.n1135 dvdd.n1120 0.753441
R9102 dvdd.n1401 dvdd.n1398 0.753441
R9103 dvdd.n1557 dvdd.n1556 0.753441
R9104 dvdd.n1764 dvdd.n1499 0.753441
R9105 dvdd.n1617 dvdd.n1507 0.753441
R9106 dvdd.n1595 dvdd.n1514 0.753441
R9107 dvdd.n1748 dvdd.n1747 0.753441
R9108 dvdd.n1720 dvdd.n1719 0.753441
R9109 dvdd.n1882 dvdd.n1881 0.753441
R9110 dvdd.n1907 dvdd.n1906 0.753441
R9111 dvdd.n2635 dvdd.n2379 0.753441
R9112 dvdd.n2483 dvdd.n2482 0.740996
R9113 dvdd.n2466 dvdd.n2400 0.740996
R9114 dvdd.n2455 dvdd.n2454 0.740996
R9115 dvdd.n750 dvdd.n749 0.731929
R9116 dvdd.n808 dvdd.n807 0.731929
R9117 dvdd.n1919 dvdd.n1918 0.711611
R9118 dvdd.t1027 dvdd.t522 0.710363
R9119 dvdd.n2952 dvdd.n2951 0.705857
R9120 dvdd.n2953 dvdd.n2952 0.705857
R9121 dvdd.n2959 dvdd.n2958 0.705857
R9122 dvdd.n2958 dvdd.n2957 0.705857
R9123 dvdd.n2957 dvdd.n2944 0.705857
R9124 dvdd.n2943 dvdd.n2872 0.691906
R9125 dvdd.n2077 dvdd.n1798 0.681097
R9126 dvdd.n1664 dvdd.n1635 0.660294
R9127 dvdd.n1664 dvdd.n1663 0.660294
R9128 dvdd.n2942 dvdd 0.645031
R9129 dvdd.n1531 dvdd.n1530 0.644287
R9130 dvdd.n257 dvdd.n223 0.635211
R9131 dvdd.n238 dvdd.n229 0.635211
R9132 dvdd.n276 dvdd.n275 0.635211
R9133 dvdd.n258 dvdd.n222 0.635211
R9134 dvdd.n301 dvdd.n300 0.635211
R9135 dvdd.n321 dvdd.n319 0.635211
R9136 dvdd.n100 dvdd.n98 0.635211
R9137 dvdd.n114 dvdd.n105 0.635211
R9138 dvdd.n172 dvdd.n162 0.635211
R9139 dvdd.n191 dvdd.n156 0.635211
R9140 dvdd.n456 dvdd.n455 0.635211
R9141 dvdd.n707 dvdd.n706 0.635211
R9142 dvdd.n725 dvdd.n636 0.635211
R9143 dvdd.n682 dvdd.n650 0.635211
R9144 dvdd.n880 dvdd.n879 0.635211
R9145 dvdd.n1292 dvdd.n1236 0.635211
R9146 dvdd.n1314 dvdd.n1229 0.635211
R9147 dvdd.n1844 dvdd.n1843 0.635211
R9148 dvdd.n2063 dvdd.n2062 0.635211
R9149 dvdd.n2004 dvdd.n2003 0.635211
R9150 dvdd.n2312 dvdd.n2127 0.635211
R9151 dvdd.n2318 dvdd.n2317 0.635211
R9152 dvdd.n2202 dvdd.n2183 0.635211
R9153 dvdd.n2468 dvdd.n2467 0.635211
R9154 dvdd.n2422 dvdd.n2411 0.635211
R9155 dvdd.n2942 dvdd.n2941 0.633614
R9156 dvdd.n2849 dvdd.n2848 0.591269
R9157 dvdd.n145 dvdd.n95 0.539826
R9158 dvdd.n2960 dvdd.n2953 0.529518
R9159 dvdd.n410 dvdd.n369 0.529426
R9160 dvdd.n2008 dvdd.n2007 0.529426
R9161 dvdd.n2915 dvdd.n2914 0.526527
R9162 dvdd.n3069 dvdd.n3068 0.519419
R9163 dvdd.n3012 dvdd.n3011 0.519419
R9164 dvdd.n2941 dvdd.n2929 0.517903
R9165 dvdd.n3122 dvdd.n3121 0.514219
R9166 dvdd.n3135 dvdd.n3134 0.492878
R9167 dvdd.n3120 dvdd.n3098 0.482207
R9168 dvdd.n3131 dvdd.n3123 0.482207
R9169 dvdd.n3132 dvdd.n3131 0.482207
R9170 dvdd.n3133 dvdd.n3132 0.482207
R9171 dvdd.n3106 dvdd.n3105 0.448442
R9172 dvdd.n3107 dvdd.n3106 0.448442
R9173 dvdd.n3114 dvdd.n3104 0.448442
R9174 dvdd.n3110 dvdd.n3104 0.448442
R9175 dvdd.n3151 dvdd.n3098 0.447146
R9176 dvdd.n708 dvdd.n641 0.42364
R9177 dvdd.n3136 dvdd.n3135 0.419707
R9178 dvdd.n3134 dvdd.n3133 0.386171
R9179 dvdd.n498 dvdd.n497 0.384032
R9180 dvdd.n732 dvdd.n729 0.376971
R9181 dvdd.n1092 dvdd.n1055 0.376971
R9182 dvdd.n1081 dvdd.n1080 0.376971
R9183 dvdd.n1180 dvdd.n925 0.376971
R9184 dvdd.n1563 dvdd.n1562 0.376971
R9185 dvdd.n1874 dvdd.n1873 0.376971
R9186 dvdd.n2345 dvdd.n2113 0.376971
R9187 dvdd.n2628 dvdd.n2561 0.376971
R9188 dvdd.n2627 dvdd.n2626 0.376971
R9189 dvdd.n3151 dvdd.n3150 0.372451
R9190 dvdd.n387 dvdd.n376 0.369731
R9191 dvdd.n406 dvdd.n370 0.369731
R9192 dvdd.n416 dvdd.n415 0.369731
R9193 dvdd.n433 dvdd.n431 0.369731
R9194 dvdd.n574 dvdd.n540 0.369731
R9195 dvdd.n555 dvdd.n546 0.369731
R9196 dvdd.n863 dvdd.n829 0.369731
R9197 dvdd.n844 dvdd.n835 0.369731
R9198 dvdd.n2246 dvdd.n2235 0.369731
R9199 dvdd.n2262 dvdd.n2144 0.369731
R9200 dvdd.n2298 dvdd.n2132 0.369731
R9201 dvdd.n2311 dvdd.n2128 0.369731
R9202 dvdd.n2291 dvdd.n2290 0.369731
R9203 dvdd.n2296 dvdd.n2133 0.369731
R9204 dvdd.n2275 dvdd.n2139 0.369731
R9205 dvdd.n2285 dvdd.n2135 0.369731
R9206 dvdd.n2221 dvdd.n2220 0.369731
R9207 dvdd.n2207 dvdd.n2180 0.369731
R9208 dvdd.n2441 dvdd.n2440 0.369731
R9209 dvdd.n2445 dvdd.n2405 0.369731
R9210 dvdd.n1361 dvdd.n1342 0.366214
R9211 dvdd.n3121 dvdd.n3120 0.361781
R9212 dvdd.n2325 dvdd.n2324 0.356056
R9213 dvdd.n2968 dvdd.n2944 0.346482
R9214 dvdd.n2545 dvdd.n2517 0.323189
R9215 dvdd.n2616 dvdd.n2615 0.323189
R9216 dvdd.n2961 dvdd.n2960 0.3105
R9217 dvdd.n2967 dvdd.n2966 0.3105
R9218 dvdd.n3137 dvdd.n3123 0.307565
R9219 dvdd.n237 dvdd.n230 0.305262
R9220 dvdd.n209 dvdd.n208 0.305262
R9221 dvdd.n212 dvdd.n195 0.305262
R9222 dvdd.n294 dvdd.n293 0.305262
R9223 dvdd.n299 dvdd.n83 0.305262
R9224 dvdd.n135 dvdd.n134 0.305262
R9225 dvdd.n90 dvdd.n88 0.305262
R9226 dvdd.n151 dvdd.n150 0.305262
R9227 dvdd.n165 dvdd.n163 0.305262
R9228 dvdd.n507 dvdd.n506 0.305262
R9229 dvdd.n500 dvdd.n499 0.305262
R9230 dvdd.n681 dvdd.n651 0.305262
R9231 dvdd.n664 dvdd.n655 0.305262
R9232 dvdd.n768 dvdd.n765 0.305262
R9233 dvdd.n893 dvdd.n892 0.305262
R9234 dvdd.n886 dvdd.n624 0.305262
R9235 dvdd.n964 dvdd.n963 0.305262
R9236 dvdd.n968 dvdd.n952 0.305262
R9237 dvdd.n1159 dvdd.n1112 0.305262
R9238 dvdd.n1144 dvdd.n1117 0.305262
R9239 dvdd.n1602 dvdd.n1601 0.305262
R9240 dvdd.n1586 dvdd.n1523 0.305262
R9241 dvdd.n1918 dvdd.n1917 0.305262
R9242 dvdd.n1922 dvdd.n1808 0.305262
R9243 dvdd.n1988 dvdd.n1927 0.305262
R9244 dvdd.n2077 dvdd.n2076 0.305262
R9245 dvdd.n2070 dvdd.n2069 0.305262
R9246 dvdd.n2335 dvdd.n2334 0.305262
R9247 dvdd.n2340 dvdd.n2116 0.305262
R9248 dvdd.n2322 dvdd.n2321 0.305262
R9249 dvdd.n2326 dvdd.n2121 0.305262
R9250 dvdd.n2570 dvdd.n2567 0.305262
R9251 dvdd.n2602 dvdd.n2601 0.305262
R9252 dvdd.n2599 dvdd.n2576 0.305262
R9253 dvdd.n2590 dvdd.n2589 0.305262
R9254 dvdd dvdd.n2224 0.2951
R9255 dvdd.n3148 dvdd.n3137 0.272821
R9256 dvdd.n1659 dvdd.n1636 0.264418
R9257 dvdd.n2224 dvdd 0.256072
R9258 dvdd.n777 dvdd.n776 0.254468
R9259 dvdd.n2571 dvdd.n2570 0.254468
R9260 dvdd.n3150 dvdd.n3149 0.252732
R9261 dvdd.n732 dvdd.n731 0.25148
R9262 dvdd.n803 dvdd.n801 0.246654
R9263 dvdd.n695 dvdd.n694 0.227049
R9264 dvdd.n701 dvdd.n700 0.227049
R9265 dvdd.n1858 dvdd.n1857 0.227049
R9266 dvdd.n1865 dvdd.n1864 0.227049
R9267 dvdd.n2426 dvdd.n2425 0.227049
R9268 dvdd.n2439 dvdd.n2407 0.227049
R9269 dvdd.n553 dvdd 0.217591
R9270 dvdd.n842 dvdd 0.217591
R9271 dvdd.n149 dvdd.n92 0.21623
R9272 dvdd.n824 dvdd.n822 0.21207
R9273 dvdd.n2399 dvdd.n2398 0.21207
R9274 dvdd.n2446 dvdd.n2404 0.21207
R9275 dvdd.n3135 dvdd.n3126 0.206229
R9276 dvdd.n2759 dvdd.n2758 0.204363
R9277 dvdd.n1600 dvdd.n1512 0.203675
R9278 dvdd.n1608 dvdd.n1607 0.203675
R9279 dvdd.n1610 dvdd.n1609 0.203675
R9280 dvdd.n1981 dvdd.n1930 0.203675
R9281 dvdd.n2071 dvdd.n1806 0.203675
R9282 dvdd.n1071 dvdd.n1064 0.180304
R9283 dvdd.n1241 dvdd.n1239 0.180304
R9284 dvdd.n2507 dvdd.n2503 0.180304
R9285 dvdd.n1582 dvdd.n1581 0.180304
R9286 dvdd dvdd.n1130 0.17983
R9287 dvdd dvdd.n1421 0.17983
R9288 dvdd.n1713 dvdd 0.17983
R9289 dvdd.n2024 dvdd 0.17983
R9290 dvdd.n2194 dvdd 0.17983
R9291 dvdd.n2587 dvdd 0.17983
R9292 dvdd dvdd.n2223 0.17983
R9293 dvdd.n2462 dvdd 0.17983
R9294 dvdd.n2478 dvdd 0.17983
R9295 dvdd.n828 dvdd 0.179485
R9296 dvdd dvdd.n2065 0.179485
R9297 dvdd dvdd.n2106 0.179485
R9298 dvdd.n3140 dvdd.n3099 0.179346
R9299 dvdd.n3148 dvdd.n3147 0.179346
R9300 dvdd.n2960 dvdd.n2959 0.176839
R9301 dvdd dvdd.n384 0.172576
R9302 dvdd.n659 dvdd 0.172576
R9303 dvdd dvdd.n961 0.172576
R9304 dvdd dvdd.n1264 0.172576
R9305 dvdd.n1547 dvdd 0.172576
R9306 dvdd dvdd.n1840 0.172576
R9307 dvdd dvdd.n2243 0.172576
R9308 dvdd dvdd.n2419 0.172576
R9309 dvdd.n611 dvdd.n328 0.1603
R9310 dvdd.n912 dvdd.n611 0.1603
R9311 dvdd.n1201 dvdd.n912 0.1603
R9312 dvdd.n1485 dvdd.n1201 0.1603
R9313 dvdd.n1786 dvdd.n1485 0.1603
R9314 dvdd.n2088 dvdd.n1786 0.1603
R9315 dvdd.n2358 dvdd.n2088 0.1603
R9316 dvdd.n2646 dvdd.n2358 0.1603
R9317 dvdd.n435 dvdd 0.158169
R9318 dvdd.n1581 dvdd 0.158169
R9319 dvdd.n1034 dvdd.n1033 0.152881
R9320 dvdd.n1033 dvdd.n1032 0.152881
R9321 dvdd.n1042 dvdd.n1039 0.152881
R9322 dvdd.n1043 dvdd.n1042 0.152881
R9323 dvdd.n3133 dvdd.n3128 0.152674
R9324 dvdd.n142 dvdd.n141 0.14432
R9325 dvdd dvdd.n828 0.14207
R9326 dvdd.n2065 dvdd 0.14207
R9327 dvdd.n2106 dvdd 0.14207
R9328 dvdd.n553 dvdd 0.141725
R9329 dvdd.n842 dvdd 0.141725
R9330 dvdd.n1130 dvdd 0.141725
R9331 dvdd.n1421 dvdd 0.141725
R9332 dvdd.n1713 dvdd 0.141725
R9333 dvdd.n2024 dvdd 0.141725
R9334 dvdd.n2223 dvdd 0.141725
R9335 dvdd.n2194 dvdd 0.141725
R9336 dvdd dvdd.n2462 0.141725
R9337 dvdd dvdd.n2478 0.141725
R9338 dvdd.n2587 dvdd 0.141725
R9339 dvdd.n2758 dvdd.n0 0.122113
R9340 dvdd.n3093 dvdd 0.121114
R9341 dvdd.n2765 dvdd 0.121114
R9342 dvdd.n2769 dvdd 0.121114
R9343 dvdd.n2773 dvdd 0.121114
R9344 dvdd.n2777 dvdd 0.121114
R9345 dvdd.n2781 dvdd 0.121114
R9346 dvdd.n2785 dvdd 0.121114
R9347 dvdd.n2789 dvdd 0.121114
R9348 dvdd.n2793 dvdd 0.121114
R9349 dvdd.n2797 dvdd 0.121114
R9350 dvdd.n2801 dvdd 0.121114
R9351 dvdd.n2753 dvdd 0.121114
R9352 dvdd.n2749 dvdd 0.121114
R9353 dvdd.n2745 dvdd 0.121114
R9354 dvdd.n2741 dvdd 0.121114
R9355 dvdd.n2737 dvdd 0.121114
R9356 dvdd.n2733 dvdd 0.121114
R9357 dvdd.n2729 dvdd 0.121114
R9358 dvdd.n2725 dvdd 0.121114
R9359 dvdd.n2721 dvdd 0.121114
R9360 dvdd.n2717 dvdd 0.121114
R9361 dvdd.n539 dvdd 0.120408
R9362 dvdd.n2510 dvdd 0.120408
R9363 dvdd.n2384 dvdd 0.120408
R9364 dvdd.n703 dvdd 0.120408
R9365 dvdd.n2487 dvdd 0.120408
R9366 dvdd.n169 dvdd.n168 0.120292
R9367 dvdd.n174 dvdd.n173 0.120292
R9368 dvdd.n174 dvdd.n161 0.120292
R9369 dvdd.n178 dvdd.n161 0.120292
R9370 dvdd.n179 dvdd.n178 0.120292
R9371 dvdd.n179 dvdd.n159 0.120292
R9372 dvdd.n183 dvdd.n159 0.120292
R9373 dvdd.n184 dvdd.n183 0.120292
R9374 dvdd.n185 dvdd.n184 0.120292
R9375 dvdd.n185 dvdd.n157 0.120292
R9376 dvdd.n189 dvdd.n157 0.120292
R9377 dvdd.n190 dvdd.n189 0.120292
R9378 dvdd.n154 dvdd.n153 0.120292
R9379 dvdd.n153 dvdd.n89 0.120292
R9380 dvdd.n148 dvdd.n147 0.120292
R9381 dvdd.n147 dvdd.n93 0.120292
R9382 dvdd.n140 dvdd.n93 0.120292
R9383 dvdd.n140 dvdd.n139 0.120292
R9384 dvdd.n139 dvdd.n138 0.120292
R9385 dvdd.n138 dvdd.n97 0.120292
R9386 dvdd.n133 dvdd.n97 0.120292
R9387 dvdd.n132 dvdd.n131 0.120292
R9388 dvdd.n131 dvdd.n99 0.120292
R9389 dvdd.n127 dvdd.n99 0.120292
R9390 dvdd.n127 dvdd.n126 0.120292
R9391 dvdd.n126 dvdd.n102 0.120292
R9392 dvdd.n122 dvdd.n102 0.120292
R9393 dvdd.n122 dvdd.n121 0.120292
R9394 dvdd.n121 dvdd.n120 0.120292
R9395 dvdd.n120 dvdd.n104 0.120292
R9396 dvdd.n116 dvdd.n104 0.120292
R9397 dvdd.n116 dvdd.n115 0.120292
R9398 dvdd.n111 dvdd.n110 0.120292
R9399 dvdd.n110 dvdd.n108 0.120292
R9400 dvdd.n290 dvdd.n289 0.120292
R9401 dvdd.n291 dvdd.n290 0.120292
R9402 dvdd.n297 dvdd 0.120292
R9403 dvdd.n298 dvdd.n297 0.120292
R9404 dvdd.n303 dvdd.n302 0.120292
R9405 dvdd.n304 dvdd.n303 0.120292
R9406 dvdd.n304 dvdd.n81 0.120292
R9407 dvdd.n309 dvdd.n81 0.120292
R9408 dvdd.n310 dvdd.n309 0.120292
R9409 dvdd.n311 dvdd.n310 0.120292
R9410 dvdd.n311 dvdd.n79 0.120292
R9411 dvdd.n315 dvdd.n79 0.120292
R9412 dvdd.n316 dvdd.n315 0.120292
R9413 dvdd.n317 dvdd.n316 0.120292
R9414 dvdd.n207 dvdd.n196 0.120292
R9415 dvdd.n214 dvdd.n196 0.120292
R9416 dvdd.n215 dvdd.n214 0.120292
R9417 dvdd.n277 dvdd.n216 0.120292
R9418 dvdd.n272 dvdd.n216 0.120292
R9419 dvdd.n272 dvdd.n271 0.120292
R9420 dvdd.n271 dvdd.n270 0.120292
R9421 dvdd.n270 dvdd.n218 0.120292
R9422 dvdd.n266 dvdd.n218 0.120292
R9423 dvdd.n266 dvdd.n265 0.120292
R9424 dvdd.n265 dvdd.n264 0.120292
R9425 dvdd.n264 dvdd.n221 0.120292
R9426 dvdd.n260 dvdd.n221 0.120292
R9427 dvdd.n260 dvdd.n259 0.120292
R9428 dvdd.n256 dvdd.n255 0.120292
R9429 dvdd.n255 dvdd.n224 0.120292
R9430 dvdd.n251 dvdd.n224 0.120292
R9431 dvdd.n251 dvdd.n250 0.120292
R9432 dvdd.n250 dvdd.n226 0.120292
R9433 dvdd.n246 dvdd.n226 0.120292
R9434 dvdd.n246 dvdd.n245 0.120292
R9435 dvdd.n245 dvdd.n244 0.120292
R9436 dvdd.n244 dvdd.n228 0.120292
R9437 dvdd.n240 dvdd.n228 0.120292
R9438 dvdd.n240 dvdd.n239 0.120292
R9439 dvdd.n236 dvdd.n235 0.120292
R9440 dvdd.n235 dvdd.n231 0.120292
R9441 dvdd.n389 dvdd.n388 0.120292
R9442 dvdd.n389 dvdd.n375 0.120292
R9443 dvdd.n393 dvdd.n375 0.120292
R9444 dvdd.n394 dvdd.n393 0.120292
R9445 dvdd.n394 dvdd.n373 0.120292
R9446 dvdd.n398 dvdd.n373 0.120292
R9447 dvdd.n399 dvdd.n398 0.120292
R9448 dvdd.n400 dvdd.n399 0.120292
R9449 dvdd.n400 dvdd.n371 0.120292
R9450 dvdd.n404 dvdd.n371 0.120292
R9451 dvdd.n405 dvdd.n404 0.120292
R9452 dvdd.n419 dvdd.n368 0.120292
R9453 dvdd.n420 dvdd.n419 0.120292
R9454 dvdd.n421 dvdd.n420 0.120292
R9455 dvdd.n421 dvdd.n366 0.120292
R9456 dvdd.n426 dvdd.n366 0.120292
R9457 dvdd.n427 dvdd.n426 0.120292
R9458 dvdd.n428 dvdd.n427 0.120292
R9459 dvdd.n428 dvdd.n364 0.120292
R9460 dvdd.n434 dvdd.n364 0.120292
R9461 dvdd.n436 dvdd.n361 0.120292
R9462 dvdd.n442 dvdd.n361 0.120292
R9463 dvdd.n443 dvdd.n442 0.120292
R9464 dvdd.n443 dvdd.n358 0.120292
R9465 dvdd.n449 dvdd.n358 0.120292
R9466 dvdd.n450 dvdd.n449 0.120292
R9467 dvdd.n451 dvdd.n450 0.120292
R9468 dvdd.n451 dvdd.n355 0.120292
R9469 dvdd.n457 dvdd.n355 0.120292
R9470 dvdd.n459 dvdd.n458 0.120292
R9471 dvdd.n459 dvdd.n353 0.120292
R9472 dvdd.n464 dvdd.n353 0.120292
R9473 dvdd.n521 dvdd.n520 0.120292
R9474 dvdd.n517 dvdd.n516 0.120292
R9475 dvdd.n516 dvdd.n467 0.120292
R9476 dvdd.n468 dvdd.n467 0.120292
R9477 dvdd.n509 dvdd.n468 0.120292
R9478 dvdd.n503 dvdd.n502 0.120292
R9479 dvdd.n502 dvdd.n473 0.120292
R9480 dvdd.n496 dvdd.n495 0.120292
R9481 dvdd.n495 dvdd.n494 0.120292
R9482 dvdd.n494 dvdd.n476 0.120292
R9483 dvdd.n490 dvdd.n476 0.120292
R9484 dvdd.n490 dvdd.n489 0.120292
R9485 dvdd.n489 dvdd.n481 0.120292
R9486 dvdd.n600 dvdd.n347 0.120292
R9487 dvdd.n600 dvdd.n599 0.120292
R9488 dvdd.n599 dvdd.n598 0.120292
R9489 dvdd.n591 dvdd.n590 0.120292
R9490 dvdd.n590 dvdd.n528 0.120292
R9491 dvdd.n585 dvdd.n528 0.120292
R9492 dvdd.n585 dvdd.n584 0.120292
R9493 dvdd.n584 dvdd.n583 0.120292
R9494 dvdd.n580 dvdd.n579 0.120292
R9495 dvdd.n579 dvdd.n578 0.120292
R9496 dvdd.n578 dvdd.n533 0.120292
R9497 dvdd.n573 dvdd.n572 0.120292
R9498 dvdd.n572 dvdd.n541 0.120292
R9499 dvdd.n568 dvdd.n541 0.120292
R9500 dvdd.n568 dvdd.n567 0.120292
R9501 dvdd.n567 dvdd.n543 0.120292
R9502 dvdd.n563 dvdd.n543 0.120292
R9503 dvdd.n563 dvdd.n562 0.120292
R9504 dvdd.n562 dvdd.n561 0.120292
R9505 dvdd.n561 dvdd.n545 0.120292
R9506 dvdd.n557 dvdd.n545 0.120292
R9507 dvdd.n557 dvdd.n556 0.120292
R9508 dvdd.n666 dvdd.n653 0.120292
R9509 dvdd.n672 dvdd.n653 0.120292
R9510 dvdd.n673 dvdd.n672 0.120292
R9511 dvdd.n680 dvdd.n679 0.120292
R9512 dvdd.n684 dvdd.n683 0.120292
R9513 dvdd.n684 dvdd.n648 0.120292
R9514 dvdd.n690 dvdd.n648 0.120292
R9515 dvdd.n691 dvdd.n690 0.120292
R9516 dvdd.n697 dvdd.n696 0.120292
R9517 dvdd.n697 dvdd.n644 0.120292
R9518 dvdd.n702 dvdd.n644 0.120292
R9519 dvdd.n711 dvdd.n642 0.120292
R9520 dvdd.n712 dvdd.n711 0.120292
R9521 dvdd.n713 dvdd.n712 0.120292
R9522 dvdd.n713 dvdd.n640 0.120292
R9523 dvdd.n718 dvdd.n640 0.120292
R9524 dvdd.n719 dvdd.n718 0.120292
R9525 dvdd.n719 dvdd.n637 0.120292
R9526 dvdd.n723 dvdd.n637 0.120292
R9527 dvdd.n724 dvdd.n723 0.120292
R9528 dvdd.n635 dvdd.n633 0.120292
R9529 dvdd.n733 dvdd.n633 0.120292
R9530 dvdd.n734 dvdd.n733 0.120292
R9531 dvdd.n735 dvdd.n734 0.120292
R9532 dvdd.n735 dvdd.n630 0.120292
R9533 dvdd.n741 dvdd.n630 0.120292
R9534 dvdd.n742 dvdd.n741 0.120292
R9535 dvdd.n742 dvdd.n628 0.120292
R9536 dvdd.n751 dvdd.n628 0.120292
R9537 dvdd.n752 dvdd.n751 0.120292
R9538 dvdd.n806 dvdd.n805 0.120292
R9539 dvdd.n805 dvdd.n756 0.120292
R9540 dvdd.n799 dvdd.n756 0.120292
R9541 dvdd.n799 dvdd.n798 0.120292
R9542 dvdd.n798 dvdd.n797 0.120292
R9543 dvdd.n797 dvdd.n759 0.120292
R9544 dvdd.n789 dvdd.n762 0.120292
R9545 dvdd.n783 dvdd.n762 0.120292
R9546 dvdd.n782 dvdd.n781 0.120292
R9547 dvdd.n781 dvdd.n766 0.120292
R9548 dvdd.n775 dvdd.n766 0.120292
R9549 dvdd.n894 dvdd.n623 0.120292
R9550 dvdd.n888 dvdd.n623 0.120292
R9551 dvdd.n888 dvdd.n887 0.120292
R9552 dvdd.n881 dvdd.n816 0.120292
R9553 dvdd.n876 dvdd.n816 0.120292
R9554 dvdd.n876 dvdd.n875 0.120292
R9555 dvdd.n875 dvdd.n874 0.120292
R9556 dvdd.n874 dvdd.n820 0.120292
R9557 dvdd.n869 dvdd.n820 0.120292
R9558 dvdd.n869 dvdd.n868 0.120292
R9559 dvdd.n868 dvdd.n867 0.120292
R9560 dvdd.n862 dvdd.n861 0.120292
R9561 dvdd.n861 dvdd.n830 0.120292
R9562 dvdd.n857 dvdd.n830 0.120292
R9563 dvdd.n857 dvdd.n856 0.120292
R9564 dvdd.n856 dvdd.n832 0.120292
R9565 dvdd.n852 dvdd.n832 0.120292
R9566 dvdd.n852 dvdd.n851 0.120292
R9567 dvdd.n851 dvdd.n850 0.120292
R9568 dvdd.n850 dvdd.n834 0.120292
R9569 dvdd.n846 dvdd.n834 0.120292
R9570 dvdd.n846 dvdd.n845 0.120292
R9571 dvdd.n971 dvdd.n953 0.120292
R9572 dvdd.n972 dvdd.n971 0.120292
R9573 dvdd.n980 dvdd.n951 0.120292
R9574 dvdd.n982 dvdd.n949 0.120292
R9575 dvdd.n988 dvdd.n946 0.120292
R9576 dvdd.n996 dvdd.n995 0.120292
R9577 dvdd.n997 dvdd.n996 0.120292
R9578 dvdd.n997 dvdd.n941 0.120292
R9579 dvdd.n1004 dvdd.n941 0.120292
R9580 dvdd.n1005 dvdd.n1004 0.120292
R9581 dvdd.n1006 dvdd.n1005 0.120292
R9582 dvdd.n1006 dvdd.n939 0.120292
R9583 dvdd.n1011 dvdd.n939 0.120292
R9584 dvdd.n1012 dvdd.n1011 0.120292
R9585 dvdd.n1012 dvdd.n936 0.120292
R9586 dvdd.n1018 dvdd.n936 0.120292
R9587 dvdd.n1019 dvdd.n1018 0.120292
R9588 dvdd.n1020 dvdd.n1019 0.120292
R9589 dvdd.n1020 dvdd.n934 0.120292
R9590 dvdd.n1024 dvdd.n934 0.120292
R9591 dvdd.n1025 dvdd.n1024 0.120292
R9592 dvdd.n1026 dvdd.n1025 0.120292
R9593 dvdd.n1036 dvdd.n1035 0.120292
R9594 dvdd.n1049 dvdd.n929 0.120292
R9595 dvdd.n1050 dvdd.n1049 0.120292
R9596 dvdd.n1096 dvdd.n1053 0.120292
R9597 dvdd.n1091 dvdd.n1053 0.120292
R9598 dvdd.n1086 dvdd.n1085 0.120292
R9599 dvdd.n1085 dvdd.n1084 0.120292
R9600 dvdd.n1078 dvdd.n1060 0.120292
R9601 dvdd.n1078 dvdd.n1077 0.120292
R9602 dvdd.n1077 dvdd.n1076 0.120292
R9603 dvdd.n1072 dvdd.n1071 0.120292
R9604 dvdd.n1186 dvdd.n1185 0.120292
R9605 dvdd.n1182 dvdd.n1181 0.120292
R9606 dvdd.n1181 dvdd.n926 0.120292
R9607 dvdd.n1170 dvdd.n1103 0.120292
R9608 dvdd.n1170 dvdd.n1169 0.120292
R9609 dvdd.n1163 dvdd.n1109 0.120292
R9610 dvdd.n1163 dvdd.n1162 0.120292
R9611 dvdd.n1162 dvdd.n1161 0.120292
R9612 dvdd.n1158 dvdd.n1157 0.120292
R9613 dvdd.n1157 dvdd.n1113 0.120292
R9614 dvdd.n1152 dvdd.n1113 0.120292
R9615 dvdd.n1152 dvdd.n1151 0.120292
R9616 dvdd.n1151 dvdd.n1116 0.120292
R9617 dvdd.n1146 dvdd.n1116 0.120292
R9618 dvdd.n1146 dvdd.n1145 0.120292
R9619 dvdd.n1141 dvdd.n1140 0.120292
R9620 dvdd.n1136 dvdd.n1121 0.120292
R9621 dvdd.n1131 dvdd.n1121 0.120292
R9622 dvdd.n1266 dvdd.n1265 0.120292
R9623 dvdd.n1271 dvdd.n1270 0.120292
R9624 dvdd.n1271 dvdd.n1253 0.120292
R9625 dvdd.n1277 dvdd.n1250 0.120292
R9626 dvdd.n1278 dvdd.n1277 0.120292
R9627 dvdd.n1279 dvdd.n1278 0.120292
R9628 dvdd.n1279 dvdd.n1246 0.120292
R9629 dvdd.n1284 dvdd.n1246 0.120292
R9630 dvdd.n1242 dvdd.n1241 0.120292
R9631 dvdd.n1294 dvdd.n1293 0.120292
R9632 dvdd.n1294 dvdd.n1235 0.120292
R9633 dvdd.n1299 dvdd.n1235 0.120292
R9634 dvdd.n1300 dvdd.n1299 0.120292
R9635 dvdd.n1300 dvdd.n1232 0.120292
R9636 dvdd.n1305 dvdd.n1232 0.120292
R9637 dvdd.n1306 dvdd.n1305 0.120292
R9638 dvdd.n1307 dvdd.n1306 0.120292
R9639 dvdd.n1307 dvdd.n1230 0.120292
R9640 dvdd.n1312 dvdd.n1230 0.120292
R9641 dvdd.n1313 dvdd.n1312 0.120292
R9642 dvdd.n1317 dvdd.n1227 0.120292
R9643 dvdd.n1318 dvdd.n1317 0.120292
R9644 dvdd.n1323 dvdd.n1222 0.120292
R9645 dvdd.n1377 dvdd.n1376 0.120292
R9646 dvdd.n1376 dvdd.n1375 0.120292
R9647 dvdd.n1375 dvdd.n1328 0.120292
R9648 dvdd.n1336 dvdd.n1333 0.120292
R9649 dvdd.n1337 dvdd.n1336 0.120292
R9650 dvdd.n1365 dvdd.n1337 0.120292
R9651 dvdd.n1365 dvdd.n1364 0.120292
R9652 dvdd.n1359 dvdd.n1343 0.120292
R9653 dvdd.n1353 dvdd.n1343 0.120292
R9654 dvdd.n1353 dvdd.n1352 0.120292
R9655 dvdd.n1352 dvdd.n1348 0.120292
R9656 dvdd.n1470 dvdd.n1469 0.120292
R9657 dvdd.n1469 dvdd.n1211 0.120292
R9658 dvdd.n1463 dvdd.n1211 0.120292
R9659 dvdd.n1463 dvdd.n1462 0.120292
R9660 dvdd.n1457 dvdd.n1456 0.120292
R9661 dvdd.n1456 dvdd.n1389 0.120292
R9662 dvdd.n1450 dvdd.n1389 0.120292
R9663 dvdd.n1450 dvdd.n1449 0.120292
R9664 dvdd.n1449 dvdd.n1448 0.120292
R9665 dvdd.n1448 dvdd.n1395 0.120292
R9666 dvdd.n1396 dvdd.n1395 0.120292
R9667 dvdd.n1397 dvdd.n1396 0.120292
R9668 dvdd.n1442 dvdd.n1397 0.120292
R9669 dvdd.n1442 dvdd.n1441 0.120292
R9670 dvdd.n1441 dvdd.n1440 0.120292
R9671 dvdd.n1437 dvdd.n1436 0.120292
R9672 dvdd.n1435 dvdd.n1404 0.120292
R9673 dvdd.n1431 dvdd.n1404 0.120292
R9674 dvdd.n1431 dvdd.n1430 0.120292
R9675 dvdd.n1430 dvdd.n1429 0.120292
R9676 dvdd.n1429 dvdd.n1407 0.120292
R9677 dvdd.n1423 dvdd.n1422 0.120292
R9678 dvdd.n1558 dvdd.n1541 0.120292
R9679 dvdd.n1559 dvdd.n1558 0.120292
R9680 dvdd.n1565 dvdd.n1564 0.120292
R9681 dvdd.n1571 dvdd.n1535 0.120292
R9682 dvdd.n1572 dvdd.n1571 0.120292
R9683 dvdd.n1572 dvdd.n1532 0.120292
R9684 dvdd.n1578 dvdd.n1532 0.120292
R9685 dvdd.n1582 dvdd.n1524 0.120292
R9686 dvdd.n1589 dvdd.n1524 0.120292
R9687 dvdd.n1590 dvdd.n1589 0.120292
R9688 dvdd.n1521 dvdd.n1515 0.120292
R9689 dvdd.n1597 dvdd.n1515 0.120292
R9690 dvdd.n1598 dvdd.n1597 0.120292
R9691 dvdd.n1604 dvdd.n1603 0.120292
R9692 dvdd.n1605 dvdd.n1604 0.120292
R9693 dvdd.n1612 dvdd.n1511 0.120292
R9694 dvdd.n1613 dvdd.n1612 0.120292
R9695 dvdd.n1614 dvdd.n1508 0.120292
R9696 dvdd.n1618 dvdd.n1508 0.120292
R9697 dvdd.n1619 dvdd.n1618 0.120292
R9698 dvdd.n1619 dvdd.n1505 0.120292
R9699 dvdd.n1505 dvdd.n1503 0.120292
R9700 dvdd.n1624 dvdd.n1503 0.120292
R9701 dvdd.n1625 dvdd.n1624 0.120292
R9702 dvdd.n1677 dvdd.n1676 0.120292
R9703 dvdd.n1676 dvdd.n1627 0.120292
R9704 dvdd.n1672 dvdd.n1627 0.120292
R9705 dvdd.n1671 dvdd.n1670 0.120292
R9706 dvdd.n1670 dvdd.n1631 0.120292
R9707 dvdd.n1666 dvdd.n1631 0.120292
R9708 dvdd.n1666 dvdd.n1665 0.120292
R9709 dvdd.n1665 dvdd.n1634 0.120292
R9710 dvdd.n1655 dvdd.n1639 0.120292
R9711 dvdd.n1655 dvdd.n1654 0.120292
R9712 dvdd.n1651 dvdd.n1650 0.120292
R9713 dvdd.n1650 dvdd.n1649 0.120292
R9714 dvdd.n1649 dvdd.n1641 0.120292
R9715 dvdd.n1643 dvdd.n1641 0.120292
R9716 dvdd.n1769 dvdd.n1768 0.120292
R9717 dvdd.n1768 dvdd.n1497 0.120292
R9718 dvdd.n1763 dvdd.n1497 0.120292
R9719 dvdd.n1763 dvdd.n1762 0.120292
R9720 dvdd.n1757 dvdd.n1756 0.120292
R9721 dvdd.n1750 dvdd.n1689 0.120292
R9722 dvdd.n1745 dvdd.n1689 0.120292
R9723 dvdd.n1745 dvdd.n1744 0.120292
R9724 dvdd.n1744 dvdd.n1692 0.120292
R9725 dvdd.n1739 dvdd.n1692 0.120292
R9726 dvdd.n1739 dvdd.n1738 0.120292
R9727 dvdd.n1738 dvdd.n1737 0.120292
R9728 dvdd.n1737 dvdd.n1695 0.120292
R9729 dvdd.n1731 dvdd.n1695 0.120292
R9730 dvdd.n1731 dvdd.n1730 0.120292
R9731 dvdd.n1730 dvdd.n1699 0.120292
R9732 dvdd.n1726 dvdd.n1699 0.120292
R9733 dvdd.n1726 dvdd.n1725 0.120292
R9734 dvdd.n1725 dvdd.n1724 0.120292
R9735 dvdd.n1724 dvdd.n1702 0.120292
R9736 dvdd.n1718 dvdd.n1702 0.120292
R9737 dvdd.n1718 dvdd.n1717 0.120292
R9738 dvdd.n1717 dvdd.n1716 0.120292
R9739 dvdd.n1847 dvdd.n1846 0.120292
R9740 dvdd.n1847 dvdd.n1830 0.120292
R9741 dvdd.n1853 dvdd.n1830 0.120292
R9742 dvdd.n1854 dvdd.n1853 0.120292
R9743 dvdd.n1860 dvdd.n1859 0.120292
R9744 dvdd.n1861 dvdd.n1860 0.120292
R9745 dvdd.n1861 dvdd.n1827 0.120292
R9746 dvdd.n1866 dvdd.n1827 0.120292
R9747 dvdd.n1871 dvdd.n1870 0.120292
R9748 dvdd.n1872 dvdd.n1871 0.120292
R9749 dvdd.n1878 dvdd.n1877 0.120292
R9750 dvdd.n1878 dvdd.n1821 0.120292
R9751 dvdd.n1884 dvdd.n1821 0.120292
R9752 dvdd.n1885 dvdd.n1884 0.120292
R9753 dvdd.n1886 dvdd.n1885 0.120292
R9754 dvdd.n1886 dvdd.n1818 0.120292
R9755 dvdd.n1892 dvdd.n1818 0.120292
R9756 dvdd.n1893 dvdd.n1892 0.120292
R9757 dvdd.n1894 dvdd.n1893 0.120292
R9758 dvdd.n1894 dvdd.n1816 0.120292
R9759 dvdd.n1900 dvdd.n1816 0.120292
R9760 dvdd.n1901 dvdd.n1900 0.120292
R9761 dvdd.n1902 dvdd.n1901 0.120292
R9762 dvdd.n1902 dvdd.n1814 0.120292
R9763 dvdd.n1908 dvdd.n1814 0.120292
R9764 dvdd.n1909 dvdd.n1908 0.120292
R9765 dvdd.n1914 dvdd.n1812 0.120292
R9766 dvdd.n1916 dvdd.n1809 0.120292
R9767 dvdd.n1924 dvdd.n1809 0.120292
R9768 dvdd.n1925 dvdd.n1924 0.120292
R9769 dvdd.n1987 dvdd.n1986 0.120292
R9770 dvdd.n1983 dvdd.n1982 0.120292
R9771 dvdd.n1978 dvdd.n1932 0.120292
R9772 dvdd.n1972 dvdd.n1932 0.120292
R9773 dvdd.n1972 dvdd.n1971 0.120292
R9774 dvdd.n1971 dvdd.n1970 0.120292
R9775 dvdd.n1970 dvdd.n1938 0.120292
R9776 dvdd.n1964 dvdd.n1938 0.120292
R9777 dvdd.n1964 dvdd.n1963 0.120292
R9778 dvdd.n1963 dvdd.n1942 0.120292
R9779 dvdd.n1957 dvdd.n1942 0.120292
R9780 dvdd.n1957 dvdd.n1956 0.120292
R9781 dvdd.n1956 dvdd.n1955 0.120292
R9782 dvdd.n1955 dvdd.n1947 0.120292
R9783 dvdd.n1949 dvdd.n1947 0.120292
R9784 dvdd.n2073 dvdd.n2072 0.120292
R9785 dvdd.n2072 dvdd.n1807 0.120292
R9786 dvdd.n2064 dvdd.n1999 0.120292
R9787 dvdd.n2058 dvdd.n1999 0.120292
R9788 dvdd.n2058 dvdd.n2057 0.120292
R9789 dvdd.n2057 dvdd.n2056 0.120292
R9790 dvdd.n2056 dvdd.n2001 0.120292
R9791 dvdd.n2052 dvdd.n2001 0.120292
R9792 dvdd.n2052 dvdd.n2051 0.120292
R9793 dvdd.n2051 dvdd.n2050 0.120292
R9794 dvdd.n2050 dvdd.n2006 0.120292
R9795 dvdd.n2045 dvdd.n2006 0.120292
R9796 dvdd.n2045 dvdd.n2044 0.120292
R9797 dvdd.n2034 dvdd.n2033 0.120292
R9798 dvdd.n2033 dvdd.n2015 0.120292
R9799 dvdd.n2029 dvdd.n2015 0.120292
R9800 dvdd.n2028 dvdd.n2027 0.120292
R9801 dvdd.n2248 dvdd.n2247 0.120292
R9802 dvdd.n2248 dvdd.n2234 0.120292
R9803 dvdd.n2252 dvdd.n2234 0.120292
R9804 dvdd.n2253 dvdd.n2252 0.120292
R9805 dvdd.n2253 dvdd.n2232 0.120292
R9806 dvdd.n2257 dvdd.n2232 0.120292
R9807 dvdd.n2258 dvdd.n2257 0.120292
R9808 dvdd.n2259 dvdd.n2258 0.120292
R9809 dvdd.n2259 dvdd.n2230 0.120292
R9810 dvdd.n2264 dvdd.n2230 0.120292
R9811 dvdd.n2265 dvdd.n2264 0.120292
R9812 dvdd.n2271 dvdd.n2270 0.120292
R9813 dvdd.n2272 dvdd.n2271 0.120292
R9814 dvdd.n2277 dvdd.n2276 0.120292
R9815 dvdd.n2277 dvdd.n2138 0.120292
R9816 dvdd.n2281 dvdd.n2138 0.120292
R9817 dvdd.n2282 dvdd.n2281 0.120292
R9818 dvdd.n2282 dvdd.n2136 0.120292
R9819 dvdd.n2287 dvdd.n2136 0.120292
R9820 dvdd.n2288 dvdd.n2287 0.120292
R9821 dvdd.n2289 dvdd.n2134 0.120292
R9822 dvdd.n2294 dvdd.n2134 0.120292
R9823 dvdd.n2295 dvdd.n2294 0.120292
R9824 dvdd.n2300 dvdd.n2299 0.120292
R9825 dvdd.n2300 dvdd.n2131 0.120292
R9826 dvdd.n2304 dvdd.n2131 0.120292
R9827 dvdd.n2305 dvdd.n2304 0.120292
R9828 dvdd.n2305 dvdd.n2129 0.120292
R9829 dvdd.n2309 dvdd.n2129 0.120292
R9830 dvdd.n2310 dvdd.n2309 0.120292
R9831 dvdd.n2314 dvdd.n2313 0.120292
R9832 dvdd.n2314 dvdd.n2125 0.120292
R9833 dvdd dvdd.n2125 0.120292
R9834 dvdd.n2320 dvdd.n2122 0.120292
R9835 dvdd.n2328 dvdd.n2122 0.120292
R9836 dvdd.n2120 dvdd.n2118 0.120292
R9837 dvdd.n2338 dvdd.n2117 0.120292
R9838 dvdd.n2339 dvdd.n2338 0.120292
R9839 dvdd.n2343 dvdd.n2114 0.120292
R9840 dvdd.n2344 dvdd.n2111 0.120292
R9841 dvdd.n2348 dvdd.n2111 0.120292
R9842 dvdd.n2349 dvdd.n2348 0.120292
R9843 dvdd.n2155 dvdd.n2095 0.120292
R9844 dvdd.n2155 dvdd.n2151 0.120292
R9845 dvdd.n2160 dvdd.n2151 0.120292
R9846 dvdd.n2222 dvdd.n2174 0.120292
R9847 dvdd.n2216 dvdd.n2174 0.120292
R9848 dvdd.n2216 dvdd.n2215 0.120292
R9849 dvdd.n2215 dvdd.n2214 0.120292
R9850 dvdd.n2214 dvdd.n2177 0.120292
R9851 dvdd.n2210 dvdd.n2177 0.120292
R9852 dvdd.n2210 dvdd.n2209 0.120292
R9853 dvdd.n2209 dvdd.n2208 0.120292
R9854 dvdd.n2204 dvdd.n2203 0.120292
R9855 dvdd.n2199 dvdd.n2198 0.120292
R9856 dvdd.n2198 dvdd.n2187 0.120292
R9857 dvdd.n2424 dvdd.n2410 0.120292
R9858 dvdd.n2431 dvdd.n2410 0.120292
R9859 dvdd.n2432 dvdd.n2431 0.120292
R9860 dvdd.n2433 dvdd.n2432 0.120292
R9861 dvdd.n2433 dvdd.n2408 0.120292
R9862 dvdd.n2437 dvdd.n2408 0.120292
R9863 dvdd.n2438 dvdd.n2437 0.120292
R9864 dvdd.n2443 dvdd.n2406 0.120292
R9865 dvdd.n2444 dvdd.n2443 0.120292
R9866 dvdd.n2452 dvdd.n2451 0.120292
R9867 dvdd.n2452 dvdd.n2402 0.120292
R9868 dvdd.n2457 dvdd.n2402 0.120292
R9869 dvdd.n2470 dvdd.n2469 0.120292
R9870 dvdd.n2471 dvdd.n2470 0.120292
R9871 dvdd.n2480 dvdd.n2479 0.120292
R9872 dvdd.n2480 dvdd.n2396 0.120292
R9873 dvdd.n2486 dvdd.n2396 0.120292
R9874 dvdd.n2496 dvdd.n2390 0.120292
R9875 dvdd.n2497 dvdd.n2496 0.120292
R9876 dvdd.n2498 dvdd.n2497 0.120292
R9877 dvdd.n2502 dvdd.n2501 0.120292
R9878 dvdd.n2552 dvdd.n2551 0.120292
R9879 dvdd.n2551 dvdd.n2503 0.120292
R9880 dvdd.n2544 dvdd.n2515 0.120292
R9881 dvdd.n2544 dvdd.n2543 0.120292
R9882 dvdd.n2543 dvdd.n2518 0.120292
R9883 dvdd.n2538 dvdd.n2518 0.120292
R9884 dvdd.n2538 dvdd.n2537 0.120292
R9885 dvdd.n2533 dvdd.n2532 0.120292
R9886 dvdd.n2532 dvdd.n2523 0.120292
R9887 dvdd.n2636 dvdd.n2378 0.120292
R9888 dvdd.n2630 dvdd.n2629 0.120292
R9889 dvdd.n2629 dvdd.n2559 0.120292
R9890 dvdd.n2624 dvdd.n2559 0.120292
R9891 dvdd.n2624 dvdd.n2623 0.120292
R9892 dvdd.n2618 dvdd.n2617 0.120292
R9893 dvdd.n2617 dvdd.n2566 0.120292
R9894 dvdd.n2610 dvdd.n2609 0.120292
R9895 dvdd.n2609 dvdd.n2568 0.120292
R9896 dvdd.n2605 dvdd.n2568 0.120292
R9897 dvdd.n2605 dvdd.n2604 0.120292
R9898 dvdd.n2604 dvdd.n2574 0.120292
R9899 dvdd.n2598 dvdd.n2597 0.120292
R9900 dvdd.n2593 dvdd.n2592 0.120292
R9901 dvdd.n2592 dvdd.n2579 0.120292
R9902 dvdd.n2894 dvdd.n2893 0.120292
R9903 dvdd.n2895 dvdd.n2894 0.120292
R9904 dvdd.n2895 dvdd.n2884 0.120292
R9905 dvdd.n2902 dvdd.n2884 0.120292
R9906 dvdd.n2903 dvdd.n2902 0.120292
R9907 dvdd.n2904 dvdd.n2903 0.120292
R9908 dvdd.n2904 dvdd.n2881 0.120292
R9909 dvdd.n2911 dvdd.n2881 0.120292
R9910 dvdd.n2912 dvdd.n2911 0.120292
R9911 dvdd.n2912 dvdd.n2877 0.120292
R9912 dvdd.n2917 dvdd.n2877 0.120292
R9913 dvdd.n2918 dvdd.n2917 0.120292
R9914 dvdd.n2923 dvdd.n2922 0.120292
R9915 dvdd.n2924 dvdd.n2923 0.120292
R9916 dvdd.n2924 dvdd.n2873 0.120292
R9917 dvdd.n2928 dvdd.n2873 0.120292
R9918 dvdd.n3048 dvdd.n3047 0.120292
R9919 dvdd.n3049 dvdd.n3048 0.120292
R9920 dvdd.n3049 dvdd.n3038 0.120292
R9921 dvdd.n3056 dvdd.n3038 0.120292
R9922 dvdd.n3057 dvdd.n3056 0.120292
R9923 dvdd.n3058 dvdd.n3057 0.120292
R9924 dvdd.n3058 dvdd.n3035 0.120292
R9925 dvdd.n3065 dvdd.n3035 0.120292
R9926 dvdd.n3066 dvdd.n3065 0.120292
R9927 dvdd.n3066 dvdd.n3031 0.120292
R9928 dvdd.n3071 dvdd.n3031 0.120292
R9929 dvdd.n3072 dvdd.n3071 0.120292
R9930 dvdd.n3077 dvdd.n3076 0.120292
R9931 dvdd.n3078 dvdd.n3077 0.120292
R9932 dvdd.n3078 dvdd.n3027 0.120292
R9933 dvdd.n3082 dvdd.n3027 0.120292
R9934 dvdd.n2991 dvdd.n2990 0.120292
R9935 dvdd.n2992 dvdd.n2991 0.120292
R9936 dvdd.n2992 dvdd.n2981 0.120292
R9937 dvdd.n2999 dvdd.n2981 0.120292
R9938 dvdd.n3000 dvdd.n2999 0.120292
R9939 dvdd.n3001 dvdd.n3000 0.120292
R9940 dvdd.n3001 dvdd.n2978 0.120292
R9941 dvdd.n3008 dvdd.n2978 0.120292
R9942 dvdd.n3009 dvdd.n3008 0.120292
R9943 dvdd.n3009 dvdd.n2974 0.120292
R9944 dvdd.n3014 dvdd.n2974 0.120292
R9945 dvdd.n3015 dvdd.n3014 0.120292
R9946 dvdd.n3020 dvdd.n3019 0.120292
R9947 dvdd.n3021 dvdd.n3020 0.120292
R9948 dvdd.n3021 dvdd.n2970 0.120292
R9949 dvdd.n3025 dvdd.n2970 0.120292
R9950 dvdd.n2828 dvdd.n2827 0.120292
R9951 dvdd.n2829 dvdd.n2828 0.120292
R9952 dvdd.n2829 dvdd.n2818 0.120292
R9953 dvdd.n2836 dvdd.n2818 0.120292
R9954 dvdd.n2837 dvdd.n2836 0.120292
R9955 dvdd.n2838 dvdd.n2837 0.120292
R9956 dvdd.n2838 dvdd.n2815 0.120292
R9957 dvdd.n2843 dvdd.n2815 0.120292
R9958 dvdd.n2844 dvdd.n2843 0.120292
R9959 dvdd.n2844 dvdd.n2811 0.120292
R9960 dvdd.n2851 dvdd.n2811 0.120292
R9961 dvdd.n2852 dvdd.n2851 0.120292
R9962 dvdd.n2856 dvdd.n2855 0.120292
R9963 dvdd.n2856 dvdd.n2807 0.120292
R9964 dvdd.n2860 dvdd.n2807 0.120292
R9965 dvdd.n2861 dvdd.n2860 0.120292
R9966 dvdd.n2866 dvdd.n2865 0.120292
R9967 dvdd.n2867 dvdd.n2866 0.120292
R9968 dvdd.n2867 dvdd.n2803 0.120292
R9969 dvdd.n2871 dvdd.n2803 0.120292
R9970 dvdd.n411 dvdd.n410 0.106285
R9971 dvdd.n2043 dvdd.n2008 0.106285
R9972 dvdd.n384 dvdd 0.105238
R9973 dvdd.n659 dvdd 0.105238
R9974 dvdd.n961 dvdd 0.105238
R9975 dvdd.n1264 dvdd 0.105238
R9976 dvdd.n1547 dvdd 0.105238
R9977 dvdd.n1840 dvdd 0.105238
R9978 dvdd.n2243 dvdd 0.105238
R9979 dvdd.n2419 dvdd 0.105238
R9980 dvdd.n1609 dvdd.n1510 0.102087
R9981 dvdd.n1930 dvdd.n1929 0.102087
R9982 dvdd.n2157 dvdd.n2156 0.102087
R9983 dvdd.n2596 dvdd.n2577 0.102087
R9984 dvdd.n982 dvdd 0.0994583
R9985 dvdd dvdd.n946 0.0994583
R9986 dvdd.n168 dvdd 0.0981562
R9987 dvdd dvdd.n155 0.0981562
R9988 dvdd.n112 dvdd 0.0981562
R9989 dvdd dvdd.n111 0.0981562
R9990 dvdd.n289 dvdd 0.0981562
R9991 dvdd.n256 dvdd 0.0981562
R9992 dvdd.n236 dvdd 0.0981562
R9993 dvdd.n412 dvdd 0.0981562
R9994 dvdd.n436 dvdd 0.0981562
R9995 dvdd.n458 dvdd 0.0981562
R9996 dvdd.n679 dvdd 0.0981562
R9997 dvdd dvdd.n642 0.0981562
R9998 dvdd dvdd.n635 0.0981562
R9999 dvdd dvdd.n953 0.0981562
R10000 dvdd.n1044 dvdd 0.0981562
R10001 dvdd dvdd.n929 0.0981562
R10002 dvdd.n1109 dvdd 0.0981562
R10003 dvdd dvdd.n1141 0.0981562
R10004 dvdd dvdd.n1250 0.0981562
R10005 dvdd dvdd.n1227 0.0981562
R10006 dvdd dvdd.n1224 0.0981562
R10007 dvdd.n1325 dvdd 0.0981562
R10008 dvdd dvdd.n1377 0.0981562
R10009 dvdd.n1333 dvdd 0.0981562
R10010 dvdd dvdd.n1359 0.0981562
R10011 dvdd.n1411 dvdd 0.0981562
R10012 dvdd.n1564 dvdd 0.0981562
R10013 dvdd dvdd.n1521 0.0981562
R10014 dvdd dvdd.n1750 0.0981562
R10015 dvdd.n1867 dvdd 0.0981562
R10016 dvdd dvdd.n1978 0.0981562
R10017 dvdd.n2040 dvdd 0.0981562
R10018 dvdd dvdd.n2038 0.0981562
R10019 dvdd.n2266 dvdd 0.0981562
R10020 dvdd.n2289 dvdd 0.0981562
R10021 dvdd.n2299 dvdd 0.0981562
R10022 dvdd.n2313 dvdd 0.0981562
R10023 dvdd dvdd.n2120 0.0981562
R10024 dvdd.n2205 dvdd 0.0981562
R10025 dvdd dvdd.n2204 0.0981562
R10026 dvdd dvdd.n2199 0.0981562
R10027 dvdd.n2450 dvdd 0.0981562
R10028 dvdd.n2469 dvdd 0.0981562
R10029 dvdd.n2488 dvdd 0.0981562
R10030 dvdd dvdd.n2630 0.0981562
R10031 dvdd.n806 dvdd 0.0968542
R10032 dvdd.n1086 dvdd 0.0968542
R10033 dvdd.n1270 dvdd 0.0968542
R10034 dvdd.n1757 dvdd 0.0968542
R10035 dvdd dvdd.n2034 0.0968542
R10036 dvdd.n326 dvdd.n325 0.0950946
R10037 dvdd.n204 dvdd.n203 0.0950946
R10038 dvdd.n609 dvdd.n608 0.0950946
R10039 dvdd.n345 dvdd.n344 0.0950946
R10040 dvdd.n910 dvdd.n909 0.0950946
R10041 dvdd.n900 dvdd.n899 0.0950946
R10042 dvdd.n1199 dvdd.n1198 0.0950946
R10043 dvdd.n1191 dvdd.n1190 0.0950946
R10044 dvdd.n1483 dvdd.n1482 0.0950946
R10045 dvdd.n1475 dvdd.n1474 0.0950946
R10046 dvdd.n1784 dvdd.n1783 0.0950946
R10047 dvdd.n1774 dvdd.n1773 0.0950946
R10048 dvdd.n2086 dvdd.n2085 0.0950946
R10049 dvdd.n1804 dvdd.n1803 0.0950946
R10050 dvdd.n2356 dvdd.n2355 0.0950946
R10051 dvdd.n2101 dvdd.n2100 0.0950946
R10052 dvdd.n2644 dvdd.n2643 0.0950946
R10053 dvdd.n2376 dvdd.n2375 0.0950946
R10054 dvdd dvdd.n2646 0.08745
R10055 dvdd.n343 dvdd.n334 0.0838333
R10056 dvdd.n622 dvdd.n617 0.0838333
R10057 dvdd.n1496 dvdd.n1491 0.0838333
R10058 dvdd.n1802 dvdd.n1792 0.0838333
R10059 dvdd.n2096 dvdd.n2094 0.0838333
R10060 dvdd.n2374 dvdd.n2364 0.0838333
R10061 dvdd.n539 dvdd 0.082648
R10062 dvdd dvdd.n1064 0.082648
R10063 dvdd.n1239 dvdd 0.082648
R10064 dvdd dvdd.n2507 0.082648
R10065 dvdd.n2384 dvdd 0.082648
R10066 dvdd dvdd.n435 0.082648
R10067 dvdd.n703 dvdd 0.082648
R10068 dvdd dvdd.n2487 0.082648
R10069 dvdd.n2510 dvdd 0.0813459
R10070 dvdd.n324 dvdd.n323 0.0812292
R10071 dvdd.n607 dvdd.n606 0.0812292
R10072 dvdd.n908 dvdd.n907 0.0812292
R10073 dvdd.n1197 dvdd.n1196 0.0812292
R10074 dvdd.n1782 dvdd.n1781 0.0812292
R10075 dvdd.n2084 dvdd.n2083 0.0812292
R10076 dvdd.n2354 dvdd.n2353 0.0812292
R10077 dvdd.n2642 dvdd.n2641 0.0812292
R10078 dvdd.n3153 dvdd.n3151 0.0789314
R10079 dvdd.n317 dvdd.n74 0.0760208
R10080 dvdd.n485 dvdd.n331 0.0760208
R10081 dvdd.n773 dvdd.n614 0.0760208
R10082 dvdd.n1348 dvdd.n1204 0.0760208
R10083 dvdd.n1949 dvdd.n1789 0.0760208
R10084 dvdd.n2759 dvdd.n2647 0.074995
R10085 dvdd.n206 dvdd.n205 0.0708125
R10086 dvdd.n347 dvdd.n346 0.0708125
R10087 dvdd.n1476 dvdd.n1470 0.0708125
R10088 dvdd.n1775 dvdd.n1769 0.0708125
R10089 dvdd.n2102 dvdd.n2095 0.0708125
R10090 dvdd.n199 dvdd.n75 0.0680676
R10091 dvdd.n201 dvdd.n199 0.0680676
R10092 dvdd.n340 dvdd.n332 0.0680676
R10093 dvdd.n342 dvdd.n340 0.0680676
R10094 dvdd.n896 dvdd.n615 0.0680676
R10095 dvdd.n898 dvdd.n896 0.0680676
R10096 dvdd.n1187 dvdd.n916 0.0680676
R10097 dvdd.n1189 dvdd.n1187 0.0680676
R10098 dvdd.n1471 dvdd.n1205 0.0680676
R10099 dvdd.n1473 dvdd.n1471 0.0680676
R10100 dvdd.n1770 dvdd.n1489 0.0680676
R10101 dvdd.n1772 dvdd.n1770 0.0680676
R10102 dvdd.n1799 dvdd.n1790 0.0680676
R10103 dvdd.n1801 dvdd.n1799 0.0680676
R10104 dvdd.n2097 dvdd.n2092 0.0680676
R10105 dvdd.n2099 dvdd.n2097 0.0680676
R10106 dvdd.n2371 dvdd.n2362 0.0680676
R10107 dvdd.n2373 dvdd.n2371 0.0680676
R10108 dvdd.n202 dvdd 0.0656042
R10109 dvdd.n2761 dvdd.n2760 0.063
R10110 dvdd dvdd.n169 0.0603958
R10111 dvdd.n170 dvdd 0.0603958
R10112 dvdd.n173 dvdd 0.0603958
R10113 dvdd dvdd.n154 0.0603958
R10114 dvdd.n148 dvdd 0.0603958
R10115 dvdd dvdd.n132 0.0603958
R10116 dvdd.n108 dvdd 0.0603958
R10117 dvdd.n284 dvdd 0.0603958
R10118 dvdd.n285 dvdd 0.0603958
R10119 dvdd.n286 dvdd 0.0603958
R10120 dvdd.n291 dvdd 0.0603958
R10121 dvdd.n302 dvdd 0.0603958
R10122 dvdd dvdd.n206 0.0603958
R10123 dvdd.n207 dvdd 0.0603958
R10124 dvdd.n279 dvdd 0.0603958
R10125 dvdd dvdd.n278 0.0603958
R10126 dvdd dvdd.n277 0.0603958
R10127 dvdd.n385 dvdd 0.0603958
R10128 dvdd.n388 dvdd 0.0603958
R10129 dvdd.n413 dvdd 0.0603958
R10130 dvdd dvdd.n368 0.0603958
R10131 dvdd.n522 dvdd 0.0603958
R10132 dvdd dvdd.n521 0.0603958
R10133 dvdd.n517 dvdd 0.0603958
R10134 dvdd dvdd.n508 0.0603958
R10135 dvdd.n503 dvdd 0.0603958
R10136 dvdd.n496 dvdd 0.0603958
R10137 dvdd.n485 dvdd 0.0603958
R10138 dvdd.n595 dvdd 0.0603958
R10139 dvdd dvdd.n594 0.0603958
R10140 dvdd.n591 dvdd 0.0603958
R10141 dvdd.n580 dvdd 0.0603958
R10142 dvdd dvdd.n538 0.0603958
R10143 dvdd.n573 dvdd 0.0603958
R10144 dvdd.n665 dvdd 0.0603958
R10145 dvdd.n666 dvdd 0.0603958
R10146 dvdd.n674 dvdd 0.0603958
R10147 dvdd.n683 dvdd 0.0603958
R10148 dvdd dvdd.n691 0.0603958
R10149 dvdd.n692 dvdd 0.0603958
R10150 dvdd.n696 dvdd 0.0603958
R10151 dvdd.n811 dvdd 0.0603958
R10152 dvdd dvdd.n810 0.0603958
R10153 dvdd.n791 dvdd 0.0603958
R10154 dvdd.n791 dvdd 0.0603958
R10155 dvdd dvdd.n790 0.0603958
R10156 dvdd dvdd.n789 0.0603958
R10157 dvdd dvdd.n782 0.0603958
R10158 dvdd dvdd.n774 0.0603958
R10159 dvdd dvdd.n773 0.0603958
R10160 dvdd dvdd.n895 0.0603958
R10161 dvdd dvdd.n894 0.0603958
R10162 dvdd.n883 dvdd 0.0603958
R10163 dvdd dvdd.n882 0.0603958
R10164 dvdd dvdd.n881 0.0603958
R10165 dvdd.n862 dvdd 0.0603958
R10166 dvdd.n962 dvdd 0.0603958
R10167 dvdd.n973 dvdd 0.0603958
R10168 dvdd dvdd.n951 0.0603958
R10169 dvdd dvdd.n980 0.0603958
R10170 dvdd.n981 dvdd 0.0603958
R10171 dvdd.n949 dvdd 0.0603958
R10172 dvdd dvdd.n948 0.0603958
R10173 dvdd.n989 dvdd 0.0603958
R10174 dvdd.n990 dvdd 0.0603958
R10175 dvdd.n995 dvdd 0.0603958
R10176 dvdd.n1035 dvdd 0.0603958
R10177 dvdd.n1037 dvdd 0.0603958
R10178 dvdd dvdd.n1050 0.0603958
R10179 dvdd.n1051 dvdd 0.0603958
R10180 dvdd.n1097 dvdd 0.0603958
R10181 dvdd dvdd.n1096 0.0603958
R10182 dvdd dvdd.n1090 0.0603958
R10183 dvdd.n1084 dvdd 0.0603958
R10184 dvdd.n1058 dvdd 0.0603958
R10185 dvdd.n1060 dvdd 0.0603958
R10186 dvdd.n1073 dvdd 0.0603958
R10187 dvdd dvdd.n1072 0.0603958
R10188 dvdd.n1067 dvdd 0.0603958
R10189 dvdd dvdd.n1186 0.0603958
R10190 dvdd.n1182 dvdd 0.0603958
R10191 dvdd.n1176 dvdd 0.0603958
R10192 dvdd dvdd.n1175 0.0603958
R10193 dvdd.n1103 dvdd 0.0603958
R10194 dvdd.n1106 dvdd 0.0603958
R10195 dvdd.n1108 dvdd 0.0603958
R10196 dvdd.n1158 dvdd 0.0603958
R10197 dvdd.n1142 dvdd 0.0603958
R10198 dvdd.n1140 dvdd 0.0603958
R10199 dvdd.n1137 dvdd 0.0603958
R10200 dvdd dvdd.n1136 0.0603958
R10201 dvdd.n1265 dvdd 0.0603958
R10202 dvdd.n1269 dvdd 0.0603958
R10203 dvdd dvdd.n1252 0.0603958
R10204 dvdd.n1285 dvdd 0.0603958
R10205 dvdd.n1286 dvdd 0.0603958
R10206 dvdd dvdd.n1242 0.0603958
R10207 dvdd dvdd.n1238 0.0603958
R10208 dvdd.n1293 dvdd 0.0603958
R10209 dvdd dvdd.n1222 0.0603958
R10210 dvdd dvdd.n1323 0.0603958
R10211 dvdd.n1324 dvdd 0.0603958
R10212 dvdd.n1384 dvdd 0.0603958
R10213 dvdd dvdd.n1383 0.0603958
R10214 dvdd dvdd.n1382 0.0603958
R10215 dvdd.n1382 dvdd 0.0603958
R10216 dvdd.n1379 dvdd 0.0603958
R10217 dvdd dvdd.n1328 0.0603958
R10218 dvdd.n1332 dvdd 0.0603958
R10219 dvdd.n1364 dvdd 0.0603958
R10220 dvdd.n1360 dvdd 0.0603958
R10221 dvdd dvdd.n1480 0.0603958
R10222 dvdd.n1217 dvdd 0.0603958
R10223 dvdd.n1458 dvdd 0.0603958
R10224 dvdd dvdd.n1457 0.0603958
R10225 dvdd.n1437 dvdd 0.0603958
R10226 dvdd dvdd.n1435 0.0603958
R10227 dvdd.n1410 dvdd 0.0603958
R10228 dvdd.n1423 dvdd 0.0603958
R10229 dvdd dvdd.n1543 0.0603958
R10230 dvdd dvdd.n1541 0.0603958
R10231 dvdd.n1560 dvdd 0.0603958
R10232 dvdd dvdd.n1537 0.0603958
R10233 dvdd dvdd.n1535 0.0603958
R10234 dvdd.n1579 dvdd 0.0603958
R10235 dvdd.n1580 dvdd 0.0603958
R10236 dvdd.n1591 dvdd 0.0603958
R10237 dvdd dvdd.n1522 0.0603958
R10238 dvdd.n1598 dvdd 0.0603958
R10239 dvdd.n1603 dvdd 0.0603958
R10240 dvdd.n1605 dvdd 0.0603958
R10241 dvdd dvdd.n1511 0.0603958
R10242 dvdd.n1614 dvdd 0.0603958
R10243 dvdd.n1681 dvdd 0.0603958
R10244 dvdd dvdd.n1680 0.0603958
R10245 dvdd.n1677 dvdd 0.0603958
R10246 dvdd dvdd.n1671 0.0603958
R10247 dvdd.n1639 dvdd 0.0603958
R10248 dvdd.n1651 dvdd 0.0603958
R10249 dvdd.n1500 dvdd 0.0603958
R10250 dvdd.n1686 dvdd 0.0603958
R10251 dvdd dvdd.n1755 0.0603958
R10252 dvdd.n1755 dvdd 0.0603958
R10253 dvdd.n1752 dvdd 0.0603958
R10254 dvdd dvdd.n1751 0.0603958
R10255 dvdd.n1841 dvdd 0.0603958
R10256 dvdd.n1845 dvdd 0.0603958
R10257 dvdd.n1846 dvdd 0.0603958
R10258 dvdd.n1855 dvdd 0.0603958
R10259 dvdd.n1859 dvdd 0.0603958
R10260 dvdd.n1870 dvdd 0.0603958
R10261 dvdd.n1877 dvdd 0.0603958
R10262 dvdd dvdd.n1812 0.0603958
R10263 dvdd.n1915 dvdd 0.0603958
R10264 dvdd.n1916 dvdd 0.0603958
R10265 dvdd.n1926 dvdd 0.0603958
R10266 dvdd.n1987 dvdd 0.0603958
R10267 dvdd.n1986 dvdd 0.0603958
R10268 dvdd.n1983 dvdd 0.0603958
R10269 dvdd.n1979 dvdd 0.0603958
R10270 dvdd.n2079 dvdd 0.0603958
R10271 dvdd dvdd.n2078 0.0603958
R10272 dvdd.n2078 dvdd 0.0603958
R10273 dvdd.n2073 dvdd 0.0603958
R10274 dvdd.n2066 dvdd 0.0603958
R10275 dvdd dvdd.n2064 0.0603958
R10276 dvdd dvdd.n2039 0.0603958
R10277 dvdd.n2035 dvdd 0.0603958
R10278 dvdd.n2029 dvdd 0.0603958
R10279 dvdd dvdd.n2028 0.0603958
R10280 dvdd.n2244 dvdd 0.0603958
R10281 dvdd.n2247 dvdd 0.0603958
R10282 dvdd.n2270 dvdd 0.0603958
R10283 dvdd.n2276 dvdd 0.0603958
R10284 dvdd.n2319 dvdd 0.0603958
R10285 dvdd.n2320 dvdd 0.0603958
R10286 dvdd.n2329 dvdd 0.0603958
R10287 dvdd.n2330 dvdd 0.0603958
R10288 dvdd.n2118 dvdd 0.0603958
R10289 dvdd dvdd.n2117 0.0603958
R10290 dvdd dvdd.n2114 0.0603958
R10291 dvdd dvdd.n2343 0.0603958
R10292 dvdd.n2344 dvdd 0.0603958
R10293 dvdd.n2161 dvdd 0.0603958
R10294 dvdd dvdd.n2149 0.0603958
R10295 dvdd.n2225 dvdd 0.0603958
R10296 dvdd dvdd.n2222 0.0603958
R10297 dvdd.n2200 dvdd 0.0603958
R10298 dvdd dvdd.n2187 0.0603958
R10299 dvdd.n2420 dvdd 0.0603958
R10300 dvdd.n2423 dvdd 0.0603958
R10301 dvdd.n2424 dvdd 0.0603958
R10302 dvdd dvdd.n2406 0.0603958
R10303 dvdd.n2451 dvdd 0.0603958
R10304 dvdd.n2463 dvdd 0.0603958
R10305 dvdd.n2479 dvdd 0.0603958
R10306 dvdd dvdd.n2390 0.0603958
R10307 dvdd.n2501 dvdd 0.0603958
R10308 dvdd.n2553 dvdd 0.0603958
R10309 dvdd dvdd.n2552 0.0603958
R10310 dvdd dvdd.n2509 0.0603958
R10311 dvdd.n2515 dvdd 0.0603958
R10312 dvdd.n2534 dvdd 0.0603958
R10313 dvdd dvdd.n2533 0.0603958
R10314 dvdd.n2527 dvdd 0.0603958
R10315 dvdd.n2637 dvdd 0.0603958
R10316 dvdd dvdd.n2636 0.0603958
R10317 dvdd dvdd.n2383 0.0603958
R10318 dvdd.n2631 dvdd 0.0603958
R10319 dvdd dvdd.n2622 0.0603958
R10320 dvdd.n2619 dvdd 0.0603958
R10321 dvdd dvdd.n2618 0.0603958
R10322 dvdd dvdd.n2566 0.0603958
R10323 dvdd.n2611 dvdd 0.0603958
R10324 dvdd dvdd.n2610 0.0603958
R10325 dvdd.n2575 dvdd 0.0603958
R10326 dvdd.n2598 dvdd 0.0603958
R10327 dvdd.n2594 dvdd 0.0603958
R10328 dvdd dvdd.n2593 0.0603958
R10329 dvdd.n2922 dvdd 0.0603958
R10330 dvdd.n3076 dvdd 0.0603958
R10331 dvdd.n3019 dvdd 0.0603958
R10332 dvdd.n2855 dvdd 0.0603958
R10333 dvdd.n2865 dvdd 0.0603958
R10334 dvdd.n200 dvdd.n73 0.0574697
R10335 dvdd.n341 dvdd.n330 0.0574697
R10336 dvdd.n897 dvdd.n613 0.0574697
R10337 dvdd.n1188 dvdd.n914 0.0574697
R10338 dvdd.n1472 dvdd.n1203 0.0574697
R10339 dvdd.n1771 dvdd.n1487 0.0574697
R10340 dvdd.n1800 dvdd.n1788 0.0574697
R10341 dvdd.n2098 dvdd.n2090 0.0574697
R10342 dvdd.n2372 dvdd.n2360 0.0574697
R10343 dvdd dvdd.n915 0.0538854
R10344 dvdd dvdd.n2361 0.0538854
R10345 dvdd.n778 dvdd.n777 0.0512937
R10346 dvdd.n205 dvdd.n198 0.0499792
R10347 dvdd.n346 dvdd.n337 0.0499792
R10348 dvdd.n902 dvdd.n901 0.0499792
R10349 dvdd.n1193 dvdd.n1192 0.0499792
R10350 dvdd.n1477 dvdd.n1476 0.0499792
R10351 dvdd.n1776 dvdd.n1775 0.0499792
R10352 dvdd.n2103 dvdd.n2102 0.0499792
R10353 dvdd.n2377 dvdd.n2368 0.0499792
R10354 dvdd.n320 dvdd.n74 0.0447708
R10355 dvdd.n333 dvdd.n331 0.0447708
R10356 dvdd.n616 dvdd.n614 0.0447708
R10357 dvdd.n917 dvdd.n915 0.0447708
R10358 dvdd.n1206 dvdd.n1204 0.0447708
R10359 dvdd.n1490 dvdd.n1488 0.0447708
R10360 dvdd.n1791 dvdd.n1789 0.0447708
R10361 dvdd.n2093 dvdd.n2091 0.0447708
R10362 dvdd.n2363 dvdd.n2361 0.0447708
R10363 dvdd.n325 dvdd.n75 0.0410405
R10364 dvdd.n203 dvdd.n201 0.0410405
R10365 dvdd.n608 dvdd.n332 0.0410405
R10366 dvdd.n344 dvdd.n342 0.0410405
R10367 dvdd.n909 dvdd.n615 0.0410405
R10368 dvdd.n899 dvdd.n898 0.0410405
R10369 dvdd.n1198 dvdd.n916 0.0410405
R10370 dvdd.n1190 dvdd.n1189 0.0410405
R10371 dvdd.n1482 dvdd.n1205 0.0410405
R10372 dvdd.n1474 dvdd.n1473 0.0410405
R10373 dvdd.n1783 dvdd.n1489 0.0410405
R10374 dvdd.n1773 dvdd.n1772 0.0410405
R10375 dvdd.n2085 dvdd.n1790 0.0410405
R10376 dvdd.n1803 dvdd.n1801 0.0410405
R10377 dvdd.n2355 dvdd.n2092 0.0410405
R10378 dvdd.n2100 dvdd.n2099 0.0410405
R10379 dvdd.n2643 dvdd.n2362 0.0410405
R10380 dvdd.n2375 dvdd.n2373 0.0410405
R10381 dvdd.n607 dvdd.n333 0.0395625
R10382 dvdd.n908 dvdd.n616 0.0395625
R10383 dvdd.n1197 dvdd.n917 0.0395625
R10384 dvdd.n1481 dvdd.n1206 0.0395625
R10385 dvdd.n1782 dvdd.n1490 0.0395625
R10386 dvdd.n2084 dvdd.n1791 0.0395625
R10387 dvdd.n2354 dvdd.n2093 0.0395625
R10388 dvdd.n2642 dvdd.n2363 0.0395625
R10389 dvdd dvdd.n3093 0.0377807
R10390 dvdd.n2762 dvdd 0.0377807
R10391 dvdd dvdd.n2765 0.0377807
R10392 dvdd.n2766 dvdd 0.0377807
R10393 dvdd dvdd.n2769 0.0377807
R10394 dvdd.n2770 dvdd 0.0377807
R10395 dvdd dvdd.n2773 0.0377807
R10396 dvdd.n2774 dvdd 0.0377807
R10397 dvdd dvdd.n2777 0.0377807
R10398 dvdd.n2778 dvdd 0.0377807
R10399 dvdd dvdd.n2781 0.0377807
R10400 dvdd.n2782 dvdd 0.0377807
R10401 dvdd dvdd.n2785 0.0377807
R10402 dvdd.n2786 dvdd 0.0377807
R10403 dvdd dvdd.n2789 0.0377807
R10404 dvdd.n2790 dvdd 0.0377807
R10405 dvdd dvdd.n2793 0.0377807
R10406 dvdd.n2794 dvdd 0.0377807
R10407 dvdd dvdd.n2797 0.0377807
R10408 dvdd.n2798 dvdd 0.0377807
R10409 dvdd dvdd.n2801 0.0377807
R10410 dvdd.n2756 dvdd 0.0377807
R10411 dvdd.n2753 dvdd 0.0377807
R10412 dvdd.n2752 dvdd 0.0377807
R10413 dvdd.n2749 dvdd 0.0377807
R10414 dvdd.n2748 dvdd 0.0377807
R10415 dvdd.n2745 dvdd 0.0377807
R10416 dvdd.n2744 dvdd 0.0377807
R10417 dvdd.n2741 dvdd 0.0377807
R10418 dvdd.n2740 dvdd 0.0377807
R10419 dvdd.n2737 dvdd 0.0377807
R10420 dvdd.n2736 dvdd 0.0377807
R10421 dvdd.n2733 dvdd 0.0377807
R10422 dvdd.n2732 dvdd 0.0377807
R10423 dvdd.n2729 dvdd 0.0377807
R10424 dvdd.n2728 dvdd 0.0377807
R10425 dvdd.n2725 dvdd 0.0377807
R10426 dvdd.n2724 dvdd 0.0377807
R10427 dvdd.n2721 dvdd 0.0377807
R10428 dvdd.n2720 dvdd 0.0377807
R10429 dvdd.n2717 dvdd 0.0377807
R10430 dvdd.n202 dvdd.n198 0.0343542
R10431 dvdd.n343 dvdd.n337 0.0343542
R10432 dvdd.n902 dvdd.n622 0.0343542
R10433 dvdd.n1193 dvdd.n924 0.0343542
R10434 dvdd.n1477 dvdd.n1210 0.0343542
R10435 dvdd.n1776 dvdd.n1496 0.0343542
R10436 dvdd.n1802 dvdd.n1797 0.0343542
R10437 dvdd.n2103 dvdd.n2096 0.0343542
R10438 dvdd.n2374 dvdd.n2368 0.0343542
R10439 dvdd.n520 dvdd 0.0330521
R10440 dvdd.n1185 dvdd 0.0330521
R10441 dvdd.n1266 dvdd 0.0330521
R10442 dvdd.n1286 dvdd 0.0330521
R10443 dvdd.n1224 dvdd 0.0330521
R10444 dvdd.n1436 dvdd 0.0330521
R10445 dvdd.n1422 dvdd 0.0330521
R10446 dvdd dvdd.n1845 0.0330521
R10447 dvdd dvdd.n1914 0.0330521
R10448 dvdd.n2027 dvdd 0.0330521
R10449 dvdd dvdd.n2423 0.0330521
R10450 dvdd dvdd.n2502 0.0330521
R10451 dvdd.n170 dvdd 0.03175
R10452 dvdd.n155 dvdd 0.03175
R10453 dvdd dvdd.n284 0.03175
R10454 dvdd dvdd.n285 0.03175
R10455 dvdd.n279 dvdd 0.03175
R10456 dvdd.n278 dvdd 0.03175
R10457 dvdd.n385 dvdd 0.03175
R10458 dvdd dvdd.n412 0.03175
R10459 dvdd.n413 dvdd 0.03175
R10460 dvdd.n522 dvdd 0.03175
R10461 dvdd.n595 dvdd 0.03175
R10462 dvdd.n594 dvdd 0.03175
R10463 dvdd dvdd.n665 0.03175
R10464 dvdd.n692 dvdd 0.03175
R10465 dvdd.n811 dvdd 0.03175
R10466 dvdd.n790 dvdd 0.03175
R10467 dvdd.n895 dvdd 0.03175
R10468 dvdd.n883 dvdd 0.03175
R10469 dvdd.n882 dvdd 0.03175
R10470 dvdd dvdd.n989 0.03175
R10471 dvdd.n990 dvdd 0.03175
R10472 dvdd dvdd.n1051 0.03175
R10473 dvdd.n1097 dvdd 0.03175
R10474 dvdd dvdd.n1058 0.03175
R10475 dvdd.n1073 dvdd 0.03175
R10476 dvdd.n1176 dvdd 0.03175
R10477 dvdd.n1137 dvdd 0.03175
R10478 dvdd dvdd.n1285 0.03175
R10479 dvdd.n1238 dvdd 0.03175
R10480 dvdd.n1384 dvdd 0.03175
R10481 dvdd.n1383 dvdd 0.03175
R10482 dvdd dvdd.n1217 0.03175
R10483 dvdd.n1458 dvdd 0.03175
R10484 dvdd.n1543 dvdd 0.03175
R10485 dvdd dvdd.n1579 0.03175
R10486 dvdd.n1681 dvdd 0.03175
R10487 dvdd.n1680 dvdd 0.03175
R10488 dvdd dvdd.n1500 0.03175
R10489 dvdd.n1752 dvdd 0.03175
R10490 dvdd.n1841 dvdd 0.03175
R10491 dvdd.n1855 dvdd 0.03175
R10492 dvdd dvdd.n1926 0.03175
R10493 dvdd.n2079 dvdd 0.03175
R10494 dvdd.n2066 dvdd 0.03175
R10495 dvdd.n2244 dvdd 0.03175
R10496 dvdd.n2266 dvdd 0.03175
R10497 dvdd dvdd.n2319 0.03175
R10498 dvdd dvdd.n2149 0.03175
R10499 dvdd.n2225 dvdd 0.03175
R10500 dvdd.n2420 dvdd 0.03175
R10501 dvdd dvdd.n2450 0.03175
R10502 dvdd.n2553 dvdd 0.03175
R10503 dvdd.n2534 dvdd 0.03175
R10504 dvdd.n2637 dvdd 0.03175
R10505 dvdd.n2622 dvdd 0.03175
R10506 dvdd.n2611 dvdd 0.03175
R10507 dvdd dvdd.n2575 0.03175
R10508 dvdd.n2594 dvdd 0.03175
R10509 dvdd.n2645 dvdd.n2360 0.0292489
R10510 dvdd.n2372 dvdd.n2359 0.0292489
R10511 dvdd.n2357 dvdd.n2090 0.0292489
R10512 dvdd.n2098 dvdd.n2089 0.0292489
R10513 dvdd.n2087 dvdd.n1788 0.0292489
R10514 dvdd.n1800 dvdd.n1787 0.0292489
R10515 dvdd.n1785 dvdd.n1487 0.0292489
R10516 dvdd.n1771 dvdd.n1486 0.0292489
R10517 dvdd.n1484 dvdd.n1203 0.0292489
R10518 dvdd.n1472 dvdd.n1202 0.0292489
R10519 dvdd.n1200 dvdd.n914 0.0292489
R10520 dvdd.n1188 dvdd.n913 0.0292489
R10521 dvdd.n911 dvdd.n613 0.0292489
R10522 dvdd.n897 dvdd.n612 0.0292489
R10523 dvdd.n610 dvdd.n330 0.0292489
R10524 dvdd.n341 dvdd.n329 0.0292489
R10525 dvdd.n327 dvdd.n73 0.0292489
R10526 dvdd.n200 dvdd.n72 0.0292489
R10527 dvdd dvdd.n2523 0.0291458
R10528 dvdd dvdd.n2378 0.0291458
R10529 dvdd.n1805 dvdd 0.0278438
R10530 dvdd.n924 dvdd 0.0265417
R10531 dvdd.n1210 dvdd 0.0265417
R10532 dvdd dvdd.n1284 0.0252396
R10533 dvdd.n3115 dvdd.n3114 0.0243462
R10534 dvdd.n3105 dvdd.n3100 0.0243462
R10535 dvdd.n810 dvdd 0.0239375
R10536 dvdd.n774 dvdd 0.0239375
R10537 dvdd.n973 dvdd 0.0239375
R10538 dvdd.n1091 dvdd 0.0239375
R10539 dvdd.n1090 dvdd 0.0239375
R10540 dvdd.n1169 dvdd 0.0239375
R10541 dvdd dvdd.n1269 0.0239375
R10542 dvdd dvdd.n1625 0.0239375
R10543 dvdd dvdd.n1686 0.0239375
R10544 dvdd.n1872 dvdd 0.0239375
R10545 dvdd.n2035 dvdd 0.0239375
R10546 dvdd.n190 dvdd 0.0226354
R10547 dvdd dvdd.n89 0.0226354
R10548 dvdd.n133 dvdd 0.0226354
R10549 dvdd.n115 dvdd 0.0226354
R10550 dvdd.n112 dvdd 0.0226354
R10551 dvdd.n286 dvdd 0.0226354
R10552 dvdd.n298 dvdd 0.0226354
R10553 dvdd.n320 dvdd 0.0226354
R10554 dvdd dvdd.n215 0.0226354
R10555 dvdd.n259 dvdd 0.0226354
R10556 dvdd.n239 dvdd 0.0226354
R10557 dvdd.n231 dvdd 0.0226354
R10558 dvdd.n405 dvdd 0.0226354
R10559 dvdd dvdd.n434 0.0226354
R10560 dvdd dvdd.n457 0.0226354
R10561 dvdd.n509 dvdd 0.0226354
R10562 dvdd.n508 dvdd 0.0226354
R10563 dvdd dvdd.n473 0.0226354
R10564 dvdd.n583 dvdd 0.0226354
R10565 dvdd dvdd.n533 0.0226354
R10566 dvdd dvdd.n538 0.0226354
R10567 dvdd.n556 dvdd 0.0226354
R10568 dvdd dvdd.n673 0.0226354
R10569 dvdd.n674 dvdd 0.0226354
R10570 dvdd.n680 dvdd 0.0226354
R10571 dvdd dvdd.n702 0.0226354
R10572 dvdd.n724 dvdd 0.0226354
R10573 dvdd dvdd.n752 0.0226354
R10574 dvdd dvdd.n759 0.0226354
R10575 dvdd.n775 dvdd 0.0226354
R10576 dvdd.n887 dvdd 0.0226354
R10577 dvdd.n867 dvdd 0.0226354
R10578 dvdd.n845 dvdd 0.0226354
R10579 dvdd.n962 dvdd 0.0226354
R10580 dvdd dvdd.n972 0.0226354
R10581 dvdd dvdd.n988 0.0226354
R10582 dvdd.n1026 dvdd 0.0226354
R10583 dvdd dvdd.n1036 0.0226354
R10584 dvdd.n1037 dvdd 0.0226354
R10585 dvdd dvdd.n1044 0.0226354
R10586 dvdd.n1067 dvdd 0.0226354
R10587 dvdd dvdd.n926 0.0226354
R10588 dvdd.n1175 dvdd 0.0226354
R10589 dvdd dvdd.n1108 0.0226354
R10590 dvdd.n1161 dvdd 0.0226354
R10591 dvdd.n1145 dvdd 0.0226354
R10592 dvdd.n1142 dvdd 0.0226354
R10593 dvdd.n1131 dvdd 0.0226354
R10594 dvdd.n1253 dvdd 0.0226354
R10595 dvdd.n1252 dvdd 0.0226354
R10596 dvdd.n1313 dvdd 0.0226354
R10597 dvdd dvdd.n1324 0.0226354
R10598 dvdd dvdd.n1325 0.0226354
R10599 dvdd.n1379 dvdd 0.0226354
R10600 dvdd dvdd.n1332 0.0226354
R10601 dvdd.n1360 dvdd 0.0226354
R10602 dvdd.n1440 dvdd 0.0226354
R10603 dvdd dvdd.n1407 0.0226354
R10604 dvdd dvdd.n1410 0.0226354
R10605 dvdd dvdd.n1411 0.0226354
R10606 dvdd dvdd.n1559 0.0226354
R10607 dvdd.n1560 dvdd 0.0226354
R10608 dvdd.n1565 dvdd 0.0226354
R10609 dvdd.n1537 dvdd 0.0226354
R10610 dvdd dvdd.n1578 0.0226354
R10611 dvdd dvdd.n1580 0.0226354
R10612 dvdd dvdd.n1590 0.0226354
R10613 dvdd.n1591 dvdd 0.0226354
R10614 dvdd.n1522 dvdd 0.0226354
R10615 dvdd dvdd.n1613 0.0226354
R10616 dvdd dvdd.n1634 0.0226354
R10617 dvdd.n1654 dvdd 0.0226354
R10618 dvdd.n1751 dvdd 0.0226354
R10619 dvdd.n1716 dvdd 0.0226354
R10620 dvdd dvdd.n1854 0.0226354
R10621 dvdd dvdd.n1866 0.0226354
R10622 dvdd.n1867 dvdd 0.0226354
R10623 dvdd.n1909 dvdd 0.0226354
R10624 dvdd dvdd.n1915 0.0226354
R10625 dvdd dvdd.n1925 0.0226354
R10626 dvdd.n1982 dvdd 0.0226354
R10627 dvdd.n1979 dvdd 0.0226354
R10628 dvdd dvdd.n1797 0.0226354
R10629 dvdd dvdd.n1807 0.0226354
R10630 dvdd.n2044 dvdd 0.0226354
R10631 dvdd.n2040 dvdd 0.0226354
R10632 dvdd.n2039 dvdd 0.0226354
R10633 dvdd.n2038 dvdd 0.0226354
R10634 dvdd dvdd.n2265 0.0226354
R10635 dvdd.n2272 dvdd 0.0226354
R10636 dvdd dvdd.n2288 0.0226354
R10637 dvdd.n2295 dvdd 0.0226354
R10638 dvdd.n2310 dvdd 0.0226354
R10639 dvdd dvdd.n2328 0.0226354
R10640 dvdd dvdd.n2329 0.0226354
R10641 dvdd.n2330 dvdd 0.0226354
R10642 dvdd.n2339 dvdd 0.0226354
R10643 dvdd.n2349 dvdd 0.0226354
R10644 dvdd dvdd.n2160 0.0226354
R10645 dvdd.n2161 dvdd 0.0226354
R10646 dvdd.n2208 dvdd 0.0226354
R10647 dvdd.n2205 dvdd 0.0226354
R10648 dvdd.n2203 dvdd 0.0226354
R10649 dvdd.n2200 dvdd 0.0226354
R10650 dvdd.n2438 dvdd 0.0226354
R10651 dvdd.n2444 dvdd 0.0226354
R10652 dvdd dvdd.n2457 0.0226354
R10653 dvdd.n2463 dvdd 0.0226354
R10654 dvdd.n2471 dvdd 0.0226354
R10655 dvdd dvdd.n2486 0.0226354
R10656 dvdd.n2488 dvdd 0.0226354
R10657 dvdd.n2498 dvdd 0.0226354
R10658 dvdd dvdd.n2509 0.0226354
R10659 dvdd.n2527 dvdd 0.0226354
R10660 dvdd dvdd.n2383 0.0226354
R10661 dvdd.n2631 dvdd 0.0226354
R10662 dvdd.n2623 dvdd 0.0226354
R10663 dvdd.n2619 dvdd 0.0226354
R10664 dvdd dvdd.n2574 0.0226354
R10665 dvdd.n2597 dvdd 0.0226354
R10666 dvdd dvdd.n2579 0.0226354
R10667 dvdd.n2918 dvdd 0.0226354
R10668 dvdd dvdd.n2928 0.0226354
R10669 dvdd.n3072 dvdd 0.0226354
R10670 dvdd dvdd.n3082 0.0226354
R10671 dvdd.n3015 dvdd 0.0226354
R10672 dvdd dvdd.n3025 0.0226354
R10673 dvdd.n2852 dvdd 0.0226354
R10674 dvdd.n2861 dvdd 0.0226354
R10675 dvdd dvdd.n2871 0.0226354
R10676 dvdd dvdd.n464 0.0213333
R10677 dvdd dvdd.n481 0.0213333
R10678 dvdd.n598 dvdd 0.0213333
R10679 dvdd.n783 dvdd 0.0213333
R10680 dvdd dvdd.n981 0.0213333
R10681 dvdd.n948 dvdd 0.0213333
R10682 dvdd.n1076 dvdd 0.0213333
R10683 dvdd dvdd.n1106 0.0213333
R10684 dvdd dvdd.n1318 0.0213333
R10685 dvdd.n1481 dvdd 0.0213333
R10686 dvdd.n1462 dvdd 0.0213333
R10687 dvdd.n1672 dvdd 0.0213333
R10688 dvdd.n1643 dvdd 0.0213333
R10689 dvdd.n1762 dvdd 0.0213333
R10690 dvdd.n1756 dvdd 0.0213333
R10691 dvdd.n2537 dvdd 0.0213333
R10692 dvdd dvdd.n1207 0.0200312
R10693 dvdd dvdd.n76 0.0187292
R10694 dvdd dvdd.n918 0.0187292
R10695 dvdd.n324 dvdd 0.0174271
R10696 dvdd dvdd.n1488 0.016125
R10697 dvdd dvdd.n2091 0.016125
R10698 dvdd.n901 dvdd 0.0109167
R10699 dvdd.n1192 dvdd 0.0109167
R10700 dvdd dvdd.n1805 0.0109167
R10701 dvdd dvdd.n2377 0.0109167
R10702 dvdd.n323 dvdd.n76 0.00310417
R10703 dvdd.n606 dvdd.n334 0.00310417
R10704 dvdd.n907 dvdd.n617 0.00310417
R10705 dvdd.n1196 dvdd.n918 0.00310417
R10706 dvdd.n1480 dvdd.n1207 0.00310417
R10707 dvdd.n1781 dvdd.n1491 0.00310417
R10708 dvdd.n2083 dvdd.n1792 0.00310417
R10709 dvdd.n2353 dvdd.n2094 0.00310417
R10710 dvdd.n2641 dvdd.n2364 0.00310417
R10711 por_ana_0.comparator_1.n0.n2 por_ana_0.comparator_1.n0.t7 227.651
R10712 por_ana_0.comparator_1.n0.n2 por_ana_0.comparator_1.n0.t5 227.173
R10713 por_ana_0.comparator_1.n0.n0 por_ana_0.comparator_1.n0.t8 224.037
R10714 por_ana_0.comparator_1.n0.n0 por_ana_0.comparator_1.n0.t6 223.559
R10715 por_ana_0.comparator_1.n0 por_ana_0.comparator_1.n0.n1 205.605
R10716 por_ana_0.comparator_1.n0 por_ana_0.comparator_1.n0.t2 96.5813
R10717 por_ana_0.comparator_1.n0 por_ana_0.comparator_1.n0.n3 70.9612
R10718 por_ana_0.comparator_1.n0.n1 por_ana_0.comparator_1.n0.t0 27.6955
R10719 por_ana_0.comparator_1.n0.n1 por_ana_0.comparator_1.n0.t1 27.6955
R10720 por_ana_0.comparator_1.n0.n3 por_ana_0.comparator_1.n0.t3 16.5305
R10721 por_ana_0.comparator_1.n0.n3 por_ana_0.comparator_1.n0.t4 16.5305
R10722 por_ana_0.comparator_1.n0.n0 por_ana_0.comparator_1.n0.n2 14.4688
R10723 por_ana_0.comparator_1.n0 por_ana_0.comparator_1.n0.n0 10.4432
R10724 por_ana_0.comparator_1.n1.n0 por_ana_0.comparator_1.n1.t16 227.657
R10725 por_ana_0.comparator_1.n1.n0 por_ana_0.comparator_1.n1.t11 227.173
R10726 por_ana_0.comparator_1.n1.n0 por_ana_0.comparator_1.n1.t5 227.173
R10727 por_ana_0.comparator_1.n1.n0 por_ana_0.comparator_1.n1.t19 227.173
R10728 por_ana_0.comparator_1.n1.n0 por_ana_0.comparator_1.n1.t12 227.173
R10729 por_ana_0.comparator_1.n1.n0 por_ana_0.comparator_1.n1.t6 227.173
R10730 por_ana_0.comparator_1.n1.n0 por_ana_0.comparator_1.n1.t18 227.173
R10731 por_ana_0.comparator_1.n1.n0 por_ana_0.comparator_1.n1.t8 227.173
R10732 por_ana_0.comparator_1.n1.n1 por_ana_0.comparator_1.n1.t14 224.042
R10733 por_ana_0.comparator_1.n1.n1 por_ana_0.comparator_1.n1.t9 223.559
R10734 por_ana_0.comparator_1.n1.n1 por_ana_0.comparator_1.n1.t17 223.559
R10735 por_ana_0.comparator_1.n1.n1 por_ana_0.comparator_1.n1.t15 223.559
R10736 por_ana_0.comparator_1.n1.n1 por_ana_0.comparator_1.n1.t10 223.559
R10737 por_ana_0.comparator_1.n1.n1 por_ana_0.comparator_1.n1.t4 223.559
R10738 por_ana_0.comparator_1.n1.n1 por_ana_0.comparator_1.n1.t13 223.559
R10739 por_ana_0.comparator_1.n1.n1 por_ana_0.comparator_1.n1.t7 223.559
R10740 por_ana_0.comparator_1.n1.n5 por_ana_0.comparator_1.n1.n4 204.31
R10741 por_ana_0.comparator_1.n1.n3 por_ana_0.comparator_1.n1.n2 71.6326
R10742 por_ana_0.comparator_1.n1.n5 por_ana_0.comparator_1.n1.t0 27.6955
R10743 por_ana_0.comparator_1.n1.t1 por_ana_0.comparator_1.n1.n5 27.6955
R10744 por_ana_0.comparator_1.n1.n2 por_ana_0.comparator_1.n1.t3 16.5305
R10745 por_ana_0.comparator_1.n1.n2 por_ana_0.comparator_1.n1.t2 16.5305
R10746 por_ana_0.comparator_1.n1.n4 por_ana_0.comparator_1.n1.n0 8.13016
R10747 por_ana_0.comparator_1.n1.n3 por_ana_0.comparator_1.n1.n1 7.46509
R10748 por_ana_0.comparator_1.n1.n4 por_ana_0.comparator_1.n1.n3 4.52617
R10749 dvss.n4825 dvss.n1237 246424
R10750 dvss.n4813 dvss.n1237 246424
R10751 dvss.n4813 dvss.n1238 246418
R10752 dvss.n4825 dvss.n1238 246418
R10753 dvss.n1687 dvss.n1686 198880
R10754 dvss.n1572 dvss.n1571 198880
R10755 dvss.n1572 dvss.t1027 192115
R10756 dvss.t126 dvss.n1686 192115
R10757 dvss.n4824 dvss.n2296 86177
R10758 dvss.n7042 dvss.n7041 82533.9
R10759 dvss.n7039 dvss.n7017 78608.8
R10760 dvss.n7018 dvss.n7017 78608.8
R10761 dvss.n7039 dvss.n7023 78608.8
R10762 dvss.n7023 dvss.n7018 78608.8
R10763 dvss.n4812 dvss.n4811 58917.7
R10764 dvss.n6610 dvss.n6609 37915.2
R10765 dvss.n4824 dvss.n4823 26879.3
R10766 dvss.n6639 dvss.n6638 22284.8
R10767 dvss.n4814 dvss.n1235 16011.3
R10768 dvss.n4826 dvss.n1236 16010.9
R10769 dvss.n4827 dvss.n4826 16010.2
R10770 dvss.n4815 dvss.n4814 16007.9
R10771 dvss.n7020 dvss.n7002 12828.2
R10772 dvss.n7043 dvss.n7002 12828.2
R10773 dvss.n7020 dvss.n7016 12822.4
R10774 dvss.n7043 dvss.n7016 12822.4
R10775 dvss.n4799 dvss.n4797 12566.2
R10776 dvss.n435 dvss 12161.8
R10777 dvss.n4807 dvss.n237 11129.1
R10778 dvss.n4807 dvss.n4806 8961.68
R10779 dvss.n6986 dvss.n8 8941.81
R10780 dvss.n434 dvss.n278 8034.33
R10781 dvss.n5610 dvss.t665 8003.11
R10782 dvss.n6647 dvss.t1408 8003.11
R10783 dvss.t1099 dvss.n6949 8003.11
R10784 dvss.n6208 dvss.t2201 8003.11
R10785 dvss.t1003 dvss.n487 8003.11
R10786 dvss.t1121 dvss.n862 8003.11
R10787 dvss.t1496 dvss.n2105 8003.11
R10788 dvss.t1307 dvss.n1985 8003.11
R10789 dvss.t259 dvss.n1530 8003.11
R10790 dvss.t663 dvss.t671 7626.67
R10791 dvss.t669 dvss.t665 7626.67
R10792 dvss.t1414 dvss.t1412 7626.67
R10793 dvss.t1410 dvss.t1408 7626.67
R10794 dvss.t1103 dvss.t1105 7626.67
R10795 dvss.t1099 dvss.t1101 7626.67
R10796 dvss.t2203 dvss.t2205 7626.67
R10797 dvss.t2197 dvss.t2201 7626.67
R10798 dvss.t1005 dvss.t1001 7626.67
R10799 dvss.t1003 dvss.t999 7626.67
R10800 dvss.t1113 dvss.t1117 7626.67
R10801 dvss.t1121 dvss.t1115 7626.67
R10802 dvss.t1492 dvss.t1490 7626.67
R10803 dvss.t1496 dvss.t1488 7626.67
R10804 dvss.t1313 dvss.t1311 7626.67
R10805 dvss.t1307 dvss.t1309 7626.67
R10806 dvss.t265 dvss.t263 7626.67
R10807 dvss.t261 dvss.t259 7626.67
R10808 dvss.n4812 dvss.n4807 7609.27
R10809 dvss.n6811 dvss.n6810 6332.05
R10810 dvss.n6728 dvss.n111 6332.05
R10811 dvss.n5923 dvss.n5922 6332.05
R10812 dvss.n5997 dvss.n5996 6332.05
R10813 dvss.n5834 dvss.n840 6332.05
R10814 dvss.n5752 dvss.n874 6332.05
R10815 dvss.n2013 dvss.n2004 6332.05
R10816 dvss.n1649 dvss.n1648 6332.05
R10817 dvss.n6120 dvss.t1545 6153.5
R10818 dvss.n6861 dvss.t1513 6153.5
R10819 dvss.t1072 dvss.n11 6153.5
R10820 dvss.t40 dvss.n849 6153.5
R10821 dvss.n5731 dvss.t40 6153.5
R10822 dvss.n2017 dvss.t40 6153.5
R10823 dvss.n1506 dvss.t40 6153.5
R10824 dvss.t1456 dvss.n3265 6153.5
R10825 dvss.n6607 dvss.n335 5792.85
R10826 dvss.n6503 dvss.n6502 5772.37
R10827 dvss.n4825 dvss.n4824 5737.8
R10828 dvss.n6502 dvss.n8 5605.26
R10829 dvss.n435 dvss.n434 5502.51
R10830 dvss.n2295 dvss.n1239 5392.4
R10831 dvss.n7038 dvss.n7024 5107.58
R10832 dvss.n7036 dvss.n7024 5107.58
R10833 dvss.n7038 dvss.n7037 5107.58
R10834 dvss.n7037 dvss.n7036 5107.58
R10835 dvss.n6981 dvss.n11 5082
R10836 dvss.n6861 dvss.n6860 5082
R10837 dvss.n5989 dvss.n507 5082
R10838 dvss.n6715 dvss.n121 5082
R10839 dvss.n6716 dvss.n6715 5082
R10840 dvss.n6239 dvss.n507 5082
R10841 dvss.n6120 dvss.n6119 5082
R10842 dvss.n5822 dvss.n849 5082
R10843 dvss.n5732 dvss.n5731 5082
R10844 dvss.n2017 dvss.n2016 5082
R10845 dvss.n1652 dvss.n1506 5082
R10846 dvss dvss.t1784 4897.32
R10847 dvss dvss.t1794 4897.32
R10848 dvss.t1737 dvss 4888.89
R10849 dvss.t1860 dvss 4888.89
R10850 dvss dvss.t1734 4888.89
R10851 dvss.n6608 dvss.n6607 4826.37
R10852 dvss.n3197 dvss.n3196 4776.42
R10853 dvss.n6606 dvss.t334 4465.22
R10854 dvss.t1025 dvss.n1571 4455
R10855 dvss.n1687 dvss.t124 4455
R10856 dvss dvss.t1737 4408.43
R10857 dvss.t1784 dvss 4408.43
R10858 dvss.t1794 dvss 4408.43
R10859 dvss dvss.t1860 4408.43
R10860 dvss.t1734 dvss 4408.43
R10861 dvss.n419 dvss.n416 4160.18
R10862 dvss.n432 dvss.n416 4160.18
R10863 dvss.n419 dvss.n417 4160.18
R10864 dvss.n432 dvss.n417 4160.18
R10865 dvss.n3237 dvss.n3153 4092
R10866 dvss.n4855 dvss.n1231 3912.21
R10867 dvss.n4851 dvss.n1231 3912.21
R10868 dvss.n4851 dvss.n1229 3912.21
R10869 dvss.n4855 dvss.n1229 3912.21
R10870 dvss.t1773 dvss.t1765 3877.39
R10871 dvss.n6610 dvss.n278 3708.43
R10872 dvss.n2296 dvss.n2295 3614.09
R10873 dvss.n4804 dvss.n2306 3391.9
R10874 dvss.n4804 dvss.n2307 3391.9
R10875 dvss.n4800 dvss.n2307 3391.9
R10876 dvss.n4800 dvss.n2306 3391.9
R10877 dvss dvss.t1726 3363.22
R10878 dvss.n6607 dvss.n6606 3328.76
R10879 dvss.n1570 dvss.n1239 3302.54
R10880 dvss.n6638 dvss.n237 3196.46
R10881 dvss.t1694 dvss.t1776 3101.92
R10882 dvss.n6609 dvss.n6608 2962.09
R10883 dvss.n3907 dvss.n1132 2882.92
R10884 dvss.t1717 dvss 2857.47
R10885 dvss.t1897 dvss 2857.47
R10886 dvss dvss.n278 2800
R10887 dvss dvss.n6610 2763.24
R10888 dvss dvss.t1815 2570.88
R10889 dvss.t1697 dvss 2562.45
R10890 dvss dvss.t1743 2562.45
R10891 dvss.t1881 dvss.t1697 2326.44
R10892 dvss.t1815 dvss.t1746 2326.44
R10893 dvss.t1027 dvss.t1025 2310
R10894 dvss.t124 dvss.t126 2310
R10895 dvss.t520 dvss.t1087 2149.43
R10896 dvss.t1941 dvss 2090.42
R10897 dvss.t1844 dvss 2081.99
R10898 dvss.t1743 dvss 2081.99
R10899 dvss.t1746 dvss 2081.99
R10900 dvss.n1593 dvss.t1029 2079.65
R10901 dvss.n7042 dvss.t2099 2014.07
R10902 dvss.t1191 dvss.t1872 1963.98
R10903 dvss.t1386 dvss.t799 1888.12
R10904 dvss.n4821 dvss.n2297 1830.97
R10905 dvss.n4821 dvss.n2298 1830.97
R10906 dvss.n4810 dvss.n2298 1830.97
R10907 dvss.n4810 dvss.n2297 1830.97
R10908 dvss.n3291 dvss.n237 1808.4
R10909 dvss.n6606 dvss.t227 1808.05
R10910 dvss dvss.t1926 1795.4
R10911 dvss.t1076 dvss.t1078 1778.24
R10912 dvss.t1519 dvss.t1517 1778.24
R10913 dvss.t1462 dvss.t1464 1778.24
R10914 dvss.t1537 dvss.t1539 1778.24
R10915 dvss.t1535 dvss.t1545 1778.24
R10916 dvss.t662 dvss.t1014 1753.26
R10917 dvss.t621 dvss.t283 1753.26
R10918 dvss.t117 dvss.t307 1753.26
R10919 dvss dvss.t1720 1702.68
R10920 dvss dvss.t1729 1702.68
R10921 dvss dvss.t1797 1702.68
R10922 dvss dvss.t1688 1702.68
R10923 dvss.t1723 dvss 1702.68
R10924 dvss.t1825 dvss 1702.68
R10925 dvss dvss.t1863 1694.25
R10926 dvss dvss.t827 1681.61
R10927 dvss.n6949 dvss.t1078 1652.85
R10928 dvss.n6647 dvss.t1519 1652.85
R10929 dvss.t1462 dvss.n3153 1652.85
R10930 dvss.n5610 dvss.t1537 1652.85
R10931 dvss.n4797 dvss.n4796 1647.35
R10932 dvss.n4796 dvss.n4795 1647.35
R10933 dvss.n4795 dvss.n4794 1647.35
R10934 dvss.n4794 dvss.n4793 1647.35
R10935 dvss.n4793 dvss.n4792 1647.35
R10936 dvss.n4792 dvss.n4791 1647.35
R10937 dvss.n4791 dvss.n4790 1647.35
R10938 dvss.t1572 dvss 1626.82
R10939 dvss.n7021 dvss.t2021 1589.55
R10940 dvss.t1388 dvss.t299 1584.67
R10941 dvss.t475 dvss.t1439 1584.67
R10942 dvss.t919 dvss.t2004 1576.25
R10943 dvss.t2069 dvss.t792 1576.25
R10944 dvss.n2448 dvss.t1800 1550.96
R10945 dvss.t1926 dvss.t1717 1550.96
R10946 dvss.n4789 dvss.t1828 1550.96
R10947 dvss.n4316 dvss.t1894 1550.96
R10948 dvss.t829 dvss.t1749 1534.1
R10949 dvss.t1757 dvss.t553 1517.24
R10950 dvss.t1847 dvss 1424.52
R10951 dvss dvss.t1740 1424.52
R10952 dvss dvss.t1812 1424.52
R10953 dvss.n3196 dvss.n1132 1413.96
R10954 dvss dvss.t1875 1407.66
R10955 dvss dvss.t1700 1407.66
R10956 dvss.t1706 dvss 1407.66
R10957 dvss dvss.t1787 1407.66
R10958 dvss dvss.t1853 1407.66
R10959 dvss dvss.t1703 1407.66
R10960 dvss.t1034 dvss.t721 1399.23
R10961 dvss.t687 dvss.t1055 1399.23
R10962 dvss.t18 dvss.t356 1399.23
R10963 dvss.t2211 dvss.t1135 1399.23
R10964 dvss.t1428 dvss.t2233 1399.23
R10965 dvss.t21 dvss.t1284 1399.23
R10966 dvss.t2037 dvss.t900 1399.23
R10967 dvss.n6608 dvss.t62 1395.12
R10968 dvss.n6609 dvss.t1138 1376.81
R10969 dvss.t1685 dvss 1365.52
R10970 dvss.t369 dvss.t913 1348.66
R10971 dvss dvss.t2179 1340.23
R10972 dvss.t2 dvss 1340.23
R10973 dvss.t16 dvss.t1956 1323.37
R10974 dvss.t1781 dvss.t771 1323.37
R10975 dvss.t1820 dvss 1314.94
R10976 dvss dvss.t1951 1306.51
R10977 dvss dvss.t1401 1306.51
R10978 dvss.t1776 dvss 1306.51
R10979 dvss dvss.t1181 1297.56
R10980 dvss.n4790 dvss.t2121 1297.34
R10981 dvss dvss.t811 1280.53
R10982 dvss.n434 dvss.n433 1258.81
R10983 dvss.t1568 dvss.t428 1255.94
R10984 dvss.t285 dvss.t408 1255.94
R10985 dvss.t950 dvss.t1505 1255.94
R10986 dvss dvss.t929 1247.51
R10987 dvss.n2990 dvss.n2989 1198.25
R10988 dvss.n2743 dvss.n2742 1198.25
R10989 dvss.n3412 dvss.n3338 1198.25
R10990 dvss.n3759 dvss.n3758 1198.25
R10991 dvss.n3761 dvss.n3760 1198.25
R10992 dvss.n3906 dvss.n3905 1198.25
R10993 dvss.n3977 dvss.n3908 1198.25
R10994 dvss.n3629 dvss.n3628 1198.25
R10995 dvss.n4315 dvss.n2386 1198.25
R10996 dvss.n4736 dvss.n4545 1198.25
R10997 dvss.n5003 dvss.n5002 1198.25
R10998 dvss.n5003 dvss.n1228 1198.25
R10999 dvss.n5004 dvss.n5003 1198.25
R11000 dvss.n4266 dvss.n4193 1198.25
R11001 dvss.n4192 dvss.n4191 1198.25
R11002 dvss.n3125 dvss.n2305 1197.1
R11003 dvss.n2482 dvss.n2448 1197.02
R11004 dvss.n4677 dvss.n4593 1196.86
R11005 dvss.n2630 dvss.n2566 1194.5
R11006 dvss.n3124 dvss.n3123 1194.5
R11007 dvss.n2988 dvss.n2987 1194.5
R11008 dvss.n2846 dvss.n2845 1194.5
R11009 dvss.n3567 dvss.n3527 1194.5
R11010 dvss.n4384 dvss.n4316 1194.5
R11011 dvss.n4789 dvss.n4788 1194.5
R11012 dvss.n4050 dvss.n4049 1194.5
R11013 dvss.n2989 dvss.t1444 1180.08
R11014 dvss.n2742 dvss.t970 1180.08
R11015 dvss.n3527 dvss.t730 1180.08
R11016 dvss.n4049 dvss.t988 1180.08
R11017 dvss.n4491 dvss.t307 1180.08
R11018 dvss.n4491 dvss.n4490 1178.76
R11019 dvss.n4490 dvss.n2326 1139.2
R11020 dvss.t648 dvss.n335 1124.77
R11021 dvss.n433 dvss.t650 1124.77
R11022 dvss.t1273 dvss.t944 1112.64
R11023 dvss.t406 dvss.t917 1112.64
R11024 dvss.t964 dvss.t1289 1112.64
R11025 dvss.t952 dvss.t269 1112.64
R11026 dvss.t948 dvss.t1352 1112.64
R11027 dvss dvss.t412 1095.79
R11028 dvss.t1502 dvss.t1992 1095.79
R11029 dvss.t862 dvss 1095.79
R11030 dvss.t1091 dvss.t774 1095.79
R11031 dvss.t954 dvss 1095.79
R11032 dvss.t896 dvss 1078.93
R11033 dvss.t730 dvss.t2030 1078.93
R11034 dvss.t1107 dvss.t602 1070.5
R11035 dvss dvss.t1269 1070.5
R11036 dvss.t1281 dvss 1070.5
R11037 dvss.t1053 dvss 1062.07
R11038 dvss.t233 dvss.t227 1062.07
R11039 dvss.t229 dvss.t233 1062.07
R11040 dvss.t241 dvss.t229 1062.07
R11041 dvss.t235 dvss.t241 1062.07
R11042 dvss.t231 dvss.t235 1062.07
R11043 dvss.t243 dvss.t231 1062.07
R11044 dvss.t237 dvss.t243 1062.07
R11045 dvss.t251 dvss.t237 1062.07
R11046 dvss.t247 dvss.t251 1062.07
R11047 dvss.t253 dvss.t247 1062.07
R11048 dvss.t245 dvss.t239 1062.07
R11049 dvss.t239 dvss.t255 1062.07
R11050 dvss.t255 dvss.t249 1062.07
R11051 dvss.t249 dvss.t257 1062.07
R11052 dvss.t827 dvss.t821 1062.07
R11053 dvss.t821 dvss.t823 1062.07
R11054 dvss.t823 dvss.t825 1062.07
R11055 dvss dvss.t1963 1053.64
R11056 dvss dvss.t1356 1053.64
R11057 dvss.t1570 dvss 1045.21
R11058 dvss.t1217 dvss 1045.21
R11059 dvss.t722 dvss 1045.21
R11060 dvss.t1866 dvss 1036.78
R11061 dvss dvss.t742 1036.78
R11062 dvss.t1450 dvss.t2008 1036.78
R11063 dvss.t774 dvss.t1052 1036.78
R11064 dvss.t1452 dvss.t1317 1036.78
R11065 dvss dvss.t1507 1036.78
R11066 dvss.t541 dvss.t1058 1036.78
R11067 dvss dvss.t1416 1036.78
R11068 dvss dvss.t1265 1028.35
R11069 dvss dvss.t1169 1028.35
R11070 dvss dvss.t2153 1028.35
R11071 dvss.t283 dvss 1028.35
R11072 dvss dvss.t1452 1028.35
R11073 dvss.t1951 dvss 1019.92
R11074 dvss.t1770 dvss 1019.92
R11075 dvss.t673 dvss.t885 1019.92
R11076 dvss.t985 dvss 1019.92
R11077 dvss dvss.t1897 1019.92
R11078 dvss.t1765 dvss 1019.92
R11079 dvss.t426 dvss.t454 1011.49
R11080 dvss.t1878 dvss 1011.49
R11081 dvss.t1565 dvss 1011.49
R11082 dvss.t718 dvss.t1336 1003.07
R11083 dvss.t2028 dvss.t728 1003.07
R11084 dvss.t2010 dvss 1003.07
R11085 dvss.t320 dvss 986.207
R11086 dvss dvss.t930 986.207
R11087 dvss.t80 dvss.n4315 986.207
R11088 dvss.t257 dvss 986.207
R11089 dvss.t1999 dvss.t848 977.779
R11090 dvss.t166 dvss.t1959 969.35
R11091 dvss.t1251 dvss.t1276 960.92
R11092 dvss.t1833 dvss.t80 952.49
R11093 dvss.t825 dvss 948.277
R11094 dvss dvss.t831 935.633
R11095 dvss dvss.n2565 927.203
R11096 dvss.t1584 dvss.t648 920.795
R11097 dvss.t819 dvss.t1584 920.795
R11098 dvss.t819 dvss.t652 920.795
R11099 dvss.t652 dvss.t650 920.795
R11100 dvss.t1800 dvss 918.774
R11101 dvss.t1875 dvss 918.774
R11102 dvss.t1700 dvss 918.774
R11103 dvss.t620 dvss.t526 918.774
R11104 dvss dvss.t1706 918.774
R11105 dvss.t1272 dvss.t1056 918.774
R11106 dvss.t1787 dvss 918.774
R11107 dvss.t19 dvss.t519 918.774
R11108 dvss dvss.t1847 918.774
R11109 dvss.t1853 dvss 918.774
R11110 dvss.t1740 dvss 918.774
R11111 dvss dvss.t1714 918.774
R11112 dvss.t1703 dvss 918.774
R11113 dvss.t2036 dvss.t26 918.774
R11114 dvss.t1812 dvss 918.774
R11115 dvss.t715 dvss.t449 910.346
R11116 dvss.t1093 dvss.t469 910.346
R11117 dvss.t866 dvss.t2144 910.346
R11118 dvss dvss.n3759 901.917
R11119 dvss.t931 dvss.t1331 893.487
R11120 dvss.t1179 dvss 885.058
R11121 dvss.t1262 dvss.t1249 885.058
R11122 dvss.t717 dvss.t2232 885.058
R11123 dvss dvss.t2094 885.058
R11124 dvss.n2566 dvss.t440 876.629
R11125 dvss.t438 dvss.n3124 876.629
R11126 dvss.t720 dvss.t1805 868.199
R11127 dvss.n1755 dvss.t1029 867.946
R11128 dvss.n1730 dvss.t396 867.946
R11129 dvss dvss.t38 859.77
R11130 dvss.n4797 dvss 851.341
R11131 dvss.n4796 dvss 851.341
R11132 dvss.n4795 dvss 851.341
R11133 dvss.t84 dvss 851.341
R11134 dvss.n4794 dvss 851.341
R11135 dvss.t868 dvss.t1468 851.341
R11136 dvss.n4793 dvss 851.341
R11137 dvss.n4792 dvss 851.341
R11138 dvss.n4790 dvss 851.341
R11139 dvss.n4791 dvss 851.341
R11140 dvss dvss.n435 847.126
R11141 dvss.t2187 dvss.t1243 842.913
R11142 dvss.t379 dvss.t87 842.913
R11143 dvss.t925 dvss.t881 834.484
R11144 dvss.t1056 dvss.t1273 834.484
R11145 dvss.t917 dvss.t19 834.484
R11146 dvss.t1134 dvss.t2209 834.484
R11147 dvss.t269 dvss.t2036 834.484
R11148 dvss.n7045 dvss.n7044 833.506
R11149 dvss.n7045 dvss.n7001 833.506
R11150 dvss.n7044 dvss.n7015 833.13
R11151 dvss.n7015 dvss.n7001 833.13
R11152 dvss.t1956 dvss.t445 826.054
R11153 dvss.t27 dvss.t1781 826.054
R11154 dvss.t62 dvss.t68 819.513
R11155 dvss.t68 dvss.t64 819.513
R11156 dvss.t64 dvss.t76 819.513
R11157 dvss.t76 dvss.t70 819.513
R11158 dvss.t70 dvss.t66 819.513
R11159 dvss.t66 dvss.t78 819.513
R11160 dvss.t78 dvss.t72 819.513
R11161 dvss.t72 dvss.t54 819.513
R11162 dvss.t54 dvss.t50 819.513
R11163 dvss.t50 dvss.t56 819.513
R11164 dvss.t48 dvss.t74 819.513
R11165 dvss.t74 dvss.t58 819.513
R11166 dvss.t58 dvss.t52 819.513
R11167 dvss.t52 dvss.t60 819.513
R11168 dvss.t1181 dvss.t1187 819.513
R11169 dvss.t1187 dvss.t1185 819.513
R11170 dvss.t1185 dvss.t1183 819.513
R11171 dvss.t794 dvss.t854 817.625
R11172 dvss.t857 dvss.t790 817.625
R11173 dvss.t1399 dvss.t1572 809.196
R11174 dvss.t448 dvss.t1568 809.196
R11175 dvss.t721 dvss.t447 809.196
R11176 dvss.t991 dvss.t1016 809.196
R11177 dvss.t885 dvss.t726 809.196
R11178 dvss.t1574 dvss.t451 809.196
R11179 dvss.t1265 dvss.t1576 809.196
R11180 dvss.t1576 dvss.t637 809.196
R11181 dvss.t1267 dvss.t1221 809.196
R11182 dvss.t1222 dvss.t1208 809.196
R11183 dvss.t831 dvss.t1272 809.196
R11184 dvss.t1055 dvss.t1271 809.196
R11185 dvss.t100 dvss.t927 809.196
R11186 dvss.t519 dvss.t285 809.196
R11187 dvss.t522 dvss.t18 809.196
R11188 dvss.t2008 dvss.t2093 809.196
R11189 dvss.t458 dvss.t1094 809.196
R11190 dvss.t1173 dvss.t458 809.196
R11191 dvss.t1237 dvss.t692 809.196
R11192 dvss.t1972 dvss.t695 809.196
R11193 dvss.t1507 dvss.t1259 809.196
R11194 dvss.t1420 dvss.t24 809.196
R11195 dvss.t26 dvss.t309 809.196
R11196 dvss.t29 dvss.t2037 809.196
R11197 dvss.t1280 dvss.t541 809.196
R11198 dvss.t1138 dvss.t1144 808.754
R11199 dvss.t1144 dvss.t1140 808.754
R11200 dvss.t1140 dvss.t1152 808.754
R11201 dvss.t1152 dvss.t1146 808.754
R11202 dvss.t1146 dvss.t1142 808.754
R11203 dvss.t1142 dvss.t1154 808.754
R11204 dvss.t1154 dvss.t1148 808.754
R11205 dvss.t1148 dvss.t1162 808.754
R11206 dvss.t1162 dvss.t1158 808.754
R11207 dvss.t1158 dvss.t1164 808.754
R11208 dvss.t1156 dvss.t1150 808.754
R11209 dvss.t1150 dvss.t1166 808.754
R11210 dvss.t1166 dvss.t1160 808.754
R11211 dvss.t1160 dvss.t1136 808.754
R11212 dvss.t811 dvss.t801 808.754
R11213 dvss.t801 dvss.t803 808.754
R11214 dvss.t803 dvss.t809 808.754
R11215 dvss.t447 dvss.t16 800.766
R11216 dvss.t1271 dvss.t896 800.766
R11217 dvss.t1087 dvss.t522 800.766
R11218 dvss.t459 dvss.t983 800.766
R11219 dvss.t1992 dvss.t472 800.766
R11220 dvss.t2090 dvss.t1502 800.766
R11221 dvss.t2044 dvss.t1189 800.766
R11222 dvss.t2101 dvss.t688 800.766
R11223 dvss.t1201 dvss.t836 800.766
R11224 dvss.t87 dvss.t2015 800.766
R11225 dvss.t898 dvss.t746 800.766
R11226 dvss.t799 dvss.t971 800.766
R11227 dvss.t771 dvss.t29 800.766
R11228 dvss.t2074 dvss.t1981 800.766
R11229 dvss.t622 dvss.t2078 800.766
R11230 dvss.t881 dvss.t641 792.337
R11231 dvss.t543 dvss.t1833 792.337
R11232 dvss.t1754 dvss.t1878 775.48
R11233 dvss.t299 dvss.t302 775.48
R11234 dvss.t24 dvss.t1197 775.48
R11235 dvss.t1726 dvss.t1844 775.48
R11236 dvss.t2226 dvss.t696 775.48
R11237 dvss.n3335 dvss.n3334 769.572
R11238 dvss.n5494 dvss.n5493 769.572
R11239 dvss.n6987 dvss.n6986 769.572
R11240 dvss.t412 dvss.t662 767.051
R11241 dvss.t992 dvss.t414 767.051
R11242 dvss.t525 dvss.t2152 767.051
R11243 dvss.t914 dvss.t958 767.051
R11244 dvss.t408 dvss.t621 767.051
R11245 dvss.t741 dvss.t420 767.051
R11246 dvss.t833 dvss.t416 767.051
R11247 dvss.t946 dvss.t117 767.051
R11248 dvss.t962 dvss.t383 767.051
R11249 dvss.n6949 dvss.t1233 761.905
R11250 dvss.t361 dvss.n487 761.905
R11251 dvss.n6208 dvss.t780 761.905
R11252 dvss.t6 dvss.n862 761.905
R11253 dvss.n2105 dvss.t1340 761.905
R11254 dvss.n1985 dvss.t973 761.905
R11255 dvss.t2214 dvss.n1530 761.905
R11256 dvss.n6647 dvss.t1130 761.905
R11257 dvss.n5610 dvss.t1293 761.905
R11258 dvss.t60 dvss 760.976
R11259 dvss.t1711 dvss.t1217 758.621
R11260 dvss.t1136 dvss 750.986
R11261 dvss.t35 dvss.t868 750.192
R11262 dvss.n6900 dvss.n65 747.437
R11263 dvss.n662 dvss.n608 747.437
R11264 dvss.n6159 dvss.n789 747.437
R11265 dvss.n1007 dvss.n1006 747.437
R11266 dvss.n2056 dvss.n1439 747.437
R11267 dvss.n1878 dvss.n1503 747.437
R11268 dvss.n201 dvss.n189 747.437
R11269 dvss.n1059 dvss.n972 747.437
R11270 dvss.t396 dvss.t400 745.433
R11271 dvss.t2153 dvss.t1323 741.763
R11272 dvss.t1331 dvss.t601 741.763
R11273 dvss.t102 dvss.t379 741.763
R11274 dvss.t724 dvss.t735 741.763
R11275 dvss.t1416 dvss.t634 741.763
R11276 dvss.t177 dvss.t1215 741.763
R11277 dvss.t879 dvss.t1007 733.333
R11278 dvss.t993 dvss.t620 733.333
R11279 dvss dvss.t2006 733.333
R11280 dvss.t1183 dvss 731.707
R11281 dvss.t647 dvss.t1404 724.904
R11282 dvss.t996 dvss.t2208 724.904
R11283 dvss.t773 dvss.t1053 724.904
R11284 dvss.t575 dvss.t585 724.904
R11285 dvss.t585 dvss.t571 724.904
R11286 dvss.t591 dvss.t573 724.904
R11287 dvss.t2128 dvss.t2132 724.904
R11288 dvss.t1963 dvss.t1039 724.904
R11289 dvss.t2027 dvss.t2048 724.904
R11290 dvss.t1193 dvss.t2027 724.904
R11291 dvss.t144 dvss.t158 724.904
R11292 dvss.t164 dvss.t150 724.904
R11293 dvss.t162 dvss.t138 724.904
R11294 dvss.t156 dvss.t136 724.904
R11295 dvss.t890 dvss.t886 724.904
R11296 dvss.t733 dvss.t2146 724.904
R11297 dvss.t1243 dvss.t1239 724.904
R11298 dvss.t304 dvss.t1968 724.904
R11299 dvss.t1915 dvss.t475 724.904
R11300 dvss.t1850 dvss.t1285 724.904
R11301 dvss.t2126 dvss.t2136 724.904
R11302 dvss.t189 dvss.t2126 724.904
R11303 dvss.t181 dvss.t203 724.904
R11304 dvss.t179 dvss.t199 724.904
R11305 dvss.t185 dvss.t205 724.904
R11306 dvss.t193 dvss.t183 724.904
R11307 dvss.t809 dvss 722.101
R11308 dvss dvss.t643 716.476
R11309 dvss.t840 dvss.t1998 716.476
R11310 dvss.t587 dvss.n2846 716.476
R11311 dvss.t1039 dvss.t842 716.476
R11312 dvss.t134 dvss.t152 716.476
R11313 dvss.t2146 dvss.t838 716.476
R11314 dvss.t1418 dvss.t1358 716.476
R11315 dvss.t1317 dvss.t1472 716.476
R11316 dvss.t197 dvss.t179 716.476
R11317 dvss.t1110 dvss.t1009 708.047
R11318 dvss.t2149 dvss.t2147 708.047
R11319 dvss.t445 dvss.t707 708.047
R11320 dvss.t1014 dvss.t1012 708.047
R11321 dvss.t555 dvss.t561 708.047
R11322 dvss.t527 dvss.t711 708.047
R11323 dvss.t639 dvss.t638 708.047
R11324 dvss.t602 dvss.t1334 708.047
R11325 dvss.t1169 dvss.t2181 708.047
R11326 dvss.t1959 dvss.t1044 708.047
R11327 dvss.t702 dvss.t520 708.047
R11328 dvss.t1978 dvss 708.047
R11329 dvss.t1530 dvss.t175 708.047
R11330 dvss.t302 dvss.t1531 708.047
R11331 dvss.t864 dvss.t2067 708.047
R11332 dvss.t2017 dvss.t91 708.047
R11333 dvss.t1096 dvss.t1549 708.047
R11334 dvss.t460 dvss.t1096 708.047
R11335 dvss.t315 dvss.t1511 708.047
R11336 dvss.t89 dvss.t932 708.047
R11337 dvss.t988 dvss.t300 708.047
R11338 dvss.t1259 dvss.t508 708.047
R11339 dvss.t1500 dvss.t1498 708.047
R11340 dvss.t796 dvss.t2123 708.047
R11341 dvss.t859 dvss.t796 708.047
R11342 dvss.t1448 dvss.t2115 708.047
R11343 dvss.t2115 dvss.t857 708.047
R11344 dvss.t4 dvss.t2 708.047
R11345 dvss.t1356 dvss.t1354 708.047
R11346 dvss.t2230 dvss.t2228 708.047
R11347 dvss.t500 dvss.t27 708.047
R11348 dvss.t372 dvss.t374 708.047
R11349 dvss.t1048 dvss.t372 708.047
R11350 dvss.t921 dvss.t1168 708.047
R11351 dvss.t2078 dvss.t2076 708.047
R11352 dvss.t2134 dvss.t549 699.617
R11353 dvss.t875 dvss.t1112 699.617
R11354 dvss.t154 dvss.t442 699.617
R11355 dvss.t1393 dvss.t164 699.617
R11356 dvss.t1582 dvss 699.617
R11357 dvss.t32 dvss.t834 699.617
R11358 dvss.t1931 dvss.t583 691.188
R11359 dvss.t1398 dvss.t1526 691.188
R11360 dvss dvss.t1394 691.188
R11361 dvss.t187 dvss 691.188
R11362 dvss dvss.t1448 691.188
R11363 dvss.t309 dvss.t1921 691.188
R11364 dvss.t170 dvss 682.76
R11365 dvss.t1454 dvss.t1390 682.76
R11366 dvss.t211 dvss 682.76
R11367 dvss.t848 dvss.t2113 682.76
R11368 dvss.n436 dvss.t245 682.76
R11369 dvss.t641 dvss.t1760 674.331
R11370 dvss.t2208 dvss.t750 674.331
R11371 dvss.t1170 dvss.t626 674.331
R11372 dvss.t465 dvss.t1237 674.331
R11373 dvss.t1275 dvss.t990 674.331
R11374 dvss.t98 dvss.t381 674.331
R11375 dvss.t2013 dvss.t935 674.331
R11376 dvss.t2002 dvss.t1199 674.331
R11377 dvss.t569 dvss 665.9
R11378 dvss.t844 dvss.t1219 657.471
R11379 dvss.t317 dvss.t2177 657.471
R11380 dvss.t1135 dvss.t693 657.471
R11381 dvss.t213 dvss.t1351 657.471
R11382 dvss.t1304 dvss.t1971 649.043
R11383 dvss.t932 dvss.t2191 649.043
R11384 dvss.n2565 dvss 640.614
R11385 dvss.t452 dvss.t1397 640.614
R11386 dvss.t1470 dvss.t140 640.614
R11387 dvss.t384 dvss.t2083 640.614
R11388 dvss.t1276 dvss.t173 640.614
R11389 dvss.t2155 dvss.t1283 640.614
R11390 dvss.t498 dvss.t2169 640.614
R11391 dvss.n4806 dvss.n2305 640.361
R11392 dvss.n4806 dvss.n4805 637.461
R11393 dvss.t1720 dvss 632.184
R11394 dvss.n2448 dvss 632.184
R11395 dvss.t1729 dvss 632.184
R11396 dvss.n2988 dvss 632.184
R11397 dvss.t1797 dvss 632.184
R11398 dvss.n3338 dvss 632.184
R11399 dvss.t1863 dvss 632.184
R11400 dvss.t1872 dvss 632.184
R11401 dvss.n3527 dvss 632.184
R11402 dvss.t2065 dvss.t690 632.184
R11403 dvss.t2186 dvss.t1245 632.184
R11404 dvss.n3908 dvss 632.184
R11405 dvss.t1688 dvss 632.184
R11406 dvss dvss.t1723 632.184
R11407 dvss dvss.n4789 632.184
R11408 dvss.n4545 dvss 632.184
R11409 dvss.n4593 dvss 632.184
R11410 dvss dvss.t1825 632.184
R11411 dvss dvss.n4491 632.184
R11412 dvss.n4316 dvss 632.184
R11413 dvss.t93 dvss.t166 623.755
R11414 dvss.t583 dvss 615.327
R11415 dvss.n3759 dvss 615.327
R11416 dvss.t160 dvss.t1977 615.327
R11417 dvss.t892 dvss.t1174 615.327
R11418 dvss dvss.t370 615.327
R11419 dvss.t1257 dvss.n1572 610.777
R11420 dvss.n3337 dvss.n3126 608.452
R11421 dvss.n6359 dvss.n6358 607.51
R11422 dvss.n6408 dvss.n6401 607.51
R11423 dvss.t640 dvss.t870 606.898
R11424 dvss.t1402 dvss.t640 606.898
R11425 dvss.t748 dvss.t563 606.898
R11426 dvss.t750 dvss.t424 606.898
R11427 dvss.t713 dvss.t941 606.898
R11428 dvss.t453 dvss.t642 606.898
R11429 dvss.t1525 dvss.t2175 606.898
R11430 dvss.t636 dvss.t456 606.898
R11431 dvss.t356 dvss.t406 606.898
R11432 dvss.t430 dvss.t148 606.898
R11433 dvss.t418 dvss.t1582 606.898
R11434 dvss.t1330 dvss.t597 606.898
R11435 dvss.t386 dvss.t1994 606.898
R11436 dvss.t956 dvss.t1965 606.898
R11437 dvss.t2113 dvss.t2069 606.898
R11438 dvss.t852 dvss.t1910 606.898
R11439 dvss.t104 dvss.t798 606.898
R11440 dvss.n236 dvss.t1517 604.145
R11441 dvss.n2565 dvss.n2564 599.125
R11442 dvss.n4193 dvss.t432 598.467
R11443 dvss.n3300 dvss.n3159 593.402
R11444 dvss.n6357 dvss.n235 592.001
R11445 dvss.n6517 dvss.n6516 592.001
R11446 dvss.n6816 dvss.n6815 590.068
R11447 dvss.n6742 dvss.n6741 590.068
R11448 dvss.n5928 dvss.n5927 590.068
R11449 dvss.n6001 dvss.n6000 590.068
R11450 dvss.n5848 dvss.n5847 590.068
R11451 dvss.n5767 dvss.n5766 590.068
R11452 dvss.n2010 dvss.n2009 590.068
R11453 dvss.n1641 dvss.n1640 590.068
R11454 dvss.n1667 dvss.n1666 590.068
R11455 dvss.t589 dvss.t704 590.038
R11456 dvss.t2181 dvss 590.038
R11457 dvss.t1044 dvss.t1338 590.038
R11458 dvss.n3760 dvss.t1471 590.038
R11459 dvss.t1431 dvss.t477 590.038
R11460 dvss.t1983 dvss.t1509 590.038
R11461 dvss.t1350 dvss.t390 590.038
R11462 dvss.n3126 dvss.n3125 588.648
R11463 dvss.n6518 dvss.n6400 588.516
R11464 dvss.n3303 dvss.n3302 587.614
R11465 dvss.n6819 dvss.n6818 587.271
R11466 dvss.n6755 dvss.n102 587.271
R11467 dvss.n5931 dvss.n5918 587.271
R11468 dvss.n6004 dvss.n5976 587.271
R11469 dvss.n5861 dvss.n831 587.271
R11470 dvss.n5768 dvss.n863 587.271
R11471 dvss.n2008 dvss.n2007 587.271
R11472 dvss.n1637 dvss.n1636 587.271
R11473 dvss.n1665 dvss.n1633 587.271
R11474 dvss.n3301 dvss.n3154 586.313
R11475 dvss.n5602 dvss.n1131 585.389
R11476 dvss.n5604 dvss.n5603 585.197
R11477 dvss.n504 dvss.n503 585
R11478 dvss.n503 dvss.n502 585
R11479 dvss.n6249 dvss.n6248 585
R11480 dvss.n6250 dvss.n6249 585
R11481 dvss.n501 dvss.n500 585
R11482 dvss.n6251 dvss.n501 585
R11483 dvss.n6255 dvss.n6254 585
R11484 dvss.n6254 dvss.n6253 585
R11485 dvss.n498 dvss.n497 585
R11486 dvss.n6252 dvss.n497 585
R11487 dvss.n6265 dvss.n6264 585
R11488 dvss.n6266 dvss.n6265 585
R11489 dvss.n496 dvss.n495 585
R11490 dvss.n6267 dvss.n496 585
R11491 dvss.n6270 dvss.n6269 585
R11492 dvss.n6269 dvss.n6268 585
R11493 dvss.n494 dvss.n493 585
R11494 dvss.n493 dvss.n492 585
R11495 dvss.n6276 dvss.n6275 585
R11496 dvss.n6277 dvss.n6276 585
R11497 dvss.n491 dvss.n490 585
R11498 dvss.n6278 dvss.n491 585
R11499 dvss.n6282 dvss.n6281 585
R11500 dvss.n6281 dvss.n6280 585
R11501 dvss.n489 dvss.n488 585
R11502 dvss.n6279 dvss.n488 585
R11503 dvss.n6290 dvss.n6289 585
R11504 dvss.n6291 dvss.n6290 585
R11505 dvss.n486 dvss.n485 585
R11506 dvss.n6292 dvss.n486 585
R11507 dvss.n6295 dvss.n6294 585
R11508 dvss.n6294 dvss.n6293 585
R11509 dvss.n479 dvss.n478 585
R11510 dvss.n478 dvss.n477 585
R11511 dvss.n6307 dvss.n6306 585
R11512 dvss.n6308 dvss.n6307 585
R11513 dvss.n480 dvss.n476 585
R11514 dvss.n6309 dvss.n476 585
R11515 dvss.n6311 dvss.n475 585
R11516 dvss.n6311 dvss.n6310 585
R11517 dvss.n6317 dvss.n6316 585
R11518 dvss.n6316 dvss.n6315 585
R11519 dvss.n6312 dvss.n472 585
R11520 dvss.n6314 dvss.n6312 585
R11521 dvss.n6321 dvss.n473 585
R11522 dvss.n6313 dvss.n473 585
R11523 dvss.n6322 dvss.n470 585
R11524 dvss.n470 dvss.n469 585
R11525 dvss.n6333 dvss.n6332 585
R11526 dvss.n6334 dvss.n6333 585
R11527 dvss.n471 dvss.n467 585
R11528 dvss.n6335 dvss.n467 585
R11529 dvss.n6337 dvss.n468 585
R11530 dvss.n6337 dvss.n6336 585
R11531 dvss.n6338 dvss.n459 585
R11532 dvss.n6339 dvss.n6338 585
R11533 dvss.n6577 dvss.n460 585
R11534 dvss.n6340 dvss.n460 585
R11535 dvss.n6576 dvss.n461 585
R11536 dvss.n6341 dvss.n461 585
R11537 dvss.n6342 dvss.n462 585
R11538 dvss.n6343 dvss.n6342 585
R11539 dvss.n6572 dvss.n463 585
R11540 dvss.n6344 dvss.n463 585
R11541 dvss.n5573 dvss.n5572 585
R11542 dvss.n5572 dvss.n5571 585
R11543 dvss.n523 dvss.n522 585
R11544 dvss.n524 dvss.n523 585
R11545 dvss.n6211 dvss.n6210 585
R11546 dvss.n6210 dvss.n6209 585
R11547 dvss.n521 dvss.n520 585
R11548 dvss.n525 dvss.n520 585
R11549 dvss.n6219 dvss.n6218 585
R11550 dvss.n6220 dvss.n6219 585
R11551 dvss.n518 dvss.n514 585
R11552 dvss.n6221 dvss.n518 585
R11553 dvss.n6226 dvss.n6225 585
R11554 dvss.n6225 dvss.n6224 585
R11555 dvss.n519 dvss.n517 585
R11556 dvss.n6223 dvss.n519 585
R11557 dvss.n509 dvss.n508 585
R11558 dvss.n6222 dvss.n508 585
R11559 dvss.n6237 dvss.n6236 585
R11560 dvss.n6238 dvss.n6237 585
R11561 dvss.n506 dvss.n505 585
R11562 dvss.n6240 dvss.n506 585
R11563 dvss.n6243 dvss.n6242 585
R11564 dvss.n6242 dvss.n6241 585
R11565 dvss.n1569 dvss.n1567 585
R11566 dvss.n1593 dvss.n1569 585
R11567 dvss.n1582 dvss.n1581 585
R11568 dvss.n1580 dvss.n1579 585
R11569 dvss.n1590 dvss.n1589 585
R11570 dvss.n1591 dvss.n1554 585
R11571 dvss.n1552 dvss.n1551 585
R11572 dvss.n1577 dvss.n1551 585
R11573 dvss.n1791 dvss.n1790 585
R11574 dvss.n1792 dvss.n1791 585
R11575 dvss.n1548 dvss.n1547 585
R11576 dvss.n1795 dvss.n1548 585
R11577 dvss.n1799 dvss.n1798 585
R11578 dvss.n1798 dvss.n1797 585
R11579 dvss.n1542 dvss.n1541 585
R11580 dvss.n1796 dvss.n1541 585
R11581 dvss.n1813 dvss.n1812 585
R11582 dvss.n1814 dvss.n1813 585
R11583 dvss.n1537 dvss.n1536 585
R11584 dvss.n1817 dvss.n1537 585
R11585 dvss.n1822 dvss.n1821 585
R11586 dvss.n1821 dvss.n1820 585
R11587 dvss.n1532 dvss.n1531 585
R11588 dvss.n1538 dvss.n1531 585
R11589 dvss.n1833 dvss.n1832 585
R11590 dvss.n1834 dvss.n1833 585
R11591 dvss.n1527 dvss.n1526 585
R11592 dvss.n1526 dvss.n1524 585
R11593 dvss.n1847 dvss.n1846 585
R11594 dvss.n1848 dvss.n1847 585
R11595 dvss.n1522 dvss.n1516 585
R11596 dvss.n1849 dvss.n1522 585
R11597 dvss.n1855 dvss.n1854 585
R11598 dvss.n1854 dvss.n1853 585
R11599 dvss.n1523 dvss.n1510 585
R11600 dvss.n1852 dvss.n1523 585
R11601 dvss.n1867 dvss.n1511 585
R11602 dvss.n1851 dvss.n1511 585
R11603 dvss.n1868 dvss.n1504 585
R11604 dvss.n1873 dvss.n1504 585
R11605 dvss.n1875 dvss.n1505 585
R11606 dvss.n1875 dvss.n1874 585
R11607 dvss.n1876 dvss.n1496 585
R11608 dvss.n1498 dvss.n1497 585
R11609 dvss.n1881 dvss.n1880 585
R11610 dvss.n1499 dvss.n1488 585
R11611 dvss.n1501 dvss.n1500 585
R11612 dvss.n1502 dvss.n1501 585
R11613 dvss.n1484 dvss.n1483 585
R11614 dvss.n1901 dvss.n1484 585
R11615 dvss.n1904 dvss.n1903 585
R11616 dvss.n1903 dvss.n1902 585
R11617 dvss.n1480 dvss.n1479 585
R11618 dvss.n1914 dvss.n1480 585
R11619 dvss.n1917 dvss.n1916 585
R11620 dvss.n1916 dvss.n1915 585
R11621 dvss.n1476 dvss.n1472 585
R11622 dvss.n1929 dvss.n1472 585
R11623 dvss.n1932 dvss.n1473 585
R11624 dvss.n1932 dvss.n1931 585
R11625 dvss.n1933 dvss.n1466 585
R11626 dvss.n1934 dvss.n1933 585
R11627 dvss.n1460 dvss.n1458 585
R11628 dvss.n1469 dvss.n1458 585
R11629 dvss.n1983 dvss.n1982 585
R11630 dvss.n1984 dvss.n1983 585
R11631 dvss.n1461 dvss.n1459 585
R11632 dvss.n1954 dvss.n1459 585
R11633 dvss.n1952 dvss.n1945 585
R11634 dvss.n1955 dvss.n1952 585
R11635 dvss.n1959 dvss.n1953 585
R11636 dvss.n1959 dvss.n1958 585
R11637 dvss.n1960 dvss.n1949 585
R11638 dvss.n1961 dvss.n1960 585
R11639 dvss.n1455 dvss.n1454 585
R11640 dvss.n1962 dvss.n1455 585
R11641 dvss.n2020 dvss.n2019 585
R11642 dvss.n2019 dvss.n2018 585
R11643 dvss.n1444 dvss.n1442 585
R11644 dvss.n1442 dvss.n1440 585
R11645 dvss.n2054 dvss.n2053 585
R11646 dvss.n2055 dvss.n2054 585
R11647 dvss.n1445 dvss.n1443 585
R11648 dvss.n2031 dvss.n2029 585
R11649 dvss.n2035 dvss.n2034 585
R11650 dvss.n2032 dvss.n1433 585
R11651 dvss.n2062 dvss.n1434 585
R11652 dvss.n2058 dvss.n1434 585
R11653 dvss.n2063 dvss.n1430 585
R11654 dvss.n2057 dvss.n1430 585
R11655 dvss.n2070 dvss.n1429 585
R11656 dvss.n2070 dvss.n2069 585
R11657 dvss.n2072 dvss.n2071 585
R11658 dvss.n2071 dvss.n1422 585
R11659 dvss.n1425 dvss.n1420 585
R11660 dvss.n2082 dvss.n1420 585
R11661 dvss.n2084 dvss.n1421 585
R11662 dvss.n2084 dvss.n2083 585
R11663 dvss.n2085 dvss.n1412 585
R11664 dvss.n2086 dvss.n2085 585
R11665 dvss.n1353 dvss.n1351 585
R11666 dvss.n1417 dvss.n1351 585
R11667 dvss.n2103 dvss.n2102 585
R11668 dvss.n2104 dvss.n2103 585
R11669 dvss.n1354 dvss.n1352 585
R11670 dvss.n1352 dvss.n1349 585
R11671 dvss.n1378 dvss.n1377 585
R11672 dvss.n1380 dvss.n1378 585
R11673 dvss.n1383 dvss.n1382 585
R11674 dvss.n1382 dvss.n1381 585
R11675 dvss.n1370 dvss.n1365 585
R11676 dvss.n1392 dvss.n1365 585
R11677 dvss.n1394 dvss.n1366 585
R11678 dvss.n1394 dvss.n1393 585
R11679 dvss.n1395 dvss.n1361 585
R11680 dvss.n1396 dvss.n1395 585
R11681 dvss.n893 dvss.n891 585
R11682 dvss.n891 dvss.n888 585
R11683 dvss.n5729 dvss.n5728 585
R11684 dvss.n5730 dvss.n5729 585
R11685 dvss.n894 dvss.n892 585
R11686 dvss.n892 dvss.n890 585
R11687 dvss.n1004 dvss.n899 585
R11688 dvss.n1003 dvss.n900 585
R11689 dvss.n1002 dvss.n904 585
R11690 dvss.n1000 dvss.n905 585
R11691 dvss.n999 dvss.n998 585
R11692 dvss.n1015 dvss.n999 585
R11693 dvss.n1017 dvss.n909 585
R11694 dvss.n1017 dvss.n1016 585
R11695 dvss.n1018 dvss.n914 585
R11696 dvss.n1019 dvss.n1018 585
R11697 dvss.n994 dvss.n993 585
R11698 dvss.n1020 dvss.n993 585
R11699 dvss.n1024 dvss.n997 585
R11700 dvss.n1024 dvss.n1023 585
R11701 dvss.n1026 dvss.n920 585
R11702 dvss.n1027 dvss.n1026 585
R11703 dvss.n1025 dvss.n925 585
R11704 dvss.n1025 dvss.n992 585
R11705 dvss.n990 dvss.n926 585
R11706 dvss.n1030 dvss.n990 585
R11707 dvss.n1034 dvss.n991 585
R11708 dvss.n1034 dvss.n1033 585
R11709 dvss.n1036 dvss.n929 585
R11710 dvss.n1036 dvss.n1035 585
R11711 dvss.n1037 dvss.n934 585
R11712 dvss.n1037 dvss.n989 585
R11713 dvss.n1038 dvss.n935 585
R11714 dvss.n1039 dvss.n1038 585
R11715 dvss.n979 dvss.n978 585
R11716 dvss.n1040 dvss.n978 585
R11717 dvss.n1046 dvss.n1045 585
R11718 dvss.n1047 dvss.n1046 585
R11719 dvss.n980 dvss.n974 585
R11720 dvss.n1048 dvss.n974 585
R11721 dvss.n1052 dvss.n975 585
R11722 dvss.n1052 dvss.n1051 585
R11723 dvss.n1053 dvss.n944 585
R11724 dvss.n1054 dvss.n1053 585
R11725 dvss.n1056 dvss.n949 585
R11726 dvss.n1056 dvss.n1055 585
R11727 dvss.n5649 dvss.n1075 585
R11728 dvss.n1119 dvss.n1075 585
R11729 dvss.n1113 dvss.n1076 585
R11730 dvss.n1121 dvss.n1113 585
R11731 dvss.n5613 dvss.n1115 585
R11732 dvss.n5613 dvss.n5612 585
R11733 dvss.n5614 dvss.n1101 585
R11734 dvss.n5615 dvss.n5614 585
R11735 dvss.n1111 dvss.n1105 585
R11736 dvss.n5616 dvss.n1111 585
R11737 dvss.n5619 dvss.n1112 585
R11738 dvss.n5619 dvss.n5618 585
R11739 dvss.n5620 dvss.n1109 585
R11740 dvss.n5621 dvss.n5620 585
R11741 dvss.n805 dvss.n804 585
R11742 dvss.n5622 dvss.n805 585
R11743 dvss.n6123 dvss.n6122 585
R11744 dvss.n6122 dvss.n6121 585
R11745 dvss.n794 dvss.n792 585
R11746 dvss.n792 dvss.n790 585
R11747 dvss.n6157 dvss.n6156 585
R11748 dvss.n6158 dvss.n6157 585
R11749 dvss.n795 dvss.n793 585
R11750 dvss.n6134 dvss.n6132 585
R11751 dvss.n6138 dvss.n6137 585
R11752 dvss.n6135 dvss.n783 585
R11753 dvss.n6165 dvss.n784 585
R11754 dvss.n6161 dvss.n784 585
R11755 dvss.n6166 dvss.n780 585
R11756 dvss.n6160 dvss.n780 585
R11757 dvss.n6173 dvss.n779 585
R11758 dvss.n6173 dvss.n6172 585
R11759 dvss.n6175 dvss.n6174 585
R11760 dvss.n6174 dvss.n772 585
R11761 dvss.n775 dvss.n770 585
R11762 dvss.n6185 dvss.n770 585
R11763 dvss.n6187 dvss.n771 585
R11764 dvss.n6187 dvss.n6186 585
R11765 dvss.n6188 dvss.n762 585
R11766 dvss.n6189 dvss.n6188 585
R11767 dvss.n530 dvss.n528 585
R11768 dvss.n767 dvss.n528 585
R11769 dvss.n6206 dvss.n6205 585
R11770 dvss.n6207 dvss.n6206 585
R11771 dvss.n531 dvss.n529 585
R11772 dvss.n529 dvss.n526 585
R11773 dvss.n628 dvss.n627 585
R11774 dvss.n629 dvss.n628 585
R11775 dvss.n635 dvss.n634 585
R11776 dvss.n634 dvss.n633 585
R11777 dvss.n615 dvss.n614 585
R11778 dvss.n632 dvss.n614 585
R11779 dvss.n646 dvss.n645 585
R11780 dvss.n647 dvss.n646 585
R11781 dvss.n616 dvss.n610 585
R11782 dvss.n648 dvss.n610 585
R11783 dvss.n652 dvss.n611 585
R11784 dvss.n652 dvss.n651 585
R11785 dvss.n653 dvss.n539 585
R11786 dvss.n653 dvss.n609 585
R11787 dvss.n660 dvss.n544 585
R11788 dvss.n661 dvss.n660 585
R11789 dvss.n659 dvss.n545 585
R11790 dvss.n657 dvss.n546 585
R11791 dvss.n656 dvss.n550 585
R11792 dvss.n654 dvss.n551 585
R11793 dvss.n607 dvss.n606 585
R11794 dvss.n670 dvss.n607 585
R11795 dvss.n672 dvss.n555 585
R11796 dvss.n672 dvss.n671 585
R11797 dvss.n673 dvss.n560 585
R11798 dvss.n674 dvss.n673 585
R11799 dvss.n602 dvss.n601 585
R11800 dvss.n675 dvss.n601 585
R11801 dvss.n679 dvss.n605 585
R11802 dvss.n679 dvss.n678 585
R11803 dvss.n681 dvss.n566 585
R11804 dvss.n682 dvss.n681 585
R11805 dvss.n680 dvss.n571 585
R11806 dvss.n680 dvss.n600 585
R11807 dvss.n598 dvss.n572 585
R11808 dvss.n685 dvss.n598 585
R11809 dvss.n689 dvss.n599 585
R11810 dvss.n689 dvss.n688 585
R11811 dvss.n691 dvss.n575 585
R11812 dvss.n691 dvss.n690 585
R11813 dvss.n692 dvss.n580 585
R11814 dvss.n692 dvss.n597 585
R11815 dvss.n693 dvss.n581 585
R11816 dvss.n694 dvss.n693 585
R11817 dvss.n594 dvss.n593 585
R11818 dvss.n698 dvss.n593 585
R11819 dvss.n700 dvss.n596 585
R11820 dvss.n700 dvss.n699 585
R11821 dvss.n701 dvss.n589 585
R11822 dvss.n702 dvss.n701 585
R11823 dvss.n127 dvss.n125 585
R11824 dvss.n125 dvss.n122 585
R11825 dvss.n6713 dvss.n6712 585
R11826 dvss.n6714 dvss.n6713 585
R11827 dvss.n128 dvss.n126 585
R11828 dvss.n126 dvss.n124 585
R11829 dvss.n221 dvss.n160 585
R11830 dvss.n222 dvss.n221 585
R11831 dvss.n182 dvss.n181 585
R11832 dvss.n225 dvss.n182 585
R11833 dvss.n6649 dvss.n163 585
R11834 dvss.n6649 dvss.n6648 585
R11835 dvss.n6650 dvss.n171 585
R11836 dvss.n6651 dvss.n6650 585
R11837 dvss.n179 dvss.n172 585
R11838 dvss.n6652 dvss.n179 585
R11839 dvss.n6656 dvss.n180 585
R11840 dvss.n6656 dvss.n6655 585
R11841 dvss.n6657 dvss.n176 585
R11842 dvss.n6658 dvss.n6657 585
R11843 dvss.n76 dvss.n75 585
R11844 dvss.n6659 dvss.n76 585
R11845 dvss.n6864 dvss.n6863 585
R11846 dvss.n6863 dvss.n6862 585
R11847 dvss.n70 dvss.n68 585
R11848 dvss.n68 dvss.n66 585
R11849 dvss.n6898 dvss.n6897 585
R11850 dvss.n6899 dvss.n6898 585
R11851 dvss.n71 dvss.n69 585
R11852 dvss.n6875 dvss.n6873 585
R11853 dvss.n6879 dvss.n6878 585
R11854 dvss.n6876 dvss.n59 585
R11855 dvss.n6906 dvss.n60 585
R11856 dvss.n6902 dvss.n60 585
R11857 dvss.n6907 dvss.n56 585
R11858 dvss.n6901 dvss.n56 585
R11859 dvss.n6914 dvss.n55 585
R11860 dvss.n6914 dvss.n6913 585
R11861 dvss.n6916 dvss.n6915 585
R11862 dvss.n6915 dvss.n48 585
R11863 dvss.n51 dvss.n46 585
R11864 dvss.n6926 dvss.n46 585
R11865 dvss.n6928 dvss.n47 585
R11866 dvss.n6928 dvss.n6927 585
R11867 dvss.n6929 dvss.n38 585
R11868 dvss.n6930 dvss.n6929 585
R11869 dvss.n28 dvss.n26 585
R11870 dvss.n43 dvss.n26 585
R11871 dvss.n6947 dvss.n6946 585
R11872 dvss.n6948 dvss.n6947 585
R11873 dvss.n29 dvss.n27 585
R11874 dvss.n27 dvss.n24 585
R11875 dvss.n6458 dvss.n6457 585
R11876 dvss.n6459 dvss.n6458 585
R11877 dvss.n6447 dvss.n6446 585
R11878 dvss.n6460 dvss.n6446 585
R11879 dvss.n6470 dvss.n6469 585
R11880 dvss.n6471 dvss.n6470 585
R11881 dvss.n6443 dvss.n6442 585
R11882 dvss.n6472 dvss.n6442 585
R11883 dvss.n6478 dvss.n6477 585
R11884 dvss.n6479 dvss.n6478 585
R11885 dvss.n6439 dvss.n6438 585
R11886 dvss.n6480 dvss.n6438 585
R11887 dvss.n6489 dvss.n6488 585
R11888 dvss.n6489 dvss.n6437 585
R11889 dvss.n6490 dvss.n6433 585
R11890 dvss.n6491 dvss.n6490 585
R11891 dvss.n6496 dvss.n6434 585
R11892 dvss.n6434 dvss.n6429 585
R11893 dvss.n6497 dvss.n6430 585
R11894 dvss.n6501 dvss.n6430 585
R11895 dvss.n199 dvss.n133 585
R11896 dvss.n198 dvss.n134 585
R11897 dvss.n197 dvss.n138 585
R11898 dvss.n203 dvss.n139 585
R11899 dvss.n205 dvss.n204 585
R11900 dvss.n206 dvss.n205 585
R11901 dvss.n188 dvss.n143 585
R11902 dvss.n207 dvss.n188 585
R11903 dvss.n209 dvss.n148 585
R11904 dvss.n209 dvss.n208 585
R11905 dvss.n211 dvss.n210 585
R11906 dvss.n210 dvss.n185 585
R11907 dvss.n215 dvss.n214 585
R11908 dvss.n216 dvss.n215 585
R11909 dvss.n184 dvss.n154 585
R11910 dvss.n217 dvss.n184 585
R11911 dvss.n220 dvss.n159 585
R11912 dvss.n220 dvss.n219 585
R11913 dvss.n6571 dvss.n6570 585
R11914 dvss.n6570 dvss.n6569 585
R11915 dvss.n466 dvss.n465 585
R11916 dvss.n6568 dvss.n466 585
R11917 dvss.n6566 dvss.n6565 585
R11918 dvss.n6567 dvss.n6566 585
R11919 dvss.n230 dvss.n228 585
R11920 dvss.n228 dvss.n226 585
R11921 dvss.n6645 dvss.n6644 585
R11922 dvss.n6646 dvss.n6645 585
R11923 dvss.n6643 dvss.n229 585
R11924 dvss.n229 dvss.n227 585
R11925 dvss.n6642 dvss.n6641 585
R11926 dvss.n6641 dvss.n6640 585
R11927 dvss.n235 dvss.n234 585
R11928 dvss.n6359 dvss.n6356 585
R11929 dvss.n6360 dvss.n6350 585
R11930 dvss.n6362 dvss.n6360 585
R11931 dvss.n6554 dvss.n6553 585
R11932 dvss.n6553 dvss.n6552 585
R11933 dvss.n6361 dvss.n6351 585
R11934 dvss.n6551 dvss.n6361 585
R11935 dvss.n6549 dvss.n6548 585
R11936 dvss.n6550 dvss.n6549 585
R11937 dvss.n6547 dvss.n6364 585
R11938 dvss.n6364 dvss.n6363 585
R11939 dvss.n6546 dvss.n6545 585
R11940 dvss.n6545 dvss.n6544 585
R11941 dvss.n6370 dvss.n6369 585
R11942 dvss.n6543 dvss.n6370 585
R11943 dvss.n6541 dvss.n6540 585
R11944 dvss.n6542 dvss.n6541 585
R11945 dvss.n6539 dvss.n6371 585
R11946 dvss.n6383 dvss.n6371 585
R11947 dvss.n6538 dvss.n6537 585
R11948 dvss.n6537 dvss.n6536 585
R11949 dvss.n6382 dvss.n6381 585
R11950 dvss.n6535 dvss.n6382 585
R11951 dvss.n6533 dvss.n6532 585
R11952 dvss.n6534 dvss.n6533 585
R11953 dvss.n6531 dvss.n6385 585
R11954 dvss.n6385 dvss.n6384 585
R11955 dvss.n6530 dvss.n6529 585
R11956 dvss.n6529 dvss.n6528 585
R11957 dvss.n6391 dvss.n6390 585
R11958 dvss.n6527 dvss.n6391 585
R11959 dvss.n6525 dvss.n6524 585
R11960 dvss.n6526 dvss.n6525 585
R11961 dvss.n6523 dvss.n6393 585
R11962 dvss.n6393 dvss.n6392 585
R11963 dvss.n6522 dvss.n6521 585
R11964 dvss.n6521 dvss.n6520 585
R11965 dvss.n6399 dvss.n6398 585
R11966 dvss.n6519 dvss.n6399 585
R11967 dvss.n6402 dvss.n6400 585
R11968 dvss.n6516 dvss.n6515 585
R11969 dvss.n6514 dvss.n6401 585
R11970 dvss.n6513 dvss.n6512 585
R11971 dvss.n6512 dvss.n6511 585
R11972 dvss.n6407 dvss.n6406 585
R11973 dvss.n6510 dvss.n6407 585
R11974 dvss.n6508 dvss.n6507 585
R11975 dvss.n6509 dvss.n6508 585
R11976 dvss.n6506 dvss.n6410 585
R11977 dvss.n6410 dvss.n6409 585
R11978 dvss.n6505 dvss.n6504 585
R11979 dvss.n6504 dvss.n6503 585
R11980 dvss.n3169 dvss.n3168 585
R11981 dvss.n3239 dvss.n3168 585
R11982 dvss.n3251 dvss.n3250 585
R11983 dvss.n3252 dvss.n3251 585
R11984 dvss.n3167 dvss.n3166 585
R11985 dvss.n3253 dvss.n3167 585
R11986 dvss.n3256 dvss.n3255 585
R11987 dvss.n3255 dvss.n3254 585
R11988 dvss.n3164 dvss.n3162 585
R11989 dvss.n3162 dvss.n3160 585
R11990 dvss.n3263 dvss.n3262 585
R11991 dvss.n3264 dvss.n3263 585
R11992 dvss.n3165 dvss.n3163 585
R11993 dvss.n3163 dvss.n3161 585
R11994 dvss.n240 dvss.n239 585
R11995 dvss.n239 dvss.n238 585
R11996 dvss.n6636 dvss.n6635 585
R11997 dvss.n6637 dvss.n6636 585
R11998 dvss.n3199 dvss.n3198 585
R11999 dvss.n3198 dvss.n3197 585
R12000 dvss.n3195 dvss.n3194 585
R12001 dvss.n3194 dvss.n3193 585
R12002 dvss.n3205 dvss.n3204 585
R12003 dvss.n3206 dvss.n3205 585
R12004 dvss.n3192 dvss.n3191 585
R12005 dvss.n3207 dvss.n3192 585
R12006 dvss.n3210 dvss.n3209 585
R12007 dvss.n3209 dvss.n3208 585
R12008 dvss.n3187 dvss.n3186 585
R12009 dvss.n3186 dvss.n3185 585
R12010 dvss.n3220 dvss.n3219 585
R12011 dvss.n3221 dvss.n3220 585
R12012 dvss.n3184 dvss.n3183 585
R12013 dvss.n3222 dvss.n3184 585
R12014 dvss.n3226 dvss.n3225 585
R12015 dvss.n3225 dvss.n3224 585
R12016 dvss.n3177 dvss.n3176 585
R12017 dvss.n3223 dvss.n3176 585
R12018 dvss.n3235 dvss.n3234 585
R12019 dvss.n3236 dvss.n3235 585
R12020 dvss.n3175 dvss.n3174 585
R12021 dvss.n3238 dvss.n3175 585
R12022 dvss.n3242 dvss.n3241 585
R12023 dvss.n3241 dvss.n3240 585
R12024 dvss.n3134 dvss.n3132 585
R12025 dvss.n3136 dvss.n3134 585
R12026 dvss.n3328 dvss.n3327 585
R12027 dvss.n3327 dvss.n3326 585
R12028 dvss.n3135 dvss.n3133 585
R12029 dvss.n3325 dvss.n3135 585
R12030 dvss.n3323 dvss.n3322 585
R12031 dvss.n3324 dvss.n3323 585
R12032 dvss.n3321 dvss.n3138 585
R12033 dvss.n3138 dvss.n3137 585
R12034 dvss.n3320 dvss.n3319 585
R12035 dvss.n3319 dvss.n3318 585
R12036 dvss.n3144 dvss.n3143 585
R12037 dvss.n3317 dvss.n3144 585
R12038 dvss.n3315 dvss.n3314 585
R12039 dvss.n3316 dvss.n3315 585
R12040 dvss.n3313 dvss.n3146 585
R12041 dvss.n3146 dvss.n3145 585
R12042 dvss.n3312 dvss.n3311 585
R12043 dvss.n3311 dvss.n3310 585
R12044 dvss.n3152 dvss.n3151 585
R12045 dvss.n3309 dvss.n3152 585
R12046 dvss.n3307 dvss.n3306 585
R12047 dvss.n3308 dvss.n3307 585
R12048 dvss.n3305 dvss.n3154 585
R12049 dvss.n3304 dvss.n3303 585
R12050 dvss.n3159 dvss.n3158 585
R12051 dvss.n3298 dvss.n3297 585
R12052 dvss.n3299 dvss.n3298 585
R12053 dvss.n3296 dvss.n3267 585
R12054 dvss.n3267 dvss.n3266 585
R12055 dvss.n3295 dvss.n3294 585
R12056 dvss.n3294 dvss.n3293 585
R12057 dvss.n3286 dvss.n3285 585
R12058 dvss.n3292 dvss.n3286 585
R12059 dvss.n3290 dvss.n3289 585
R12060 dvss.n3291 dvss.n3290 585
R12061 dvss.n1698 dvss.n1697 585
R12062 dvss.n1697 dvss.n1696 585
R12063 dvss.n1598 dvss.n1597 585
R12064 dvss.n1693 dvss.n1597 585
R12065 dvss.n1694 dvss.n1691 585
R12066 dvss.n1695 dvss.n1694 585
R12067 dvss.n1703 dvss.n1690 585
R12068 dvss.n1692 dvss.n1690 585
R12069 dvss.n1770 dvss.n1769 585
R12070 dvss.n1562 dvss.n1559 585
R12071 dvss.n1586 dvss.n1558 585
R12072 dvss.n1772 dvss.n1558 585
R12073 dvss.n1556 dvss.n1555 585
R12074 dvss.n1776 dvss.n1774 585
R12075 dvss.n1775 dvss.n1549 585
R12076 dvss.n1577 dvss.n1549 585
R12077 dvss.n1793 dvss.n1550 585
R12078 dvss.n1793 dvss.n1792 585
R12079 dvss.n1794 dvss.n1545 585
R12080 dvss.n1795 dvss.n1794 585
R12081 dvss.n1801 dvss.n1546 585
R12082 dvss.n1797 dvss.n1546 585
R12083 dvss.n1802 dvss.n1539 585
R12084 dvss.n1796 dvss.n1539 585
R12085 dvss.n1815 dvss.n1540 585
R12086 dvss.n1815 dvss.n1814 585
R12087 dvss.n1816 dvss.n1534 585
R12088 dvss.n1817 dvss.n1816 585
R12089 dvss.n1824 dvss.n1535 585
R12090 dvss.n1820 dvss.n1535 585
R12091 dvss.n1825 dvss.n1529 585
R12092 dvss.n1538 dvss.n1529 585
R12093 dvss.n1835 dvss.n1528 585
R12094 dvss.n1835 dvss.n1834 585
R12095 dvss.n1837 dvss.n1836 585
R12096 dvss.n1836 dvss.n1524 585
R12097 dvss.n1525 dvss.n1518 585
R12098 dvss.n1848 dvss.n1525 585
R12099 dvss.n1859 dvss.n1519 585
R12100 dvss.n1849 dvss.n1519 585
R12101 dvss.n1858 dvss.n1520 585
R12102 dvss.n1853 dvss.n1520 585
R12103 dvss.n1850 dvss.n1521 585
R12104 dvss.n1852 dvss.n1850 585
R12105 dvss.n1508 dvss.n1507 585
R12106 dvss.n1851 dvss.n1507 585
R12107 dvss.n1872 dvss.n1871 585
R12108 dvss.n1873 dvss.n1872 585
R12109 dvss.n1494 dvss.n1493 585
R12110 dvss.n1874 dvss.n1493 585
R12111 dvss.n1886 dvss.n1885 585
R12112 dvss.n1495 dvss.n1492 585
R12113 dvss.n1490 dvss.n1489 585
R12114 dvss.n1891 dvss.n1890 585
R12115 dvss.n1486 dvss.n1485 585
R12116 dvss.n1502 dvss.n1485 585
R12117 dvss.n1900 dvss.n1899 585
R12118 dvss.n1901 dvss.n1900 585
R12119 dvss.n1482 dvss.n1481 585
R12120 dvss.n1902 dvss.n1481 585
R12121 dvss.n1913 dvss.n1912 585
R12122 dvss.n1914 dvss.n1913 585
R12123 dvss.n1475 dvss.n1474 585
R12124 dvss.n1915 dvss.n1474 585
R12125 dvss.n1928 dvss.n1927 585
R12126 dvss.n1929 dvss.n1928 585
R12127 dvss.n1468 dvss.n1467 585
R12128 dvss.n1931 dvss.n1468 585
R12129 dvss.n1936 dvss.n1935 585
R12130 dvss.n1935 dvss.n1934 585
R12131 dvss.n1470 dvss.n1462 585
R12132 dvss.n1470 dvss.n1469 585
R12133 dvss.n1980 dvss.n1457 585
R12134 dvss.n1984 dvss.n1457 585
R12135 dvss.n1979 dvss.n1463 585
R12136 dvss.n1954 dvss.n1463 585
R12137 dvss.n1956 dvss.n1464 585
R12138 dvss.n1956 dvss.n1955 585
R12139 dvss.n1957 dvss.n1950 585
R12140 dvss.n1958 dvss.n1957 585
R12141 dvss.n1966 dvss.n1951 585
R12142 dvss.n1961 dvss.n1951 585
R12143 dvss.n1965 dvss.n1963 585
R12144 dvss.n1963 dvss.n1962 585
R12145 dvss.n1456 dvss.n1446 585
R12146 dvss.n2018 dvss.n1456 585
R12147 dvss.n2026 dvss.n1447 585
R12148 dvss.n1447 dvss.n1440 585
R12149 dvss.n2051 dvss.n1441 585
R12150 dvss.n2055 dvss.n1441 585
R12151 dvss.n2050 dvss.n2027 585
R12152 dvss.n2041 dvss.n2028 585
R12153 dvss.n2046 dvss.n2045 585
R12154 dvss.n1437 dvss.n1436 585
R12155 dvss.n2060 dvss.n2059 585
R12156 dvss.n2059 dvss.n2058 585
R12157 dvss.n1432 dvss.n1431 585
R12158 dvss.n2057 dvss.n1431 585
R12159 dvss.n2068 dvss.n2067 585
R12160 dvss.n2069 dvss.n2068 585
R12161 dvss.n1424 dvss.n1423 585
R12162 dvss.n1423 dvss.n1422 585
R12163 dvss.n2081 dvss.n2080 585
R12164 dvss.n2082 dvss.n2081 585
R12165 dvss.n1415 dvss.n1414 585
R12166 dvss.n2083 dvss.n1415 585
R12167 dvss.n2088 dvss.n2087 585
R12168 dvss.n2087 dvss.n2086 585
R12169 dvss.n1416 dvss.n1356 585
R12170 dvss.n1417 dvss.n1416 585
R12171 dvss.n2100 dvss.n1350 585
R12172 dvss.n2104 dvss.n1350 585
R12173 dvss.n2099 dvss.n1357 585
R12174 dvss.n1357 dvss.n1349 585
R12175 dvss.n1379 dvss.n1358 585
R12176 dvss.n1380 dvss.n1379 585
R12177 dvss.n1368 dvss.n1367 585
R12178 dvss.n1381 dvss.n1367 585
R12179 dvss.n1391 dvss.n1390 585
R12180 dvss.n1392 dvss.n1391 585
R12181 dvss.n1363 dvss.n1362 585
R12182 dvss.n1393 dvss.n1363 585
R12183 dvss.n1398 dvss.n1397 585
R12184 dvss.n1397 dvss.n1396 585
R12185 dvss.n1364 dvss.n896 585
R12186 dvss.n1364 dvss.n888 585
R12187 dvss.n5726 dvss.n889 585
R12188 dvss.n5730 dvss.n889 585
R12189 dvss.n5725 dvss.n897 585
R12190 dvss.n897 dvss.n890 585
R12191 dvss.n1009 dvss.n898 585
R12192 dvss.n5721 dvss.n901 585
R12193 dvss.n5720 dvss.n902 585
R12194 dvss.n1013 dvss.n903 585
R12195 dvss.n1014 dvss.n910 585
R12196 dvss.n1015 dvss.n1014 585
R12197 dvss.n5713 dvss.n911 585
R12198 dvss.n1016 dvss.n911 585
R12199 dvss.n5712 dvss.n912 585
R12200 dvss.n1019 dvss.n912 585
R12201 dvss.n1021 dvss.n913 585
R12202 dvss.n1021 dvss.n1020 585
R12203 dvss.n1022 dvss.n921 585
R12204 dvss.n1023 dvss.n1022 585
R12205 dvss.n5704 dvss.n922 585
R12206 dvss.n1027 dvss.n922 585
R12207 dvss.n5703 dvss.n923 585
R12208 dvss.n992 dvss.n923 585
R12209 dvss.n1031 dvss.n924 585
R12210 dvss.n1031 dvss.n1030 585
R12211 dvss.n1032 dvss.n930 585
R12212 dvss.n1033 dvss.n1032 585
R12213 dvss.n5693 dvss.n931 585
R12214 dvss.n1035 dvss.n931 585
R12215 dvss.n5692 dvss.n932 585
R12216 dvss.n989 dvss.n932 585
R12217 dvss.n988 dvss.n933 585
R12218 dvss.n1039 dvss.n988 585
R12219 dvss.n1042 dvss.n1041 585
R12220 dvss.n1041 dvss.n1040 585
R12221 dvss.n1043 dvss.n976 585
R12222 dvss.n1047 dvss.n976 585
R12223 dvss.n1049 dvss.n977 585
R12224 dvss.n1049 dvss.n1048 585
R12225 dvss.n1050 dvss.n945 585
R12226 dvss.n1051 dvss.n1050 585
R12227 dvss.n5677 dvss.n946 585
R12228 dvss.n1054 dvss.n946 585
R12229 dvss.n5676 dvss.n947 585
R12230 dvss.n1055 dvss.n947 585
R12231 dvss.n5647 dvss.n1078 585
R12232 dvss.n1119 dvss.n1078 585
R12233 dvss.n5646 dvss.n1079 585
R12234 dvss.n1121 dvss.n1079 585
R12235 dvss.n5611 dvss.n1080 585
R12236 dvss.n5612 dvss.n5611 585
R12237 dvss.n5639 dvss.n1102 585
R12238 dvss.n5615 dvss.n1102 585
R12239 dvss.n5638 dvss.n1103 585
R12240 dvss.n5616 dvss.n1103 585
R12241 dvss.n5617 dvss.n1104 585
R12242 dvss.n5618 dvss.n5617 585
R12243 dvss.n5626 dvss.n1110 585
R12244 dvss.n5621 dvss.n1110 585
R12245 dvss.n5625 dvss.n5623 585
R12246 dvss.n5623 dvss.n5622 585
R12247 dvss.n806 dvss.n796 585
R12248 dvss.n6121 dvss.n806 585
R12249 dvss.n6129 dvss.n797 585
R12250 dvss.n797 dvss.n790 585
R12251 dvss.n6154 dvss.n791 585
R12252 dvss.n6158 dvss.n791 585
R12253 dvss.n6153 dvss.n6130 585
R12254 dvss.n6144 dvss.n6131 585
R12255 dvss.n6149 dvss.n6148 585
R12256 dvss.n787 dvss.n786 585
R12257 dvss.n6163 dvss.n6162 585
R12258 dvss.n6162 dvss.n6161 585
R12259 dvss.n782 dvss.n781 585
R12260 dvss.n6160 dvss.n781 585
R12261 dvss.n6171 dvss.n6170 585
R12262 dvss.n6172 dvss.n6171 585
R12263 dvss.n774 dvss.n773 585
R12264 dvss.n773 dvss.n772 585
R12265 dvss.n6184 dvss.n6183 585
R12266 dvss.n6185 dvss.n6184 585
R12267 dvss.n765 dvss.n764 585
R12268 dvss.n6186 dvss.n765 585
R12269 dvss.n6191 dvss.n6190 585
R12270 dvss.n6190 dvss.n6189 585
R12271 dvss.n766 dvss.n533 585
R12272 dvss.n767 dvss.n766 585
R12273 dvss.n6203 dvss.n527 585
R12274 dvss.n6207 dvss.n527 585
R12275 dvss.n6202 dvss.n534 585
R12276 dvss.n534 dvss.n526 585
R12277 dvss.n630 dvss.n535 585
R12278 dvss.n630 dvss.n629 585
R12279 dvss.n631 dvss.n619 585
R12280 dvss.n633 dvss.n631 585
R12281 dvss.n642 dvss.n620 585
R12282 dvss.n632 dvss.n620 585
R12283 dvss.n643 dvss.n612 585
R12284 dvss.n647 dvss.n612 585
R12285 dvss.n649 dvss.n613 585
R12286 dvss.n649 dvss.n648 585
R12287 dvss.n650 dvss.n540 585
R12288 dvss.n651 dvss.n650 585
R12289 dvss.n754 dvss.n541 585
R12290 dvss.n609 dvss.n541 585
R12291 dvss.n753 dvss.n542 585
R12292 dvss.n661 dvss.n542 585
R12293 dvss.n664 dvss.n543 585
R12294 dvss.n749 dvss.n547 585
R12295 dvss.n748 dvss.n548 585
R12296 dvss.n668 dvss.n549 585
R12297 dvss.n669 dvss.n556 585
R12298 dvss.n670 dvss.n669 585
R12299 dvss.n741 dvss.n557 585
R12300 dvss.n671 dvss.n557 585
R12301 dvss.n740 dvss.n558 585
R12302 dvss.n674 dvss.n558 585
R12303 dvss.n676 dvss.n559 585
R12304 dvss.n676 dvss.n675 585
R12305 dvss.n677 dvss.n567 585
R12306 dvss.n678 dvss.n677 585
R12307 dvss.n732 dvss.n568 585
R12308 dvss.n682 dvss.n568 585
R12309 dvss.n731 dvss.n569 585
R12310 dvss.n600 dvss.n569 585
R12311 dvss.n686 dvss.n570 585
R12312 dvss.n686 dvss.n685 585
R12313 dvss.n687 dvss.n576 585
R12314 dvss.n688 dvss.n687 585
R12315 dvss.n721 dvss.n577 585
R12316 dvss.n690 dvss.n577 585
R12317 dvss.n720 dvss.n578 585
R12318 dvss.n597 dvss.n578 585
R12319 dvss.n695 dvss.n579 585
R12320 dvss.n695 dvss.n694 585
R12321 dvss.n697 dvss.n696 585
R12322 dvss.n698 dvss.n697 585
R12323 dvss.n591 dvss.n590 585
R12324 dvss.n699 dvss.n591 585
R12325 dvss.n704 dvss.n703 585
R12326 dvss.n703 dvss.n702 585
R12327 dvss.n592 dvss.n130 585
R12328 dvss.n592 dvss.n122 585
R12329 dvss.n6710 dvss.n123 585
R12330 dvss.n6714 dvss.n123 585
R12331 dvss.n6709 dvss.n131 585
R12332 dvss.n131 dvss.n124 585
R12333 dvss.n191 dvss.n132 585
R12334 dvss.n6705 dvss.n135 585
R12335 dvss.n6704 dvss.n136 585
R12336 dvss.n195 dvss.n137 585
R12337 dvss.n196 dvss.n144 585
R12338 dvss.n206 dvss.n196 585
R12339 dvss.n6697 dvss.n145 585
R12340 dvss.n207 dvss.n145 585
R12341 dvss.n6696 dvss.n146 585
R12342 dvss.n208 dvss.n146 585
R12343 dvss.n186 dvss.n147 585
R12344 dvss.n186 dvss.n185 585
R12345 dvss.n187 dvss.n155 585
R12346 dvss.n216 dvss.n187 585
R12347 dvss.n6688 dvss.n156 585
R12348 dvss.n217 dvss.n156 585
R12349 dvss.n6687 dvss.n157 585
R12350 dvss.n219 dvss.n157 585
R12351 dvss.n223 dvss.n158 585
R12352 dvss.n223 dvss.n222 585
R12353 dvss.n224 dvss.n164 585
R12354 dvss.n225 dvss.n224 585
R12355 dvss.n6677 dvss.n165 585
R12356 dvss.n6648 dvss.n165 585
R12357 dvss.n6676 dvss.n166 585
R12358 dvss.n6651 dvss.n166 585
R12359 dvss.n6653 dvss.n167 585
R12360 dvss.n6653 dvss.n6652 585
R12361 dvss.n6654 dvss.n177 585
R12362 dvss.n6655 dvss.n6654 585
R12363 dvss.n6663 dvss.n178 585
R12364 dvss.n6658 dvss.n178 585
R12365 dvss.n6662 dvss.n6660 585
R12366 dvss.n6660 dvss.n6659 585
R12367 dvss.n77 dvss.n72 585
R12368 dvss.n6862 dvss.n77 585
R12369 dvss.n6870 dvss.n73 585
R12370 dvss.n73 dvss.n66 585
R12371 dvss.n6895 dvss.n67 585
R12372 dvss.n6899 dvss.n67 585
R12373 dvss.n6894 dvss.n6871 585
R12374 dvss.n6885 dvss.n6872 585
R12375 dvss.n6890 dvss.n6889 585
R12376 dvss.n63 dvss.n62 585
R12377 dvss.n6904 dvss.n6903 585
R12378 dvss.n6903 dvss.n6902 585
R12379 dvss.n58 dvss.n57 585
R12380 dvss.n6901 dvss.n57 585
R12381 dvss.n6912 dvss.n6911 585
R12382 dvss.n6913 dvss.n6912 585
R12383 dvss.n50 dvss.n49 585
R12384 dvss.n49 dvss.n48 585
R12385 dvss.n6925 dvss.n6924 585
R12386 dvss.n6926 dvss.n6925 585
R12387 dvss.n41 dvss.n40 585
R12388 dvss.n6927 dvss.n41 585
R12389 dvss.n6932 dvss.n6931 585
R12390 dvss.n6931 dvss.n6930 585
R12391 dvss.n42 dvss.n31 585
R12392 dvss.n43 dvss.n42 585
R12393 dvss.n6944 dvss.n25 585
R12394 dvss.n6948 dvss.n25 585
R12395 dvss.n6943 dvss.n32 585
R12396 dvss.n32 dvss.n24 585
R12397 dvss.n6455 dvss.n33 585
R12398 dvss.n6459 dvss.n6455 585
R12399 dvss.n6462 dvss.n6461 585
R12400 dvss.n6461 dvss.n6460 585
R12401 dvss.n6445 dvss.n6444 585
R12402 dvss.n6471 dvss.n6445 585
R12403 dvss.n6474 dvss.n6473 585
R12404 dvss.n6473 dvss.n6472 585
R12405 dvss.n6441 dvss.n6440 585
R12406 dvss.n6479 dvss.n6441 585
R12407 dvss.n6482 dvss.n6481 585
R12408 dvss.n6481 dvss.n6480 585
R12409 dvss.n6436 dvss.n6435 585
R12410 dvss.n6437 dvss.n6436 585
R12411 dvss.n6493 dvss.n6492 585
R12412 dvss.n6492 dvss.n6491 585
R12413 dvss.n6432 dvss.n6431 585
R12414 dvss.n6431 dvss.n6429 585
R12415 dvss.n6500 dvss.n6499 585
R12416 dvss.n6501 dvss.n6500 585
R12417 dvss.n5669 dvss.n948 585
R12418 dvss.n5672 dvss.n5671 585
R12419 dvss.n955 dvss.n952 585
R12420 dvss.n5666 dvss.n5665 585
R12421 dvss.n1057 dvss.n950 585
R12422 dvss.n973 dvss.n951 585
R12423 dvss.n970 dvss.n969 585
R12424 dvss.n1062 dvss.n1061 585
R12425 dvss.n5664 dvss.n954 585
R12426 dvss.n971 dvss.n954 585
R12427 dvss.n5663 dvss.n5662 585
R12428 dvss.n5662 dvss.n5661 585
R12429 dvss.n965 dvss.n964 585
R12430 dvss.n1068 dvss.n965 585
R12431 dvss.n1088 dvss.n1069 585
R12432 dvss.n5655 dvss.n1069 585
R12433 dvss.n1090 dvss.n1070 585
R12434 dvss.n5654 dvss.n1070 585
R12435 dvss.n1089 dvss.n1071 585
R12436 dvss.n5653 dvss.n1071 585
R12437 dvss.n1116 dvss.n1077 585
R12438 dvss.n1117 dvss.n1116 585
R12439 dvss.n1063 dvss.n966 585
R12440 dvss.n971 dvss.n966 585
R12441 dvss.n5660 dvss.n5659 585
R12442 dvss.n5661 dvss.n5660 585
R12443 dvss.n5658 dvss.n967 585
R12444 dvss.n1068 dvss.n967 585
R12445 dvss.n5657 dvss.n5656 585
R12446 dvss.n5656 dvss.n5655 585
R12447 dvss.n1067 dvss.n1066 585
R12448 dvss.n5654 dvss.n1067 585
R12449 dvss.n5652 dvss.n5651 585
R12450 dvss.n5653 dvss.n5652 585
R12451 dvss.n5650 dvss.n1072 585
R12452 dvss.n1117 dvss.n1072 585
R12453 dvss.n5509 dvss.n5508 585
R12454 dvss.n5510 dvss.n5509 585
R12455 dvss.n1144 dvss.n1143 585
R12456 dvss.n5511 dvss.n1144 585
R12457 dvss.n5514 dvss.n5513 585
R12458 dvss.n5513 dvss.n5512 585
R12459 dvss.n1142 dvss.n1141 585
R12460 dvss.n1141 dvss.n1140 585
R12461 dvss.n5520 dvss.n5519 585
R12462 dvss.n5521 dvss.n5520 585
R12463 dvss.n1139 dvss.n1138 585
R12464 dvss.n5522 dvss.n1139 585
R12465 dvss.n5525 dvss.n5524 585
R12466 dvss.n5524 dvss.n5523 585
R12467 dvss.n1126 dvss.n1124 585
R12468 dvss.n1124 dvss.n1122 585
R12469 dvss.n5608 dvss.n5607 585
R12470 dvss.n5609 dvss.n5608 585
R12471 dvss.n5606 dvss.n1125 585
R12472 dvss.n1125 dvss.n1123 585
R12473 dvss.n5605 dvss.n5604 585
R12474 dvss.n1131 dvss.n1130 585
R12475 dvss.n5600 dvss.n5599 585
R12476 dvss.n5601 dvss.n5600 585
R12477 dvss.n5598 dvss.n1133 585
R12478 dvss.n5542 dvss.n1133 585
R12479 dvss.n5597 dvss.n5596 585
R12480 dvss.n5596 dvss.n5595 585
R12481 dvss.n5541 dvss.n5540 585
R12482 dvss.n5594 dvss.n5541 585
R12483 dvss.n5592 dvss.n5591 585
R12484 dvss.n5593 dvss.n5592 585
R12485 dvss.n5590 dvss.n5544 585
R12486 dvss.n5544 dvss.n5543 585
R12487 dvss.n5589 dvss.n5588 585
R12488 dvss.n5588 dvss.n5587 585
R12489 dvss.n5550 dvss.n5549 585
R12490 dvss.n5586 dvss.n5550 585
R12491 dvss.n5584 dvss.n5583 585
R12492 dvss.n5585 dvss.n5584 585
R12493 dvss.n5582 dvss.n5551 585
R12494 dvss.n5563 dvss.n5551 585
R12495 dvss.n5581 dvss.n5580 585
R12496 dvss.n5580 dvss.n5579 585
R12497 dvss.n5562 dvss.n5561 585
R12498 dvss.n5578 dvss.n5562 585
R12499 dvss.n5576 dvss.n5575 585
R12500 dvss.n5577 dvss.n5576 585
R12501 dvss.n5574 dvss.n5565 585
R12502 dvss.n5565 dvss.n5564 585
R12503 dvss.n3128 dvss.n3127 585
R12504 dvss.n5492 dvss.n1207 585
R12505 dvss.n5491 dvss.n1206 585
R12506 dvss.n5495 dvss.n1206 585
R12507 dvss.n5490 dvss.n5489 585
R12508 dvss.n5488 dvss.n5487 585
R12509 dvss.n5486 dvss.n5485 585
R12510 dvss.n5484 dvss.n5483 585
R12511 dvss.n5482 dvss.n5481 585
R12512 dvss.n5480 dvss.n5479 585
R12513 dvss.n5478 dvss.n5477 585
R12514 dvss.n5476 dvss.n5475 585
R12515 dvss.n5474 dvss.n5473 585
R12516 dvss.n5472 dvss.n5471 585
R12517 dvss.n5470 dvss.n5469 585
R12518 dvss.n5468 dvss.n5467 585
R12519 dvss.n5466 dvss.n5465 585
R12520 dvss.n5464 dvss.n5463 585
R12521 dvss.n5462 dvss.n5461 585
R12522 dvss.n5460 dvss.n5459 585
R12523 dvss.n5458 dvss.n5457 585
R12524 dvss.n5456 dvss.n5455 585
R12525 dvss.n5454 dvss.n5453 585
R12526 dvss.n5452 dvss.n5451 585
R12527 dvss.n5450 dvss.n5449 585
R12528 dvss.n5448 dvss.n5447 585
R12529 dvss.n5446 dvss.n5445 585
R12530 dvss.n5444 dvss.n5443 585
R12531 dvss.n5442 dvss.n5441 585
R12532 dvss.n5440 dvss.n5439 585
R12533 dvss.n5438 dvss.n5437 585
R12534 dvss.n5436 dvss.n5435 585
R12535 dvss.n5434 dvss.n5433 585
R12536 dvss.n5432 dvss.n5431 585
R12537 dvss.n5430 dvss.n5429 585
R12538 dvss.n5428 dvss.n5427 585
R12539 dvss.n5426 dvss.n5425 585
R12540 dvss.n5424 dvss.n5423 585
R12541 dvss.n5422 dvss.n5421 585
R12542 dvss.n5420 dvss.n5419 585
R12543 dvss.n5418 dvss.n5417 585
R12544 dvss.n5416 dvss.n5415 585
R12545 dvss.n5414 dvss.n5413 585
R12546 dvss.n5412 dvss.n5411 585
R12547 dvss.n5410 dvss.n5409 585
R12548 dvss.n5408 dvss.n5407 585
R12549 dvss.n5406 dvss.n5405 585
R12550 dvss.n5404 dvss.n5403 585
R12551 dvss.n5402 dvss.n5401 585
R12552 dvss.n5400 dvss.n5399 585
R12553 dvss.n5398 dvss.n5397 585
R12554 dvss.n5396 dvss.n5395 585
R12555 dvss.n5394 dvss.n5393 585
R12556 dvss.n5392 dvss.n5391 585
R12557 dvss.n5390 dvss.n5389 585
R12558 dvss.n5388 dvss.n5387 585
R12559 dvss.n5386 dvss.n5385 585
R12560 dvss.n5384 dvss.n5383 585
R12561 dvss.n5382 dvss.n5381 585
R12562 dvss.n5380 dvss.n5379 585
R12563 dvss.n5378 dvss.n5377 585
R12564 dvss.n5376 dvss.n5375 585
R12565 dvss.n5374 dvss.n5373 585
R12566 dvss.n5372 dvss.n5371 585
R12567 dvss.n5370 dvss.n5369 585
R12568 dvss.n5368 dvss.n5367 585
R12569 dvss.n5366 dvss.n5365 585
R12570 dvss.n5364 dvss.n5363 585
R12571 dvss.n5362 dvss.n5361 585
R12572 dvss.n5360 dvss.n5359 585
R12573 dvss.n5358 dvss.n5357 585
R12574 dvss.n5356 dvss.n5355 585
R12575 dvss.n5354 dvss.n5353 585
R12576 dvss.n5352 dvss.n5351 585
R12577 dvss.n5350 dvss.n5349 585
R12578 dvss.n5348 dvss.n5347 585
R12579 dvss.n5346 dvss.n5345 585
R12580 dvss.n5344 dvss.n5343 585
R12581 dvss.n5342 dvss.n5341 585
R12582 dvss.n5340 dvss.n5339 585
R12583 dvss.n5338 dvss.n5337 585
R12584 dvss.n5336 dvss.n5335 585
R12585 dvss.n5334 dvss.n5333 585
R12586 dvss.n5332 dvss.n5331 585
R12587 dvss.n5330 dvss.n5329 585
R12588 dvss.n5328 dvss.n5327 585
R12589 dvss.n5326 dvss.n5325 585
R12590 dvss.n5324 dvss.n5323 585
R12591 dvss.n5322 dvss.n5321 585
R12592 dvss.n5320 dvss.n5319 585
R12593 dvss.n5318 dvss.n5317 585
R12594 dvss.n5316 dvss.n5315 585
R12595 dvss.n5314 dvss.n5313 585
R12596 dvss.n5312 dvss.n5311 585
R12597 dvss.n5310 dvss.n5309 585
R12598 dvss.n5308 dvss.n5307 585
R12599 dvss.n5306 dvss.n5305 585
R12600 dvss.n5304 dvss.n5303 585
R12601 dvss.n5302 dvss.n5301 585
R12602 dvss.n5300 dvss.n5299 585
R12603 dvss.n5298 dvss.n5297 585
R12604 dvss.n5296 dvss.n5295 585
R12605 dvss.n5294 dvss.n5293 585
R12606 dvss.n5292 dvss.n5291 585
R12607 dvss.n5290 dvss.n5289 585
R12608 dvss.n5288 dvss.n5287 585
R12609 dvss.n1152 dvss.n1149 585
R12610 dvss.n5498 dvss.n5497 585
R12611 dvss.n1151 dvss.n1150 585
R12612 dvss.n1147 dvss.n1146 585
R12613 dvss.n1728 dvss.n1727 585
R12614 dvss.n1726 dvss.n1689 585
R12615 dvss.n1725 dvss.n1688 585
R12616 dvss.n1730 dvss.n1688 585
R12617 dvss.n1724 dvss.n1723 585
R12618 dvss.n1722 dvss.n1721 585
R12619 dvss.n1720 dvss.n1719 585
R12620 dvss.n1718 dvss.n1717 585
R12621 dvss.n1716 dvss.n1715 585
R12622 dvss.n1623 dvss.n1619 585
R12623 dvss.n1733 dvss.n1732 585
R12624 dvss.n1624 dvss.n1622 585
R12625 dvss.n1561 dvss.n1560 585
R12626 dvss.n1730 dvss.n1560 585
R12627 dvss.n1753 dvss.n1752 585
R12628 dvss.n1751 dvss.n1596 585
R12629 dvss.n1750 dvss.n1595 585
R12630 dvss.n1755 dvss.n1595 585
R12631 dvss.n1749 dvss.n1748 585
R12632 dvss.n1747 dvss.n1746 585
R12633 dvss.n1745 dvss.n1744 585
R12634 dvss.n1743 dvss.n1742 585
R12635 dvss.n1741 dvss.n1740 585
R12636 dvss.n1739 dvss.n1738 585
R12637 dvss.n1737 dvss.n1736 585
R12638 dvss.n1568 dvss.n1566 585
R12639 dvss.n1757 dvss.n1756 585
R12640 dvss.n1756 dvss.n1755 585
R12641 dvss.n2293 dvss.n0 585
R12642 dvss.n2294 dvss.n2293 585
R12643 dvss.n7055 dvss.n1 585
R12644 dvss.n2292 dvss.n1 585
R12645 dvss.n7054 dvss.n2 585
R12646 dvss.n2291 dvss.n2 585
R12647 dvss.n2289 dvss.n3 585
R12648 dvss.n2290 dvss.n2289 585
R12649 dvss.n2288 dvss.n2287 585
R12650 dvss.n2288 dvss.n1240 585
R12651 dvss.n1242 dvss.n1241 585
R12652 dvss.n1628 dvss.n1241 585
R12653 dvss.n2283 dvss.n1243 585
R12654 dvss.n1629 dvss.n1243 585
R12655 dvss.n2282 dvss.n1244 585
R12656 dvss.n1630 dvss.n1244 585
R12657 dvss.n1684 dvss.n1245 585
R12658 dvss.n1685 dvss.n1684 585
R12659 dvss.n2276 dvss.n1247 585
R12660 dvss.n1683 dvss.n1247 585
R12661 dvss.n2275 dvss.n1248 585
R12662 dvss.n1682 dvss.n1248 585
R12663 dvss.n1680 dvss.n1249 585
R12664 dvss.n1681 dvss.n1680 585
R12665 dvss.n2268 dvss.n1252 585
R12666 dvss.n1679 dvss.n1252 585
R12667 dvss.n2267 dvss.n1253 585
R12668 dvss.n1678 dvss.n1253 585
R12669 dvss.n1676 dvss.n1254 585
R12670 dvss.n1677 dvss.n1676 585
R12671 dvss.n2261 dvss.n1257 585
R12672 dvss.n1675 dvss.n1257 585
R12673 dvss.n2260 dvss.n1258 585
R12674 dvss.n1674 dvss.n1258 585
R12675 dvss.n1672 dvss.n1259 585
R12676 dvss.n1673 dvss.n1672 585
R12677 dvss.n2256 dvss.n1260 585
R12678 dvss.n1671 dvss.n1260 585
R12679 dvss.n2255 dvss.n1261 585
R12680 dvss.n1670 dvss.n1261 585
R12681 dvss.n1668 dvss.n1262 585
R12682 dvss.n1669 dvss.n1668 585
R12683 dvss.n1667 dvss.n1265 585
R12684 dvss.n2247 dvss.n1266 585
R12685 dvss.n1631 dvss.n1266 585
R12686 dvss.n2246 dvss.n1267 585
R12687 dvss.n1632 dvss.n1267 585
R12688 dvss.n1633 dvss.n1268 585
R12689 dvss.n2238 dvss.n1272 585
R12690 dvss.n1634 dvss.n1272 585
R12691 dvss.n2237 dvss.n1273 585
R12692 dvss.n1635 dvss.n1273 585
R12693 dvss.n1663 dvss.n1274 585
R12694 dvss.n1664 dvss.n1663 585
R12695 dvss.n2230 dvss.n1276 585
R12696 dvss.n1662 dvss.n1276 585
R12697 dvss.n2229 dvss.n1277 585
R12698 dvss.n1661 dvss.n1277 585
R12699 dvss.n1659 dvss.n1278 585
R12700 dvss.n1660 dvss.n1659 585
R12701 dvss.n1658 dvss.n1282 585
R12702 dvss.n1658 dvss.n1657 585
R12703 dvss.n2220 dvss.n1283 585
R12704 dvss.n1656 dvss.n1283 585
R12705 dvss.n2219 dvss.n1284 585
R12706 dvss.n1655 dvss.n1284 585
R12707 dvss.n1653 dvss.n1285 585
R12708 dvss.n1654 dvss.n1653 585
R12709 dvss.n2215 dvss.n1286 585
R12710 dvss.n1651 dvss.n1286 585
R12711 dvss.n2214 dvss.n1287 585
R12712 dvss.n1650 dvss.n1287 585
R12713 dvss.n1646 dvss.n1288 585
R12714 dvss.n2210 dvss.n1289 585
R12715 dvss.n2209 dvss.n1290 585
R12716 dvss.n1644 dvss.n1291 585
R12717 dvss.n2205 dvss.n1292 585
R12718 dvss.n1643 dvss.n1292 585
R12719 dvss.n2204 dvss.n1293 585
R12720 dvss.n1642 dvss.n1293 585
R12721 dvss.n1640 dvss.n1294 585
R12722 dvss.n2197 dvss.n1297 585
R12723 dvss.n1639 dvss.n1297 585
R12724 dvss.n2196 dvss.n1298 585
R12725 dvss.n1638 dvss.n1298 585
R12726 dvss.n1636 dvss.n1299 585
R12727 dvss.n2188 dvss.n1303 585
R12728 dvss.n1986 dvss.n1303 585
R12729 dvss.n2187 dvss.n1304 585
R12730 dvss.n1987 dvss.n1304 585
R12731 dvss.n1988 dvss.n1305 585
R12732 dvss.n1989 dvss.n1988 585
R12733 dvss.n2180 dvss.n1307 585
R12734 dvss.n1990 dvss.n1307 585
R12735 dvss.n2179 dvss.n1308 585
R12736 dvss.n1991 dvss.n1308 585
R12737 dvss.n1993 dvss.n1309 585
R12738 dvss.n1993 dvss.n1992 585
R12739 dvss.n1994 dvss.n1313 585
R12740 dvss.n1995 dvss.n1994 585
R12741 dvss.n2170 dvss.n1314 585
R12742 dvss.n1996 dvss.n1314 585
R12743 dvss.n2169 dvss.n1315 585
R12744 dvss.n1997 dvss.n1315 585
R12745 dvss.n1998 dvss.n1316 585
R12746 dvss.n1999 dvss.n1998 585
R12747 dvss.n2160 dvss.n1317 585
R12748 dvss.n2015 dvss.n1317 585
R12749 dvss.n2159 dvss.n1318 585
R12750 dvss.n2014 dvss.n1318 585
R12751 dvss.n2002 dvss.n1319 585
R12752 dvss.n2155 dvss.n1320 585
R12753 dvss.n2154 dvss.n1321 585
R12754 dvss.n2000 dvss.n1322 585
R12755 dvss.n2150 dvss.n1323 585
R12756 dvss.n2012 dvss.n1323 585
R12757 dvss.n2149 dvss.n1324 585
R12758 dvss.n2011 dvss.n1324 585
R12759 dvss.n2009 dvss.n1325 585
R12760 dvss.n2142 dvss.n1328 585
R12761 dvss.n2005 dvss.n1328 585
R12762 dvss.n2141 dvss.n1329 585
R12763 dvss.n2006 dvss.n1329 585
R12764 dvss.n2007 dvss.n1330 585
R12765 dvss.n2133 dvss.n1334 585
R12766 dvss.n1348 dvss.n1334 585
R12767 dvss.n2132 dvss.n1335 585
R12768 dvss.n1347 dvss.n1335 585
R12769 dvss.n2106 dvss.n1336 585
R12770 dvss.n2107 dvss.n2106 585
R12771 dvss.n2125 dvss.n1338 585
R12772 dvss.n2108 dvss.n1338 585
R12773 dvss.n2124 dvss.n1339 585
R12774 dvss.n2109 dvss.n1339 585
R12775 dvss.n2110 dvss.n1340 585
R12776 dvss.n2111 dvss.n2110 585
R12777 dvss.n1346 dvss.n1345 585
R12778 dvss.n2112 dvss.n1346 585
R12779 dvss.n2115 dvss.n2114 585
R12780 dvss.n2114 dvss.n2113 585
R12781 dvss.n886 dvss.n885 585
R12782 dvss.n887 dvss.n886 585
R12783 dvss.n5735 dvss.n5734 585
R12784 dvss.n5734 dvss.n5733 585
R12785 dvss.n878 dvss.n876 585
R12786 dvss.n876 dvss.n875 585
R12787 dvss.n5750 dvss.n5749 585
R12788 dvss.n5751 dvss.n5750 585
R12789 dvss.n879 dvss.n877 585
R12790 dvss.n5745 dvss.n5739 585
R12791 dvss.n5744 dvss.n5741 585
R12792 dvss.n873 dvss.n872 585
R12793 dvss.n5756 dvss.n5755 585
R12794 dvss.n5755 dvss.n5754 585
R12795 dvss.n870 dvss.n869 585
R12796 dvss.n5753 dvss.n869 585
R12797 dvss.n5766 dvss.n5765 585
R12798 dvss.n867 dvss.n866 585
R12799 dvss.n868 dvss.n867 585
R12800 dvss.n5771 dvss.n5770 585
R12801 dvss.n5770 dvss.n5769 585
R12802 dvss.n864 dvss.n863 585
R12803 dvss.n5784 dvss.n5783 585
R12804 dvss.n5785 dvss.n5784 585
R12805 dvss.n861 dvss.n860 585
R12806 dvss.n5786 dvss.n861 585
R12807 dvss.n5789 dvss.n5788 585
R12808 dvss.n5788 dvss.n5787 585
R12809 dvss.n859 dvss.n858 585
R12810 dvss.n858 dvss.n857 585
R12811 dvss.n5798 dvss.n5797 585
R12812 dvss.n5799 dvss.n5798 585
R12813 dvss.n856 dvss.n855 585
R12814 dvss.n5800 dvss.n856 585
R12815 dvss.n5803 dvss.n5802 585
R12816 dvss.n5802 dvss.n5801 585
R12817 dvss.n852 dvss.n851 585
R12818 dvss.n851 dvss.n850 585
R12819 dvss.n5819 dvss.n5818 585
R12820 dvss.n5820 dvss.n5819 585
R12821 dvss.n848 dvss.n847 585
R12822 dvss.n5821 dvss.n848 585
R12823 dvss.n5826 dvss.n5825 585
R12824 dvss.n5825 dvss.n5824 585
R12825 dvss.n846 dvss.n845 585
R12826 dvss.n5823 dvss.n845 585
R12827 dvss.n5832 dvss.n5831 585
R12828 dvss.n844 dvss.n843 585
R12829 dvss.n5837 dvss.n5836 585
R12830 dvss.n842 dvss.n841 585
R12831 dvss.n5844 dvss.n5843 585
R12832 dvss.n5845 dvss.n5844 585
R12833 dvss.n839 dvss.n838 585
R12834 dvss.n5846 dvss.n839 585
R12835 dvss.n5849 dvss.n5848 585
R12836 dvss.n834 dvss.n833 585
R12837 dvss.n833 dvss.n832 585
R12838 dvss.n5859 dvss.n5858 585
R12839 dvss.n5860 dvss.n5859 585
R12840 dvss.n831 dvss.n830 585
R12841 dvss.n5865 dvss.n5864 585
R12842 dvss.n5864 dvss.n5863 585
R12843 dvss.n824 dvss.n823 585
R12844 dvss.n5862 dvss.n823 585
R12845 dvss.n5874 dvss.n5873 585
R12846 dvss.n5875 dvss.n5874 585
R12847 dvss.n822 dvss.n821 585
R12848 dvss.n5876 dvss.n822 585
R12849 dvss.n5880 dvss.n5879 585
R12850 dvss.n5879 dvss.n5878 585
R12851 dvss.n816 dvss.n815 585
R12852 dvss.n5877 dvss.n815 585
R12853 dvss.n5889 dvss.n5888 585
R12854 dvss.n5890 dvss.n5889 585
R12855 dvss.n814 dvss.n813 585
R12856 dvss.n5891 dvss.n814 585
R12857 dvss.n5894 dvss.n5893 585
R12858 dvss.n5893 dvss.n5892 585
R12859 dvss.n811 dvss.n809 585
R12860 dvss.n809 dvss.n807 585
R12861 dvss.n6117 dvss.n6116 585
R12862 dvss.n6118 dvss.n6117 585
R12863 dvss.n812 dvss.n810 585
R12864 dvss.n810 dvss.n808 585
R12865 dvss.n6112 dvss.n5902 585
R12866 dvss.n6111 dvss.n5903 585
R12867 dvss.n5919 dvss.n5904 585
R12868 dvss.n6107 dvss.n5905 585
R12869 dvss.n6106 dvss.n5906 585
R12870 dvss.n5924 dvss.n5906 585
R12871 dvss.n5926 dvss.n5907 585
R12872 dvss.n5926 dvss.n5925 585
R12873 dvss.n5927 dvss.n5910 585
R12874 dvss.n6098 dvss.n5911 585
R12875 dvss.n5929 dvss.n5911 585
R12876 dvss.n6097 dvss.n5912 585
R12877 dvss.n5930 dvss.n5912 585
R12878 dvss.n5918 dvss.n5913 585
R12879 dvss.n6089 dvss.n5917 585
R12880 dvss.n5932 dvss.n5917 585
R12881 dvss.n6088 dvss.n5934 585
R12882 dvss.n5934 dvss.n5933 585
R12883 dvss.n5977 dvss.n5935 585
R12884 dvss.n5978 dvss.n5977 585
R12885 dvss.n6081 dvss.n5937 585
R12886 dvss.n5979 dvss.n5937 585
R12887 dvss.n6080 dvss.n5938 585
R12888 dvss.n5980 dvss.n5938 585
R12889 dvss.n5982 dvss.n5939 585
R12890 dvss.n5982 dvss.n5981 585
R12891 dvss.n5983 dvss.n5943 585
R12892 dvss.n5984 dvss.n5983 585
R12893 dvss.n6071 dvss.n5944 585
R12894 dvss.n5985 dvss.n5944 585
R12895 dvss.n6070 dvss.n5945 585
R12896 dvss.n5986 dvss.n5945 585
R12897 dvss.n5987 dvss.n5946 585
R12898 dvss.n5988 dvss.n5987 585
R12899 dvss.n6066 dvss.n5947 585
R12900 dvss.n5990 dvss.n5947 585
R12901 dvss.n6065 dvss.n5948 585
R12902 dvss.n5991 dvss.n5948 585
R12903 dvss.n5994 dvss.n5949 585
R12904 dvss.n6061 dvss.n5950 585
R12905 dvss.n6060 dvss.n5951 585
R12906 dvss.n5992 dvss.n5952 585
R12907 dvss.n6056 dvss.n5953 585
R12908 dvss.n5998 dvss.n5953 585
R12909 dvss.n6055 dvss.n5954 585
R12910 dvss.n5999 dvss.n5954 585
R12911 dvss.n6000 dvss.n5955 585
R12912 dvss.n6048 dvss.n5958 585
R12913 dvss.n6002 dvss.n5958 585
R12914 dvss.n6047 dvss.n5959 585
R12915 dvss.n6003 dvss.n5959 585
R12916 dvss.n5976 dvss.n5960 585
R12917 dvss.n6039 dvss.n5964 585
R12918 dvss.n6005 dvss.n5964 585
R12919 dvss.n6038 dvss.n5965 585
R12920 dvss.n6006 dvss.n5965 585
R12921 dvss.n6007 dvss.n5966 585
R12922 dvss.n6008 dvss.n6007 585
R12923 dvss.n6031 dvss.n5968 585
R12924 dvss.n6009 dvss.n5968 585
R12925 dvss.n6030 dvss.n5969 585
R12926 dvss.n6010 dvss.n5969 585
R12927 dvss.n6012 dvss.n5970 585
R12928 dvss.n6012 dvss.n6011 585
R12929 dvss.n6013 dvss.n5974 585
R12930 dvss.n6014 dvss.n6013 585
R12931 dvss.n6021 dvss.n5975 585
R12932 dvss.n6015 dvss.n5975 585
R12933 dvss.n6020 dvss.n6017 585
R12934 dvss.n6017 dvss.n6016 585
R12935 dvss.n119 dvss.n118 585
R12936 dvss.n120 dvss.n119 585
R12937 dvss.n6720 dvss.n6719 585
R12938 dvss.n6719 dvss.n6718 585
R12939 dvss.n117 dvss.n116 585
R12940 dvss.n6717 dvss.n116 585
R12941 dvss.n6726 dvss.n6725 585
R12942 dvss.n115 dvss.n114 585
R12943 dvss.n6731 dvss.n6730 585
R12944 dvss.n113 dvss.n112 585
R12945 dvss.n6738 dvss.n6737 585
R12946 dvss.n6739 dvss.n6738 585
R12947 dvss.n110 dvss.n109 585
R12948 dvss.n6740 dvss.n110 585
R12949 dvss.n6743 dvss.n6742 585
R12950 dvss.n105 dvss.n104 585
R12951 dvss.n104 dvss.n103 585
R12952 dvss.n6753 dvss.n6752 585
R12953 dvss.n6754 dvss.n6753 585
R12954 dvss.n102 dvss.n101 585
R12955 dvss.n6759 dvss.n6758 585
R12956 dvss.n6758 dvss.n6757 585
R12957 dvss.n95 dvss.n94 585
R12958 dvss.n6756 dvss.n94 585
R12959 dvss.n6768 dvss.n6767 585
R12960 dvss.n6769 dvss.n6768 585
R12961 dvss.n93 dvss.n92 585
R12962 dvss.n6770 dvss.n93 585
R12963 dvss.n6774 dvss.n6773 585
R12964 dvss.n6773 dvss.n6772 585
R12965 dvss.n87 dvss.n86 585
R12966 dvss.n6771 dvss.n86 585
R12967 dvss.n6783 dvss.n6782 585
R12968 dvss.n6784 dvss.n6783 585
R12969 dvss.n85 dvss.n84 585
R12970 dvss.n6785 dvss.n85 585
R12971 dvss.n6788 dvss.n6787 585
R12972 dvss.n6787 dvss.n6786 585
R12973 dvss.n82 dvss.n80 585
R12974 dvss.n80 dvss.n78 585
R12975 dvss.n6858 dvss.n6857 585
R12976 dvss.n6859 dvss.n6858 585
R12977 dvss.n83 dvss.n81 585
R12978 dvss.n81 dvss.n79 585
R12979 dvss.n6853 dvss.n6791 585
R12980 dvss.n6852 dvss.n6792 585
R12981 dvss.n6807 dvss.n6793 585
R12982 dvss.n6848 dvss.n6794 585
R12983 dvss.n6847 dvss.n6795 585
R12984 dvss.n6812 dvss.n6795 585
R12985 dvss.n6814 dvss.n6796 585
R12986 dvss.n6814 dvss.n6813 585
R12987 dvss.n6815 dvss.n6799 585
R12988 dvss.n6839 dvss.n6800 585
R12989 dvss.n6817 dvss.n6800 585
R12990 dvss.n6838 dvss.n6801 585
R12991 dvss.n6806 dvss.n6801 585
R12992 dvss.n6819 dvss.n6802 585
R12993 dvss.n6830 dvss.n6821 585
R12994 dvss.n6821 dvss.n6820 585
R12995 dvss.n6829 dvss.n6822 585
R12996 dvss.n6822 dvss.n23 585
R12997 dvss.n22 dvss.n21 585
R12998 dvss.n6950 dvss.n22 585
R12999 dvss.n6953 dvss.n6952 585
R13000 dvss.n6952 dvss.n6951 585
R13001 dvss.n20 dvss.n19 585
R13002 dvss.n19 dvss.n18 585
R13003 dvss.n6966 dvss.n6965 585
R13004 dvss.n6967 dvss.n6966 585
R13005 dvss.n17 dvss.n16 585
R13006 dvss.n6968 dvss.n17 585
R13007 dvss.n6971 dvss.n6970 585
R13008 dvss.n6970 dvss.n6969 585
R13009 dvss.n14 dvss.n13 585
R13010 dvss.n13 dvss.n12 585
R13011 dvss.n6979 dvss.n6978 585
R13012 dvss.n6980 dvss.n6979 585
R13013 dvss.n15 dvss.n9 585
R13014 dvss.n6982 dvss.n9 585
R13015 dvss.n6984 dvss.n10 585
R13016 dvss.n6984 dvss.n6983 585
R13017 dvss.n6985 dvss.n7 585
R13018 dvss.n6502 dvss.n6501 583.256
R13019 dvss dvss.t1551 581.61
R13020 dvss.t404 dvss.t465 581.61
R13021 dvss.t1285 dvss 581.61
R13022 dvss.t1199 dvss.t1424 581.61
R13023 dvss.n1696 dvss.n1239 578.14
R13024 dvss.n334 dvss.t48 575.611
R13025 dvss.t1400 dvss.t1213 573.181
R13026 dvss.t738 dvss.t1403 573.181
R13027 dvss.t34 dvss.t2063 573.181
R13028 dvss dvss.t2017 573.181
R13029 dvss.t467 dvss.t410 573.181
R13030 dvss.t199 dvss.t168 573.181
R13031 dvss.t776 dvss 573.181
R13032 dvss.n6611 dvss.t1156 568.053
R13033 dvss dvss.n2305 564.751
R13034 dvss.t1985 dvss 564.751
R13035 dvss.n3125 dvss 564.751
R13036 dvss.t553 dvss 564.751
R13037 dvss dvss.n3337 564.751
R13038 dvss.t1996 dvss 564.751
R13039 dvss.n3907 dvss 564.751
R13040 dvss dvss.n3907 564.751
R13041 dvss dvss.t122 564.751
R13042 dvss.t1263 dvss.t305 564.751
R13043 dvss.t209 dvss.t463 564.751
R13044 dvss dvss.n1145 564.751
R13045 dvss.t1354 dvss 564.751
R13046 dvss dvss.n1145 564.751
R13047 dvss.t1921 dvss.t946 564.751
R13048 dvss.t900 dvss 564.751
R13049 dvss dvss.n1145 564.751
R13050 dvss.n5668 dvss.n953 564.282
R13051 dvss.n6887 dvss.n64 564.282
R13052 dvss.n666 dvss.n663 564.282
R13053 dvss.n6146 dvss.n788 564.282
R13054 dvss.n1011 dvss.n1008 564.282
R13055 dvss.n2043 dvss.n1438 564.282
R13056 dvss.n1888 dvss.n1491 564.282
R13057 dvss.n193 dvss.n190 564.282
R13058 dvss dvss.t1034 556.322
R13059 dvss.t638 dvss.t1574 556.322
R13060 dvss dvss.t2060 556.322
R13061 dvss.t392 dvss.t154 556.322
R13062 dvss.t2091 dvss.t984 556.322
R13063 dvss.t476 dvss.t470 556.322
R13064 dvss.t31 dvss.t492 556.322
R13065 dvss dvss.t2074 556.322
R13066 dvss.t215 dvss.t1279 556.322
R13067 dvss dvss.t925 547.894
R13068 dvss.t707 dvss 547.894
R13069 dvss dvss.t709 547.894
R13070 dvss.t968 dvss.t1960 547.894
R13071 dvss dvss.t462 547.894
R13072 dvss.t1323 dvss 547.894
R13073 dvss dvss.t702 547.894
R13074 dvss.t617 dvss.t35 547.894
R13075 dvss.t888 dvss.t36 547.894
R13076 dvss dvss.t494 547.894
R13077 dvss dvss.t1255 547.894
R13078 dvss.t597 dvss 547.894
R13079 dvss dvss.t2187 547.894
R13080 dvss dvss.t1046 547.894
R13081 dvss.t1970 dvss.t1134 547.894
R13082 dvss.t496 dvss 547.894
R13083 dvss.t1966 dvss.t304 547.894
R13084 dvss.t305 dvss.t956 547.894
R13085 dvss.t2140 dvss.t1288 547.894
R13086 dvss.t1176 dvss.t201 547.894
R13087 dvss.t506 dvss 547.894
R13088 dvss dvss.t1999 547.894
R13089 dvss.t1321 dvss 547.894
R13090 dvss dvss.t500 547.894
R13091 dvss dvss.t498 547.894
R13092 dvss.t1203 dvss 539.465
R13093 dvss.t37 dvss.t444 539.465
R13094 dvss dvss.t1888 539.465
R13095 dvss.t1579 dvss 539.465
R13096 dvss.t1990 dvss 539.465
R13097 dvss.t603 dvss.t1222 539.465
R13098 dvss dvss.t100 539.465
R13099 dvss.n3629 dvss.t1550 539.465
R13100 dvss dvss.t460 539.465
R13101 dvss.t1358 dvss.t467 539.465
R13102 dvss.t1261 dvss.t171 539.465
R13103 dvss.t1289 dvss.n4192 539.465
R13104 dvss dvss.t102 539.465
R13105 dvss dvss.t850 539.465
R13106 dvss.t1168 dvss 539.465
R13107 dvss.t2076 dvss 539.465
R13108 dvss.n3134 dvss.n3127 539.294
R13109 dvss.n3327 dvss.n3134 539.294
R13110 dvss.n3327 dvss.n3135 539.294
R13111 dvss.n3323 dvss.n3135 539.294
R13112 dvss.n3323 dvss.n3138 539.294
R13113 dvss.n3319 dvss.n3138 539.294
R13114 dvss.n3319 dvss.n3144 539.294
R13115 dvss.n3315 dvss.n3144 539.294
R13116 dvss.n3315 dvss.n3146 539.294
R13117 dvss.n3311 dvss.n3146 539.294
R13118 dvss.n3311 dvss.n3152 539.294
R13119 dvss.n3307 dvss.n3152 539.294
R13120 dvss.n3307 dvss.n3154 539.294
R13121 dvss.n3303 dvss.n3154 539.294
R13122 dvss.n3303 dvss.n3159 539.294
R13123 dvss.n3298 dvss.n3159 539.294
R13124 dvss.n3298 dvss.n3267 539.294
R13125 dvss.n3294 dvss.n3267 539.294
R13126 dvss.n3294 dvss.n3286 539.294
R13127 dvss.n3290 dvss.n3286 539.294
R13128 dvss.n1207 dvss.n1206 539.294
R13129 dvss.n5489 dvss.n1206 539.294
R13130 dvss.n5487 dvss.n5486 539.294
R13131 dvss.n5483 dvss.n5482 539.294
R13132 dvss.n5479 dvss.n5478 539.294
R13133 dvss.n5475 dvss.n5474 539.294
R13134 dvss.n5471 dvss.n5470 539.294
R13135 dvss.n5467 dvss.n5466 539.294
R13136 dvss.n5463 dvss.n5462 539.294
R13137 dvss.n5459 dvss.n5458 539.294
R13138 dvss.n5455 dvss.n5454 539.294
R13139 dvss.n5451 dvss.n5450 539.294
R13140 dvss.n5447 dvss.n5446 539.294
R13141 dvss.n5443 dvss.n5442 539.294
R13142 dvss.n5439 dvss.n5438 539.294
R13143 dvss.n5435 dvss.n5434 539.294
R13144 dvss.n5431 dvss.n5430 539.294
R13145 dvss.n5427 dvss.n5426 539.294
R13146 dvss.n5423 dvss.n5422 539.294
R13147 dvss.n5419 dvss.n5418 539.294
R13148 dvss.n5415 dvss.n5414 539.294
R13149 dvss.n5411 dvss.n5410 539.294
R13150 dvss.n5407 dvss.n5406 539.294
R13151 dvss.n5403 dvss.n5402 539.294
R13152 dvss.n5399 dvss.n5398 539.294
R13153 dvss.n5395 dvss.n5394 539.294
R13154 dvss.n5391 dvss.n5390 539.294
R13155 dvss.n5387 dvss.n5386 539.294
R13156 dvss.n5383 dvss.n5382 539.294
R13157 dvss.n5379 dvss.n5378 539.294
R13158 dvss.n5375 dvss.n5374 539.294
R13159 dvss.n5371 dvss.n5370 539.294
R13160 dvss.n5367 dvss.n5366 539.294
R13161 dvss.n5363 dvss.n5362 539.294
R13162 dvss.n5359 dvss.n5358 539.294
R13163 dvss.n5355 dvss.n5354 539.294
R13164 dvss.n5351 dvss.n5350 539.294
R13165 dvss.n5347 dvss.n5346 539.294
R13166 dvss.n5343 dvss.n5342 539.294
R13167 dvss.n5339 dvss.n5338 539.294
R13168 dvss.n5335 dvss.n5334 539.294
R13169 dvss.n5331 dvss.n5330 539.294
R13170 dvss.n5327 dvss.n5326 539.294
R13171 dvss.n5323 dvss.n5322 539.294
R13172 dvss.n5319 dvss.n5318 539.294
R13173 dvss.n5315 dvss.n5314 539.294
R13174 dvss.n5311 dvss.n5310 539.294
R13175 dvss.n5307 dvss.n5306 539.294
R13176 dvss.n5303 dvss.n5302 539.294
R13177 dvss.n5299 dvss.n5298 539.294
R13178 dvss.n5295 dvss.n5294 539.294
R13179 dvss.n5291 dvss.n5290 539.294
R13180 dvss.n5287 dvss.n1152 539.294
R13181 dvss.n5497 dvss.n1151 539.294
R13182 dvss.n5509 dvss.n1146 539.294
R13183 dvss.n5509 dvss.n1144 539.294
R13184 dvss.n5513 dvss.n1144 539.294
R13185 dvss.n5513 dvss.n1141 539.294
R13186 dvss.n5520 dvss.n1141 539.294
R13187 dvss.n5520 dvss.n1139 539.294
R13188 dvss.n5524 dvss.n1139 539.294
R13189 dvss.n5524 dvss.n1124 539.294
R13190 dvss.n5608 dvss.n1124 539.294
R13191 dvss.n5608 dvss.n1125 539.294
R13192 dvss.n5604 dvss.n1125 539.294
R13193 dvss.n5604 dvss.n1131 539.294
R13194 dvss.n5600 dvss.n1131 539.294
R13195 dvss.n5600 dvss.n1133 539.294
R13196 dvss.n5596 dvss.n1133 539.294
R13197 dvss.n5596 dvss.n5541 539.294
R13198 dvss.n5592 dvss.n5541 539.294
R13199 dvss.n5592 dvss.n5544 539.294
R13200 dvss.n5588 dvss.n5544 539.294
R13201 dvss.n5588 dvss.n5550 539.294
R13202 dvss.n5584 dvss.n5550 539.294
R13203 dvss.n5584 dvss.n5551 539.294
R13204 dvss.n5580 dvss.n5551 539.294
R13205 dvss.n5580 dvss.n5562 539.294
R13206 dvss.n5576 dvss.n5562 539.294
R13207 dvss.n5576 dvss.n5565 539.294
R13208 dvss.n5572 dvss.n5565 539.294
R13209 dvss.n5572 dvss.n523 539.294
R13210 dvss.n6210 dvss.n523 539.294
R13211 dvss.n6210 dvss.n520 539.294
R13212 dvss.n6219 dvss.n520 539.294
R13213 dvss.n6219 dvss.n518 539.294
R13214 dvss.n6225 dvss.n518 539.294
R13215 dvss.n6225 dvss.n519 539.294
R13216 dvss.n519 dvss.n508 539.294
R13217 dvss.n6237 dvss.n508 539.294
R13218 dvss.n6237 dvss.n506 539.294
R13219 dvss.n6242 dvss.n506 539.294
R13220 dvss.n6242 dvss.n503 539.294
R13221 dvss.n6249 dvss.n503 539.294
R13222 dvss.n6249 dvss.n501 539.294
R13223 dvss.n6254 dvss.n501 539.294
R13224 dvss.n6254 dvss.n497 539.294
R13225 dvss.n6265 dvss.n497 539.294
R13226 dvss.n6265 dvss.n496 539.294
R13227 dvss.n6269 dvss.n496 539.294
R13228 dvss.n6269 dvss.n493 539.294
R13229 dvss.n6276 dvss.n493 539.294
R13230 dvss.n6276 dvss.n491 539.294
R13231 dvss.n6281 dvss.n491 539.294
R13232 dvss.n6281 dvss.n488 539.294
R13233 dvss.n6290 dvss.n488 539.294
R13234 dvss.n6290 dvss.n486 539.294
R13235 dvss.n6294 dvss.n486 539.294
R13236 dvss.n6294 dvss.n478 539.294
R13237 dvss.n6307 dvss.n478 539.294
R13238 dvss.n6307 dvss.n476 539.294
R13239 dvss.n6311 dvss.n476 539.294
R13240 dvss.n6316 dvss.n6311 539.294
R13241 dvss.n6316 dvss.n6312 539.294
R13242 dvss.n6312 dvss.n473 539.294
R13243 dvss.n473 dvss.n470 539.294
R13244 dvss.n6333 dvss.n470 539.294
R13245 dvss.n6333 dvss.n467 539.294
R13246 dvss.n6337 dvss.n467 539.294
R13247 dvss.n6338 dvss.n6337 539.294
R13248 dvss.n6338 dvss.n460 539.294
R13249 dvss.n461 dvss.n460 539.294
R13250 dvss.n6342 dvss.n461 539.294
R13251 dvss.n6342 dvss.n463 539.294
R13252 dvss.n6570 dvss.n463 539.294
R13253 dvss.n6570 dvss.n466 539.294
R13254 dvss.n6566 dvss.n466 539.294
R13255 dvss.n6566 dvss.n228 539.294
R13256 dvss.n6645 dvss.n228 539.294
R13257 dvss.n6645 dvss.n229 539.294
R13258 dvss.n6641 dvss.n229 539.294
R13259 dvss.n6641 dvss.n235 539.294
R13260 dvss.n6359 dvss.n235 539.294
R13261 dvss.n6360 dvss.n6359 539.294
R13262 dvss.n6553 dvss.n6360 539.294
R13263 dvss.n6553 dvss.n6361 539.294
R13264 dvss.n6549 dvss.n6361 539.294
R13265 dvss.n6549 dvss.n6364 539.294
R13266 dvss.n6545 dvss.n6364 539.294
R13267 dvss.n6545 dvss.n6370 539.294
R13268 dvss.n6541 dvss.n6370 539.294
R13269 dvss.n6541 dvss.n6371 539.294
R13270 dvss.n6537 dvss.n6371 539.294
R13271 dvss.n6537 dvss.n6382 539.294
R13272 dvss.n6533 dvss.n6382 539.294
R13273 dvss.n6533 dvss.n6385 539.294
R13274 dvss.n6529 dvss.n6385 539.294
R13275 dvss.n6529 dvss.n6391 539.294
R13276 dvss.n6525 dvss.n6391 539.294
R13277 dvss.n6525 dvss.n6393 539.294
R13278 dvss.n6521 dvss.n6393 539.294
R13279 dvss.n6521 dvss.n6399 539.294
R13280 dvss.n6400 dvss.n6399 539.294
R13281 dvss.n6516 dvss.n6400 539.294
R13282 dvss.n6516 dvss.n6401 539.294
R13283 dvss.n6512 dvss.n6401 539.294
R13284 dvss.n6512 dvss.n6407 539.294
R13285 dvss.n6508 dvss.n6407 539.294
R13286 dvss.n6508 dvss.n6410 539.294
R13287 dvss.n6504 dvss.n6410 539.294
R13288 dvss.n1697 dvss.n1597 539.294
R13289 dvss.n1753 dvss.n1597 539.294
R13290 dvss.n1596 dvss.n1595 539.294
R13291 dvss.n1748 dvss.n1595 539.294
R13292 dvss.n1746 dvss.n1745 539.294
R13293 dvss.n1742 dvss.n1741 539.294
R13294 dvss.n1738 dvss.n1737 539.294
R13295 dvss.n1756 dvss.n1568 539.294
R13296 dvss.n1756 dvss.n1569 539.294
R13297 dvss.n1581 dvss.n1569 539.294
R13298 dvss.n1590 dvss.n1579 539.294
R13299 dvss.n1591 dvss.n1551 539.294
R13300 dvss.n1791 dvss.n1551 539.294
R13301 dvss.n1791 dvss.n1548 539.294
R13302 dvss.n1798 dvss.n1548 539.294
R13303 dvss.n1798 dvss.n1541 539.294
R13304 dvss.n1813 dvss.n1541 539.294
R13305 dvss.n1813 dvss.n1537 539.294
R13306 dvss.n1821 dvss.n1537 539.294
R13307 dvss.n1821 dvss.n1531 539.294
R13308 dvss.n1833 dvss.n1531 539.294
R13309 dvss.n1833 dvss.n1526 539.294
R13310 dvss.n1847 dvss.n1526 539.294
R13311 dvss.n1847 dvss.n1522 539.294
R13312 dvss.n1854 dvss.n1522 539.294
R13313 dvss.n1854 dvss.n1523 539.294
R13314 dvss.n1523 dvss.n1511 539.294
R13315 dvss.n1511 dvss.n1504 539.294
R13316 dvss.n1875 dvss.n1504 539.294
R13317 dvss.n1876 dvss.n1875 539.294
R13318 dvss.n1880 dvss.n1498 539.294
R13319 dvss.n1501 dvss.n1499 539.294
R13320 dvss.n1501 dvss.n1484 539.294
R13321 dvss.n1903 dvss.n1484 539.294
R13322 dvss.n1903 dvss.n1480 539.294
R13323 dvss.n1916 dvss.n1480 539.294
R13324 dvss.n1916 dvss.n1472 539.294
R13325 dvss.n1932 dvss.n1472 539.294
R13326 dvss.n1933 dvss.n1932 539.294
R13327 dvss.n1933 dvss.n1458 539.294
R13328 dvss.n1983 dvss.n1458 539.294
R13329 dvss.n1983 dvss.n1459 539.294
R13330 dvss.n1952 dvss.n1459 539.294
R13331 dvss.n1959 dvss.n1952 539.294
R13332 dvss.n1960 dvss.n1959 539.294
R13333 dvss.n1960 dvss.n1455 539.294
R13334 dvss.n2019 dvss.n1455 539.294
R13335 dvss.n2019 dvss.n1442 539.294
R13336 dvss.n2054 dvss.n1442 539.294
R13337 dvss.n2054 dvss.n1443 539.294
R13338 dvss.n2034 dvss.n2031 539.294
R13339 dvss.n2032 dvss.n1434 539.294
R13340 dvss.n1434 dvss.n1430 539.294
R13341 dvss.n2070 dvss.n1430 539.294
R13342 dvss.n2071 dvss.n2070 539.294
R13343 dvss.n2071 dvss.n1420 539.294
R13344 dvss.n2084 dvss.n1420 539.294
R13345 dvss.n2085 dvss.n2084 539.294
R13346 dvss.n2085 dvss.n1351 539.294
R13347 dvss.n2103 dvss.n1351 539.294
R13348 dvss.n2103 dvss.n1352 539.294
R13349 dvss.n1378 dvss.n1352 539.294
R13350 dvss.n1382 dvss.n1378 539.294
R13351 dvss.n1382 dvss.n1365 539.294
R13352 dvss.n1394 dvss.n1365 539.294
R13353 dvss.n1395 dvss.n1394 539.294
R13354 dvss.n1395 dvss.n891 539.294
R13355 dvss.n5729 dvss.n891 539.294
R13356 dvss.n5729 dvss.n892 539.294
R13357 dvss.n1004 dvss.n892 539.294
R13358 dvss.n1003 dvss.n1002 539.294
R13359 dvss.n1000 dvss.n999 539.294
R13360 dvss.n1017 dvss.n999 539.294
R13361 dvss.n1018 dvss.n1017 539.294
R13362 dvss.n1018 dvss.n993 539.294
R13363 dvss.n1024 dvss.n993 539.294
R13364 dvss.n1026 dvss.n1024 539.294
R13365 dvss.n1026 dvss.n1025 539.294
R13366 dvss.n1025 dvss.n990 539.294
R13367 dvss.n1034 dvss.n990 539.294
R13368 dvss.n1036 dvss.n1034 539.294
R13369 dvss.n1037 dvss.n1036 539.294
R13370 dvss.n1038 dvss.n1037 539.294
R13371 dvss.n1038 dvss.n978 539.294
R13372 dvss.n1046 dvss.n978 539.294
R13373 dvss.n1046 dvss.n974 539.294
R13374 dvss.n1052 dvss.n974 539.294
R13375 dvss.n1053 dvss.n1052 539.294
R13376 dvss.n1056 dvss.n1053 539.294
R13377 dvss.n1057 dvss.n1056 539.294
R13378 dvss.n973 dvss.n970 539.294
R13379 dvss.n1061 dvss.n966 539.294
R13380 dvss.n5660 dvss.n966 539.294
R13381 dvss.n5660 dvss.n967 539.294
R13382 dvss.n5656 dvss.n967 539.294
R13383 dvss.n5656 dvss.n1067 539.294
R13384 dvss.n5652 dvss.n1067 539.294
R13385 dvss.n5652 dvss.n1072 539.294
R13386 dvss.n1075 dvss.n1072 539.294
R13387 dvss.n1113 dvss.n1075 539.294
R13388 dvss.n5613 dvss.n1113 539.294
R13389 dvss.n5614 dvss.n5613 539.294
R13390 dvss.n5614 dvss.n1111 539.294
R13391 dvss.n5619 dvss.n1111 539.294
R13392 dvss.n5620 dvss.n5619 539.294
R13393 dvss.n5620 dvss.n805 539.294
R13394 dvss.n6122 dvss.n805 539.294
R13395 dvss.n6122 dvss.n792 539.294
R13396 dvss.n6157 dvss.n792 539.294
R13397 dvss.n6157 dvss.n793 539.294
R13398 dvss.n6137 dvss.n6134 539.294
R13399 dvss.n6135 dvss.n784 539.294
R13400 dvss.n784 dvss.n780 539.294
R13401 dvss.n6173 dvss.n780 539.294
R13402 dvss.n6174 dvss.n6173 539.294
R13403 dvss.n6174 dvss.n770 539.294
R13404 dvss.n6187 dvss.n770 539.294
R13405 dvss.n6188 dvss.n6187 539.294
R13406 dvss.n6188 dvss.n528 539.294
R13407 dvss.n6206 dvss.n528 539.294
R13408 dvss.n6206 dvss.n529 539.294
R13409 dvss.n628 dvss.n529 539.294
R13410 dvss.n634 dvss.n628 539.294
R13411 dvss.n634 dvss.n614 539.294
R13412 dvss.n646 dvss.n614 539.294
R13413 dvss.n646 dvss.n610 539.294
R13414 dvss.n652 dvss.n610 539.294
R13415 dvss.n653 dvss.n652 539.294
R13416 dvss.n660 dvss.n653 539.294
R13417 dvss.n660 dvss.n659 539.294
R13418 dvss.n657 dvss.n656 539.294
R13419 dvss.n654 dvss.n607 539.294
R13420 dvss.n672 dvss.n607 539.294
R13421 dvss.n673 dvss.n672 539.294
R13422 dvss.n673 dvss.n601 539.294
R13423 dvss.n679 dvss.n601 539.294
R13424 dvss.n681 dvss.n679 539.294
R13425 dvss.n681 dvss.n680 539.294
R13426 dvss.n680 dvss.n598 539.294
R13427 dvss.n689 dvss.n598 539.294
R13428 dvss.n691 dvss.n689 539.294
R13429 dvss.n692 dvss.n691 539.294
R13430 dvss.n693 dvss.n692 539.294
R13431 dvss.n693 dvss.n593 539.294
R13432 dvss.n700 dvss.n593 539.294
R13433 dvss.n701 dvss.n700 539.294
R13434 dvss.n701 dvss.n125 539.294
R13435 dvss.n6713 dvss.n125 539.294
R13436 dvss.n6713 dvss.n126 539.294
R13437 dvss.n199 dvss.n126 539.294
R13438 dvss.n198 dvss.n197 539.294
R13439 dvss.n205 dvss.n203 539.294
R13440 dvss.n205 dvss.n188 539.294
R13441 dvss.n209 dvss.n188 539.294
R13442 dvss.n210 dvss.n209 539.294
R13443 dvss.n215 dvss.n210 539.294
R13444 dvss.n215 dvss.n184 539.294
R13445 dvss.n220 dvss.n184 539.294
R13446 dvss.n221 dvss.n220 539.294
R13447 dvss.n221 dvss.n182 539.294
R13448 dvss.n6649 dvss.n182 539.294
R13449 dvss.n6650 dvss.n6649 539.294
R13450 dvss.n6650 dvss.n179 539.294
R13451 dvss.n6656 dvss.n179 539.294
R13452 dvss.n6657 dvss.n6656 539.294
R13453 dvss.n6657 dvss.n76 539.294
R13454 dvss.n6863 dvss.n76 539.294
R13455 dvss.n6863 dvss.n68 539.294
R13456 dvss.n6898 dvss.n68 539.294
R13457 dvss.n6898 dvss.n69 539.294
R13458 dvss.n6878 dvss.n6875 539.294
R13459 dvss.n6876 dvss.n60 539.294
R13460 dvss.n60 dvss.n56 539.294
R13461 dvss.n6914 dvss.n56 539.294
R13462 dvss.n6915 dvss.n6914 539.294
R13463 dvss.n6915 dvss.n46 539.294
R13464 dvss.n6928 dvss.n46 539.294
R13465 dvss.n6929 dvss.n6928 539.294
R13466 dvss.n6929 dvss.n26 539.294
R13467 dvss.n6947 dvss.n26 539.294
R13468 dvss.n6947 dvss.n27 539.294
R13469 dvss.n6458 dvss.n27 539.294
R13470 dvss.n6458 dvss.n6446 539.294
R13471 dvss.n6470 dvss.n6446 539.294
R13472 dvss.n6470 dvss.n6442 539.294
R13473 dvss.n6478 dvss.n6442 539.294
R13474 dvss.n6478 dvss.n6438 539.294
R13475 dvss.n6489 dvss.n6438 539.294
R13476 dvss.n6490 dvss.n6489 539.294
R13477 dvss.n6490 dvss.n6434 539.294
R13478 dvss.n6434 dvss.n6430 539.294
R13479 dvss.n3198 dvss.n3194 539.294
R13480 dvss.n3205 dvss.n3194 539.294
R13481 dvss.n3205 dvss.n3192 539.294
R13482 dvss.n3209 dvss.n3192 539.294
R13483 dvss.n3209 dvss.n3186 539.294
R13484 dvss.n3220 dvss.n3186 539.294
R13485 dvss.n3220 dvss.n3184 539.294
R13486 dvss.n3225 dvss.n3184 539.294
R13487 dvss.n3225 dvss.n3176 539.294
R13488 dvss.n3235 dvss.n3176 539.294
R13489 dvss.n3235 dvss.n3175 539.294
R13490 dvss.n3241 dvss.n3175 539.294
R13491 dvss.n3241 dvss.n3168 539.294
R13492 dvss.n3251 dvss.n3168 539.294
R13493 dvss.n3251 dvss.n3167 539.294
R13494 dvss.n3255 dvss.n3167 539.294
R13495 dvss.n3255 dvss.n3162 539.294
R13496 dvss.n3263 dvss.n3162 539.294
R13497 dvss.n3263 dvss.n3163 539.294
R13498 dvss.n3163 dvss.n239 539.294
R13499 dvss.n6636 dvss.n239 539.294
R13500 dvss.n1694 dvss.n1690 539.294
R13501 dvss.n1728 dvss.n1690 539.294
R13502 dvss.n1689 dvss.n1688 539.294
R13503 dvss.n1723 dvss.n1688 539.294
R13504 dvss.n1721 dvss.n1720 539.294
R13505 dvss.n1717 dvss.n1716 539.294
R13506 dvss.n1732 dvss.n1623 539.294
R13507 dvss.n1624 dvss.n1560 539.294
R13508 dvss.n1770 dvss.n1560 539.294
R13509 dvss.n1559 dvss.n1558 539.294
R13510 dvss.n1774 dvss.n1549 539.294
R13511 dvss.n1793 dvss.n1549 539.294
R13512 dvss.n1794 dvss.n1793 539.294
R13513 dvss.n1794 dvss.n1546 539.294
R13514 dvss.n1546 dvss.n1539 539.294
R13515 dvss.n1815 dvss.n1539 539.294
R13516 dvss.n1816 dvss.n1815 539.294
R13517 dvss.n1816 dvss.n1535 539.294
R13518 dvss.n1535 dvss.n1529 539.294
R13519 dvss.n1835 dvss.n1529 539.294
R13520 dvss.n1836 dvss.n1835 539.294
R13521 dvss.n1836 dvss.n1525 539.294
R13522 dvss.n1525 dvss.n1519 539.294
R13523 dvss.n1520 dvss.n1519 539.294
R13524 dvss.n1850 dvss.n1520 539.294
R13525 dvss.n1850 dvss.n1507 539.294
R13526 dvss.n1872 dvss.n1507 539.294
R13527 dvss.n1872 dvss.n1493 539.294
R13528 dvss.n1886 dvss.n1493 539.294
R13529 dvss.n1492 dvss.n1490 539.294
R13530 dvss.n1890 dvss.n1485 539.294
R13531 dvss.n1900 dvss.n1485 539.294
R13532 dvss.n1900 dvss.n1481 539.294
R13533 dvss.n1913 dvss.n1481 539.294
R13534 dvss.n1913 dvss.n1474 539.294
R13535 dvss.n1928 dvss.n1474 539.294
R13536 dvss.n1928 dvss.n1468 539.294
R13537 dvss.n1935 dvss.n1468 539.294
R13538 dvss.n1935 dvss.n1470 539.294
R13539 dvss.n1470 dvss.n1457 539.294
R13540 dvss.n1463 dvss.n1457 539.294
R13541 dvss.n1956 dvss.n1463 539.294
R13542 dvss.n1957 dvss.n1956 539.294
R13543 dvss.n1957 dvss.n1951 539.294
R13544 dvss.n1963 dvss.n1951 539.294
R13545 dvss.n1963 dvss.n1456 539.294
R13546 dvss.n1456 dvss.n1447 539.294
R13547 dvss.n1447 dvss.n1441 539.294
R13548 dvss.n2027 dvss.n1441 539.294
R13549 dvss.n2045 dvss.n2041 539.294
R13550 dvss.n2059 dvss.n1437 539.294
R13551 dvss.n2059 dvss.n1431 539.294
R13552 dvss.n2068 dvss.n1431 539.294
R13553 dvss.n2068 dvss.n1423 539.294
R13554 dvss.n2081 dvss.n1423 539.294
R13555 dvss.n2081 dvss.n1415 539.294
R13556 dvss.n2087 dvss.n1415 539.294
R13557 dvss.n2087 dvss.n1416 539.294
R13558 dvss.n1416 dvss.n1350 539.294
R13559 dvss.n1357 dvss.n1350 539.294
R13560 dvss.n1379 dvss.n1357 539.294
R13561 dvss.n1379 dvss.n1367 539.294
R13562 dvss.n1391 dvss.n1367 539.294
R13563 dvss.n1391 dvss.n1363 539.294
R13564 dvss.n1397 dvss.n1363 539.294
R13565 dvss.n1397 dvss.n1364 539.294
R13566 dvss.n1364 dvss.n889 539.294
R13567 dvss.n897 dvss.n889 539.294
R13568 dvss.n1009 dvss.n897 539.294
R13569 dvss.n902 dvss.n901 539.294
R13570 dvss.n1014 dvss.n1013 539.294
R13571 dvss.n1014 dvss.n911 539.294
R13572 dvss.n912 dvss.n911 539.294
R13573 dvss.n1021 dvss.n912 539.294
R13574 dvss.n1022 dvss.n1021 539.294
R13575 dvss.n1022 dvss.n922 539.294
R13576 dvss.n923 dvss.n922 539.294
R13577 dvss.n1031 dvss.n923 539.294
R13578 dvss.n1032 dvss.n1031 539.294
R13579 dvss.n1032 dvss.n931 539.294
R13580 dvss.n932 dvss.n931 539.294
R13581 dvss.n988 dvss.n932 539.294
R13582 dvss.n1041 dvss.n988 539.294
R13583 dvss.n1041 dvss.n976 539.294
R13584 dvss.n1049 dvss.n976 539.294
R13585 dvss.n1050 dvss.n1049 539.294
R13586 dvss.n1050 dvss.n946 539.294
R13587 dvss.n947 dvss.n946 539.294
R13588 dvss.n5669 dvss.n947 539.294
R13589 dvss.n5671 dvss.n952 539.294
R13590 dvss.n5666 dvss.n954 539.294
R13591 dvss.n5662 dvss.n954 539.294
R13592 dvss.n5662 dvss.n965 539.294
R13593 dvss.n1069 dvss.n965 539.294
R13594 dvss.n1070 dvss.n1069 539.294
R13595 dvss.n1071 dvss.n1070 539.294
R13596 dvss.n1116 dvss.n1071 539.294
R13597 dvss.n1116 dvss.n1078 539.294
R13598 dvss.n1079 dvss.n1078 539.294
R13599 dvss.n5611 dvss.n1079 539.294
R13600 dvss.n5611 dvss.n1102 539.294
R13601 dvss.n1103 dvss.n1102 539.294
R13602 dvss.n5617 dvss.n1103 539.294
R13603 dvss.n5617 dvss.n1110 539.294
R13604 dvss.n5623 dvss.n1110 539.294
R13605 dvss.n5623 dvss.n806 539.294
R13606 dvss.n806 dvss.n797 539.294
R13607 dvss.n797 dvss.n791 539.294
R13608 dvss.n6130 dvss.n791 539.294
R13609 dvss.n6148 dvss.n6144 539.294
R13610 dvss.n6162 dvss.n787 539.294
R13611 dvss.n6162 dvss.n781 539.294
R13612 dvss.n6171 dvss.n781 539.294
R13613 dvss.n6171 dvss.n773 539.294
R13614 dvss.n6184 dvss.n773 539.294
R13615 dvss.n6184 dvss.n765 539.294
R13616 dvss.n6190 dvss.n765 539.294
R13617 dvss.n6190 dvss.n766 539.294
R13618 dvss.n766 dvss.n527 539.294
R13619 dvss.n534 dvss.n527 539.294
R13620 dvss.n630 dvss.n534 539.294
R13621 dvss.n631 dvss.n630 539.294
R13622 dvss.n631 dvss.n620 539.294
R13623 dvss.n620 dvss.n612 539.294
R13624 dvss.n649 dvss.n612 539.294
R13625 dvss.n650 dvss.n649 539.294
R13626 dvss.n650 dvss.n541 539.294
R13627 dvss.n542 dvss.n541 539.294
R13628 dvss.n664 dvss.n542 539.294
R13629 dvss.n548 dvss.n547 539.294
R13630 dvss.n669 dvss.n668 539.294
R13631 dvss.n669 dvss.n557 539.294
R13632 dvss.n558 dvss.n557 539.294
R13633 dvss.n676 dvss.n558 539.294
R13634 dvss.n677 dvss.n676 539.294
R13635 dvss.n677 dvss.n568 539.294
R13636 dvss.n569 dvss.n568 539.294
R13637 dvss.n686 dvss.n569 539.294
R13638 dvss.n687 dvss.n686 539.294
R13639 dvss.n687 dvss.n577 539.294
R13640 dvss.n578 dvss.n577 539.294
R13641 dvss.n695 dvss.n578 539.294
R13642 dvss.n697 dvss.n695 539.294
R13643 dvss.n697 dvss.n591 539.294
R13644 dvss.n703 dvss.n591 539.294
R13645 dvss.n703 dvss.n592 539.294
R13646 dvss.n592 dvss.n123 539.294
R13647 dvss.n131 dvss.n123 539.294
R13648 dvss.n191 dvss.n131 539.294
R13649 dvss.n136 dvss.n135 539.294
R13650 dvss.n196 dvss.n195 539.294
R13651 dvss.n196 dvss.n145 539.294
R13652 dvss.n146 dvss.n145 539.294
R13653 dvss.n186 dvss.n146 539.294
R13654 dvss.n187 dvss.n186 539.294
R13655 dvss.n187 dvss.n156 539.294
R13656 dvss.n157 dvss.n156 539.294
R13657 dvss.n223 dvss.n157 539.294
R13658 dvss.n224 dvss.n223 539.294
R13659 dvss.n224 dvss.n165 539.294
R13660 dvss.n166 dvss.n165 539.294
R13661 dvss.n6653 dvss.n166 539.294
R13662 dvss.n6654 dvss.n6653 539.294
R13663 dvss.n6654 dvss.n178 539.294
R13664 dvss.n6660 dvss.n178 539.294
R13665 dvss.n6660 dvss.n77 539.294
R13666 dvss.n77 dvss.n73 539.294
R13667 dvss.n73 dvss.n67 539.294
R13668 dvss.n6871 dvss.n67 539.294
R13669 dvss.n6889 dvss.n6885 539.294
R13670 dvss.n6903 dvss.n63 539.294
R13671 dvss.n6903 dvss.n57 539.294
R13672 dvss.n6912 dvss.n57 539.294
R13673 dvss.n6912 dvss.n49 539.294
R13674 dvss.n6925 dvss.n49 539.294
R13675 dvss.n6925 dvss.n41 539.294
R13676 dvss.n6931 dvss.n41 539.294
R13677 dvss.n6931 dvss.n42 539.294
R13678 dvss.n42 dvss.n25 539.294
R13679 dvss.n32 dvss.n25 539.294
R13680 dvss.n6455 dvss.n32 539.294
R13681 dvss.n6461 dvss.n6455 539.294
R13682 dvss.n6461 dvss.n6445 539.294
R13683 dvss.n6473 dvss.n6445 539.294
R13684 dvss.n6473 dvss.n6441 539.294
R13685 dvss.n6481 dvss.n6441 539.294
R13686 dvss.n6481 dvss.n6436 539.294
R13687 dvss.n6492 dvss.n6436 539.294
R13688 dvss.n6492 dvss.n6431 539.294
R13689 dvss.n6500 dvss.n6431 539.294
R13690 dvss.n2293 dvss.n1 539.294
R13691 dvss.n2 dvss.n1 539.294
R13692 dvss.n2289 dvss.n2 539.294
R13693 dvss.n2289 dvss.n2288 539.294
R13694 dvss.n2288 dvss.n1241 539.294
R13695 dvss.n1243 dvss.n1241 539.294
R13696 dvss.n1244 dvss.n1243 539.294
R13697 dvss.n1684 dvss.n1244 539.294
R13698 dvss.n1684 dvss.n1247 539.294
R13699 dvss.n1248 dvss.n1247 539.294
R13700 dvss.n1680 dvss.n1248 539.294
R13701 dvss.n1680 dvss.n1252 539.294
R13702 dvss.n1253 dvss.n1252 539.294
R13703 dvss.n1676 dvss.n1253 539.294
R13704 dvss.n1676 dvss.n1257 539.294
R13705 dvss.n1258 dvss.n1257 539.294
R13706 dvss.n1672 dvss.n1260 539.294
R13707 dvss.n1261 dvss.n1260 539.294
R13708 dvss.n1668 dvss.n1261 539.294
R13709 dvss.n1668 dvss.n1667 539.294
R13710 dvss.n1667 dvss.n1266 539.294
R13711 dvss.n1267 dvss.n1266 539.294
R13712 dvss.n1633 dvss.n1267 539.294
R13713 dvss.n1633 dvss.n1272 539.294
R13714 dvss.n1273 dvss.n1272 539.294
R13715 dvss.n1663 dvss.n1273 539.294
R13716 dvss.n1663 dvss.n1276 539.294
R13717 dvss.n1277 dvss.n1276 539.294
R13718 dvss.n1659 dvss.n1277 539.294
R13719 dvss.n1659 dvss.n1658 539.294
R13720 dvss.n1658 dvss.n1283 539.294
R13721 dvss.n1284 dvss.n1283 539.294
R13722 dvss.n1653 dvss.n1284 539.294
R13723 dvss.n1653 dvss.n1286 539.294
R13724 dvss.n1287 dvss.n1286 539.294
R13725 dvss.n1646 dvss.n1287 539.294
R13726 dvss.n1290 dvss.n1289 539.294
R13727 dvss.n1644 dvss.n1292 539.294
R13728 dvss.n1293 dvss.n1292 539.294
R13729 dvss.n1640 dvss.n1293 539.294
R13730 dvss.n1640 dvss.n1297 539.294
R13731 dvss.n1298 dvss.n1297 539.294
R13732 dvss.n1636 dvss.n1298 539.294
R13733 dvss.n1636 dvss.n1303 539.294
R13734 dvss.n1304 dvss.n1303 539.294
R13735 dvss.n1988 dvss.n1304 539.294
R13736 dvss.n1988 dvss.n1307 539.294
R13737 dvss.n1308 dvss.n1307 539.294
R13738 dvss.n1993 dvss.n1308 539.294
R13739 dvss.n1994 dvss.n1993 539.294
R13740 dvss.n1994 dvss.n1314 539.294
R13741 dvss.n1315 dvss.n1314 539.294
R13742 dvss.n1998 dvss.n1315 539.294
R13743 dvss.n1998 dvss.n1317 539.294
R13744 dvss.n1318 dvss.n1317 539.294
R13745 dvss.n2002 dvss.n1318 539.294
R13746 dvss.n1321 dvss.n1320 539.294
R13747 dvss.n2000 dvss.n1323 539.294
R13748 dvss.n1324 dvss.n1323 539.294
R13749 dvss.n2009 dvss.n1324 539.294
R13750 dvss.n2009 dvss.n1328 539.294
R13751 dvss.n1329 dvss.n1328 539.294
R13752 dvss.n2007 dvss.n1329 539.294
R13753 dvss.n2007 dvss.n1334 539.294
R13754 dvss.n1335 dvss.n1334 539.294
R13755 dvss.n2106 dvss.n1335 539.294
R13756 dvss.n2106 dvss.n1338 539.294
R13757 dvss.n1339 dvss.n1338 539.294
R13758 dvss.n2110 dvss.n1339 539.294
R13759 dvss.n2110 dvss.n1346 539.294
R13760 dvss.n2114 dvss.n1346 539.294
R13761 dvss.n2114 dvss.n886 539.294
R13762 dvss.n5734 dvss.n886 539.294
R13763 dvss.n5734 dvss.n876 539.294
R13764 dvss.n5750 dvss.n876 539.294
R13765 dvss.n5750 dvss.n877 539.294
R13766 dvss.n5741 dvss.n5739 539.294
R13767 dvss.n5755 dvss.n873 539.294
R13768 dvss.n5755 dvss.n869 539.294
R13769 dvss.n5766 dvss.n869 539.294
R13770 dvss.n5766 dvss.n867 539.294
R13771 dvss.n5770 dvss.n867 539.294
R13772 dvss.n5770 dvss.n863 539.294
R13773 dvss.n5784 dvss.n863 539.294
R13774 dvss.n5784 dvss.n861 539.294
R13775 dvss.n5788 dvss.n861 539.294
R13776 dvss.n5788 dvss.n858 539.294
R13777 dvss.n5798 dvss.n858 539.294
R13778 dvss.n5798 dvss.n856 539.294
R13779 dvss.n5802 dvss.n856 539.294
R13780 dvss.n5802 dvss.n851 539.294
R13781 dvss.n5819 dvss.n851 539.294
R13782 dvss.n5819 dvss.n848 539.294
R13783 dvss.n5825 dvss.n848 539.294
R13784 dvss.n5825 dvss.n845 539.294
R13785 dvss.n5832 dvss.n845 539.294
R13786 dvss.n5836 dvss.n844 539.294
R13787 dvss.n5844 dvss.n841 539.294
R13788 dvss.n5844 dvss.n839 539.294
R13789 dvss.n5848 dvss.n839 539.294
R13790 dvss.n5848 dvss.n833 539.294
R13791 dvss.n5859 dvss.n833 539.294
R13792 dvss.n5859 dvss.n831 539.294
R13793 dvss.n5864 dvss.n831 539.294
R13794 dvss.n5864 dvss.n823 539.294
R13795 dvss.n5874 dvss.n823 539.294
R13796 dvss.n5874 dvss.n822 539.294
R13797 dvss.n5879 dvss.n822 539.294
R13798 dvss.n5879 dvss.n815 539.294
R13799 dvss.n5889 dvss.n815 539.294
R13800 dvss.n5889 dvss.n814 539.294
R13801 dvss.n5893 dvss.n814 539.294
R13802 dvss.n5893 dvss.n809 539.294
R13803 dvss.n6117 dvss.n809 539.294
R13804 dvss.n6117 dvss.n810 539.294
R13805 dvss.n5902 dvss.n810 539.294
R13806 dvss.n5919 dvss.n5903 539.294
R13807 dvss.n5906 dvss.n5905 539.294
R13808 dvss.n5926 dvss.n5906 539.294
R13809 dvss.n5927 dvss.n5926 539.294
R13810 dvss.n5927 dvss.n5911 539.294
R13811 dvss.n5912 dvss.n5911 539.294
R13812 dvss.n5918 dvss.n5912 539.294
R13813 dvss.n5918 dvss.n5917 539.294
R13814 dvss.n5934 dvss.n5917 539.294
R13815 dvss.n5977 dvss.n5934 539.294
R13816 dvss.n5977 dvss.n5937 539.294
R13817 dvss.n5938 dvss.n5937 539.294
R13818 dvss.n5982 dvss.n5938 539.294
R13819 dvss.n5983 dvss.n5982 539.294
R13820 dvss.n5983 dvss.n5944 539.294
R13821 dvss.n5945 dvss.n5944 539.294
R13822 dvss.n5987 dvss.n5945 539.294
R13823 dvss.n5987 dvss.n5947 539.294
R13824 dvss.n5948 dvss.n5947 539.294
R13825 dvss.n5994 dvss.n5948 539.294
R13826 dvss.n5951 dvss.n5950 539.294
R13827 dvss.n5992 dvss.n5953 539.294
R13828 dvss.n5954 dvss.n5953 539.294
R13829 dvss.n6000 dvss.n5954 539.294
R13830 dvss.n6000 dvss.n5958 539.294
R13831 dvss.n5959 dvss.n5958 539.294
R13832 dvss.n5976 dvss.n5959 539.294
R13833 dvss.n5976 dvss.n5964 539.294
R13834 dvss.n5965 dvss.n5964 539.294
R13835 dvss.n6007 dvss.n5965 539.294
R13836 dvss.n6007 dvss.n5968 539.294
R13837 dvss.n5969 dvss.n5968 539.294
R13838 dvss.n6012 dvss.n5969 539.294
R13839 dvss.n6013 dvss.n6012 539.294
R13840 dvss.n6013 dvss.n5975 539.294
R13841 dvss.n6017 dvss.n5975 539.294
R13842 dvss.n6017 dvss.n119 539.294
R13843 dvss.n6719 dvss.n119 539.294
R13844 dvss.n6719 dvss.n116 539.294
R13845 dvss.n6726 dvss.n116 539.294
R13846 dvss.n6730 dvss.n115 539.294
R13847 dvss.n6738 dvss.n112 539.294
R13848 dvss.n6738 dvss.n110 539.294
R13849 dvss.n6742 dvss.n110 539.294
R13850 dvss.n6742 dvss.n104 539.294
R13851 dvss.n6753 dvss.n104 539.294
R13852 dvss.n6753 dvss.n102 539.294
R13853 dvss.n6758 dvss.n102 539.294
R13854 dvss.n6758 dvss.n94 539.294
R13855 dvss.n6768 dvss.n94 539.294
R13856 dvss.n6768 dvss.n93 539.294
R13857 dvss.n6773 dvss.n93 539.294
R13858 dvss.n6773 dvss.n86 539.294
R13859 dvss.n6783 dvss.n86 539.294
R13860 dvss.n6783 dvss.n85 539.294
R13861 dvss.n6787 dvss.n85 539.294
R13862 dvss.n6787 dvss.n80 539.294
R13863 dvss.n6858 dvss.n80 539.294
R13864 dvss.n6858 dvss.n81 539.294
R13865 dvss.n6791 dvss.n81 539.294
R13866 dvss.n6807 dvss.n6792 539.294
R13867 dvss.n6795 dvss.n6794 539.294
R13868 dvss.n6814 dvss.n6795 539.294
R13869 dvss.n6815 dvss.n6814 539.294
R13870 dvss.n6815 dvss.n6800 539.294
R13871 dvss.n6801 dvss.n6800 539.294
R13872 dvss.n6819 dvss.n6801 539.294
R13873 dvss.n6821 dvss.n6819 539.294
R13874 dvss.n6822 dvss.n6821 539.294
R13875 dvss.n6822 dvss.n22 539.294
R13876 dvss.n6952 dvss.n22 539.294
R13877 dvss.n6952 dvss.n19 539.294
R13878 dvss.n6966 dvss.n19 539.294
R13879 dvss.n6966 dvss.n17 539.294
R13880 dvss.n6970 dvss.n17 539.294
R13881 dvss.n6970 dvss.n13 539.294
R13882 dvss.n6979 dvss.n13 539.294
R13883 dvss.n6979 dvss.n9 539.294
R13884 dvss.n6984 dvss.n9 539.294
R13885 dvss.n6985 dvss.n6984 539.294
R13886 dvss.n1558 dvss.n1556 533.678
R13887 dvss.n1672 dvss.n1258 533.678
R13888 dvss dvss.t1881 531.034
R13889 dvss dvss.t1754 531.034
R13890 dvss.t420 dvss.t1996 531.034
R13891 dvss dvss.t2010 531.034
R13892 dvss dvss.t598 531.034
R13893 dvss.t2004 dvss 531.034
R13894 dvss dvss.t1841 531.034
R13895 dvss dvss.t1773 531.034
R13896 dvss dvss.t1907 531.034
R13897 dvss.t1891 dvss 531.034
R13898 dvss.t634 dvss 531.034
R13899 dvss.t2032 dvss.t2042 522.606
R13900 dvss.t2080 dvss 522.606
R13901 dvss.t2183 dvss 522.606
R13902 dvss.t1528 dvss.t85 522.606
R13903 dvss.t2040 dvss 522.606
R13904 dvss dvss.t1570 514.177
R13905 dvss dvss.t2046 514.177
R13906 dvss.t565 dvss 514.177
R13907 dvss.t97 dvss.t565 514.177
R13908 dvss dvss.t872 514.177
R13909 dvss dvss.t156 514.177
R13910 dvss dvss.t846 514.177
R13911 dvss.t1422 dvss.t1435 514.177
R13912 dvss.t207 dvss.t502 514.177
R13913 dvss.t473 dvss 514.177
R13914 dvss dvss.t543 514.177
R13915 dvss.n1594 dvss.n1593 510.284
R13916 dvss.t434 dvss.t713 505.748
R13917 dvss.t877 dvss.t567 505.748
R13918 dvss.t1328 dvss 505.748
R13919 dvss.t148 dvss.t1979 505.748
R13920 dvss.t477 dvss.t1433 505.748
R13921 dvss dvss.t1332 505.748
R13922 dvss.t1527 dvss 505.748
R13923 dvss.t1235 dvss 505.748
R13924 dvss.t2070 dvss.t187 505.748
R13925 dvss.t82 dvss.t1350 505.748
R13926 dvss.n6313 dvss.n469 498.113
R13927 dvss.n6334 dvss.n469 498.113
R13928 dvss.n6336 dvss.n6335 498.113
R13929 dvss.n6340 dvss.n6339 498.113
R13930 dvss.n6341 dvss.n6340 498.113
R13931 dvss.n6343 dvss.n6341 498.113
R13932 dvss.n6344 dvss.n6343 498.113
R13933 dvss.n6250 dvss.n502 498.113
R13934 dvss.n6251 dvss.n6250 498.113
R13935 dvss.n6253 dvss.n6252 498.113
R13936 dvss.n6267 dvss.n6266 498.113
R13937 dvss.n6268 dvss.n6267 498.113
R13938 dvss.n6268 dvss.n492 498.113
R13939 dvss.n6277 dvss.n492 498.113
R13940 dvss.n6278 dvss.n6277 498.113
R13941 dvss.t526 dvss.t624 497.318
R13942 dvss.t1171 dvss.t581 497.318
R13943 dvss dvss.t698 497.318
R13944 dvss.t195 dvss.t1286 497.318
R13945 dvss.n6569 dvss.n6344 493.485
R13946 dvss.n6501 dvss.n6429 491.163
R13947 dvss.t557 dvss.t992 488.889
R13948 dvss.t1394 dvss.t146 488.889
R13949 dvss dvss.t1191 488.889
R13950 dvss dvss.t547 488.889
R13951 dvss.t319 dvss.t1241 488.889
R13952 dvss.n1695 dvss.n1693 486.048
R13953 dvss.t995 dvss.t559 480.461
R13954 dvss.t1577 dvss 480.461
R13955 dvss.t85 dvss.t915 480.461
R13956 dvss.n6638 dvss.n6637 479.541
R13957 dvss.t322 dvss.t93 472.031
R13958 dvss.n3906 dvss.t744 472.031
R13959 dvss.t883 dvss.t118 472.031
R13960 dvss dvss.t404 472.031
R13961 dvss.t2136 dvss.t377 472.031
R13962 dvss.t1051 dvss 472.031
R13963 dvss.t504 dvss.t422 472.031
R13964 dvss.t1426 dvss.t506 472.031
R13965 dvss.t142 dvss.t1548 463.603
R13966 dvss.t2094 dvss.t1838 463.603
R13967 dvss.t370 dvss.t2171 463.603
R13968 dvss dvss.t1400 455.173
R13969 dvss.t599 dvss 455.173
R13970 dvss.t2030 dvss.t1918 455.173
R13971 dvss dvss.t950 455.173
R13972 dvss.t854 dvss.t104 455.173
R13973 dvss.n4854 dvss.n1232 451.765
R13974 dvss.n4854 dvss.n4853 451.765
R13975 dvss.n4853 dvss.n4852 451.765
R13976 dvss.t1207 dvss 446.743
R13977 dvss.t1998 dvss.t1211 446.743
R13978 dvss.t1020 dvss.t591 446.743
R13979 dvss.t1089 dvss.t1173 446.743
R13980 dvss dvss.t191 446.743
R13981 dvss.t2232 dvss 446.743
R13982 dvss.t1509 dvss 446.743
R13983 dvss.t2184 dvss 446.743
R13984 dvss.t223 dvss 446.038
R13985 dvss.t815 dvss 446.038
R13986 dvss.n1692 dvss.n1594 445.116
R13987 dvss.t1085 dvss.n6334 441.038
R13988 dvss.t1319 dvss.n6251 441.038
R13989 dvss dvss.t720 438.315
R13990 dvss.t559 dvss.t991 438.315
R13991 dvss.t436 dvss.t1170 438.315
R13992 dvss.t874 dvss.t2072 438.315
R13993 dvss.t1965 dvss.t1251 438.315
R13994 dvss.t0 dvss.t209 438.315
R13995 dvss.n6926 dvss.n48 432.788
R13996 dvss.n678 dvss.n675 432.788
R13997 dvss.n6185 dvss.n772 432.788
R13998 dvss.n1023 dvss.n1020 432.788
R13999 dvss.n2082 dvss.n1422 432.788
R14000 dvss.n1915 dvss.n1914 432.788
R14001 dvss.n1797 dvss.n1796 432.788
R14002 dvss.n216 dvss.n185 432.788
R14003 dvss.n5655 dvss.n5654 432.788
R14004 dvss.t1018 dvss.t577 429.885
R14005 dvss.t1994 dvss 429.885
R14006 dvss.t316 dvss.t185 429.885
R14007 dvss.t630 dvss.t938 429.885
R14008 dvss.t25 dvss.t1205 429.885
R14009 dvss.t1691 dvss.t320 421.457
R14010 dvss.t728 dvss.t1193 421.457
R14011 dvss dvss.t1050 421.457
R14012 dvss.n3337 dvss.n3336 417.005
R14013 dvss.t595 dvss 413.027
R14014 dvss dvss.t2138 413.027
R14015 dvss.t886 dvss 413.027
R14016 dvss dvss.t866 413.027
R14017 dvss.t924 dvss 413.027
R14018 dvss.t1498 dvss.n4545 413.027
R14019 dvss dvss.t789 413.027
R14020 dvss.t790 dvss.t1820 413.027
R14021 dvss.t2038 dvss.t1983 413.027
R14022 dvss.n6913 dvss.t1231 410.247
R14023 dvss.n674 dvss.t365 410.247
R14024 dvss.n6172 dvss.t778 410.247
R14025 dvss.n1019 dvss.t14 410.247
R14026 dvss.n2069 dvss.t1348 410.247
R14027 dvss.n1902 dvss.t981 410.247
R14028 dvss.n1795 dvss.t2222 410.247
R14029 dvss.n208 dvss.t1128 410.247
R14030 dvss.n1068 dvss.t1295 410.247
R14031 dvss.t1904 dvss.t1402 404.599
R14032 dvss.n2742 dvss.t829 404.599
R14033 dvss dvss.t1111 404.599
R14034 dvss.n3908 dvss.t2183 404.599
R14035 dvss.t2119 dvss.t2111 404.599
R14036 dvss.t1437 dvss.t948 404.599
R14037 dvss.n6637 dvss.n238 403.825
R14038 dvss.n3197 dvss.n3193 403.825
R14039 dvss.n6927 dvss.t1225 401.229
R14040 dvss.t367 dvss.n682 401.229
R14041 dvss.n6186 dvss.t786 401.229
R14042 dvss.t10 dvss.n1027 401.229
R14043 dvss.n2083 dvss.t1342 401.229
R14044 dvss.t975 dvss.n1929 401.229
R14045 dvss.n1814 dvss.t2216 401.229
R14046 dvss.t1132 dvss.n217 401.229
R14047 dvss.n5653 dvss.t1297 401.229
R14048 dvss.n6902 dvss.n6900 396.721
R14049 dvss.n670 dvss.n662 396.721
R14050 dvss.n6161 dvss.n6159 396.721
R14051 dvss.n1015 dvss.n1007 396.721
R14052 dvss.n2058 dvss.n2056 396.721
R14053 dvss.n1503 dvss.n1502 396.721
R14054 dvss.n1594 dvss.n1577 396.721
R14055 dvss.n206 dvss.n189 396.721
R14056 dvss.n972 dvss.n971 396.721
R14057 dvss.t1441 dvss 396.17
R14058 dvss.t394 dvss.t162 396.17
R14059 dvss.n3161 dvss.n238 395.663
R14060 dvss.n3254 dvss.n3253 394.031
R14061 dvss.n3254 dvss.n3160 394.031
R14062 dvss.n3264 dvss.n3161 394.031
R14063 dvss.n4803 dvss.n4802 392.283
R14064 dvss.n4802 dvss.n4801 392.283
R14065 dvss.n4801 dvss.n2325 392.283
R14066 dvss.n6280 dvss.n6278 389.37
R14067 dvss.n5571 dvss.n524 389.37
R14068 dvss.t1888 dvss.n2988 387.74
R14069 dvss.t711 dvss.t645 387.74
R14070 dvss dvss.t1223 387.74
R14071 dvss.t449 dvss.t1866 387.74
R14072 dvss.t175 dvss.t2032 387.74
R14073 dvss.t986 dvss.t954 387.74
R14074 dvss dvss.t939 387.74
R14075 dvss.t1841 dvss.t1828 387.74
R14076 dvss.t1894 dvss.t1891 387.74
R14077 dvss.n1772 dvss.n1557 380.784
R14078 dvss.n3240 dvss.n3239 379.724
R14079 dvss dvss.t1525 379.31
R14080 dvss.t136 dvss.t2081 379.31
R14081 dvss.t1241 dvss.t874 379.31
R14082 dvss.t1472 dvss.t986 379.31
R14083 dvss.t939 dvss 379.31
R14084 dvss.t2233 dvss.t630 379.31
R14085 dvss.t1205 dvss.t21 379.31
R14086 dvss.n436 dvss.t253 379.31
R14087 dvss.t30 dvss.t1970 370.882
R14088 dvss.t22 dvss.t1428 370.882
R14089 dvss.t938 dvss.t25 370.882
R14090 dvss.t1284 dvss.t936 370.882
R14091 dvss.t789 dvss 370.882
R14092 dvss.t1910 dvss.t722 370.882
R14093 dvss.t798 dvss 370.882
R14094 dvss.n6314 dvss.n6313 368.271
R14095 dvss.n6241 dvss.n502 368.271
R14096 dvss.n3206 dvss.n3193 366.872
R14097 dvss.n3207 dvss.n3206 363.512
R14098 dvss.n3221 dvss.n3185 363.512
R14099 dvss.n3224 dvss.n3223 363.512
R14100 dvss.n3240 dvss.n3238 363.512
R14101 dvss dvss.t593 362.452
R14102 dvss.t2138 dvss 362.452
R14103 dvss.t1050 dvss 362.452
R14104 dvss.n6491 dvss.n6429 358.591
R14105 dvss.n4310 dvss.n4308 358.401
R14106 dvss.n1571 dvss.t759 349.909
R14107 dvss.t400 dvss.n1687 349.909
R14108 dvss.n7012 dvss.t1649 348.875
R14109 dvss.t870 dvss.t879 345.594
R14110 dvss dvss.t1207 345.594
R14111 dvss dvss.t599 345.594
R14112 dvss.t2081 dvss.t142 345.594
R14113 dvss.t2177 dvss.t1089 345.594
R14114 dvss.t1714 dvss.t898 345.594
R14115 dvss.n3208 dvss.t535 344.579
R14116 dvss.n6280 dvss.n6279 342.301
R14117 dvss.n6293 dvss.n6292 342.301
R14118 dvss.n6308 dvss.n477 342.301
R14119 dvss.n6315 dvss.n6314 342.301
R14120 dvss.n6209 dvss.n524 342.301
R14121 dvss.n6221 dvss.n6220 342.301
R14122 dvss.n6224 dvss.n6223 342.301
R14123 dvss.n6241 dvss.n6240 342.301
R14124 dvss.t469 dvss.n3906 337.166
R14125 dvss.t1392 dvss.t2173 337.166
R14126 dvss dvss.t923 337.166
R14127 dvss.t1838 dvss.t1386 337.166
R14128 dvss.t539 dvss.n3222 337.005
R14129 dvss.n6460 dvss.n6459 332.075
R14130 dvss.n6491 dvss.n6437 332.075
R14131 dvss.n6652 dvss.n6651 332.075
R14132 dvss.n6899 dvss.n66 332.075
R14133 dvss.n694 dvss.n597 332.075
R14134 dvss.n6714 dvss.n124 332.075
R14135 dvss.n633 dvss.n629 332.075
R14136 dvss.n661 dvss.n609 332.075
R14137 dvss.n5616 dvss.n5615 332.075
R14138 dvss.n6158 dvss.n790 332.075
R14139 dvss.n1039 dvss.n989 332.075
R14140 dvss.n1055 dvss.n1054 332.075
R14141 dvss.n1381 dvss.n1380 332.075
R14142 dvss.n5730 dvss.n890 332.075
R14143 dvss.n1955 dvss.n1954 332.075
R14144 dvss.n2055 dvss.n1440 332.075
R14145 dvss.n1848 dvss.n1524 332.075
R14146 dvss.n1874 dvss.n1873 332.075
R14147 dvss.t1677 dvss.t2019 331.955
R14148 dvss.t2019 dvss.t291 331.955
R14149 dvss.n4803 dvss.n2324 329.036
R14150 dvss.t1395 dvss.t438 328.736
R14151 dvss.t150 dvss.t394 328.736
R14152 dvss.t1433 dvss.t1179 328.736
R14153 dvss.t2093 dvss.t1431 328.736
R14154 dvss.t432 dvss 328.736
R14155 dvss.t390 dvss.t1280 328.736
R14156 dvss.t1352 dvss.t82 328.736
R14157 dvss.t396 dvss.t1040 327.353
R14158 dvss.n4852 dvss.n4850 321.882
R14159 dvss.t726 dvss.t527 320.307
R14160 dvss.t958 dvss 320.307
R14161 dvss.t1938 dvss.t687 320.307
R14162 dvss.t2175 dvss.t1711 320.307
R14163 dvss.t930 dvss.t1869 320.307
R14164 dvss.t971 dvss 320.307
R14165 dvss.t1029 dvss.t757 317.724
R14166 dvss.t396 dvss.t551 317.724
R14167 dvss.t624 dvss.t557 311.877
R14168 dvss dvss.t575 311.877
R14169 dvss.t2089 dvss 311.877
R14170 dvss dvss.t2117 311.877
R14171 dvss dvss.t852 311.877
R14172 dvss.n2943 dvss.t625 307.536
R14173 dvss.n2867 dvss.t674 307.536
R14174 dvss.n3712 dvss.t618 307.536
R14175 dvss.n3724 dvss.t1088 307.536
R14176 dvss.n3724 dvss.t1962 307.536
R14177 dvss.n3933 dvss.t1210 307.536
R14178 dvss.n3939 dvss.t1436 307.536
R14179 dvss.n4123 dvss.t1196 307.536
R14180 dvss.n4177 dvss.t378 307.536
R14181 dvss.n4248 dvss.t631 307.536
R14182 dvss.n4242 dvss.t1206 307.536
R14183 dvss.t1477 dvss.n6291 306.646
R14184 dvss.n525 dvss.t1378 306.646
R14185 dvss.n2573 dvss.t17 304.238
R14186 dvss.n3111 dvss.t389 304.238
R14187 dvss.n2773 dvss.t897 304.238
R14188 dvss.n3890 dvss.t1503 304.238
R14189 dvss.n3889 dvss.t1993 304.238
R14190 dvss.n2375 dvss.t772 304.238
R14191 dvss.n4301 dvss.t2172 304.238
R14192 dvss.n2295 dvss.n2294 303.817
R14193 dvss.t2103 dvss 303.449
R14194 dvss.t424 dvss.t555 303.449
R14195 dvss dvss.t388 303.449
R14196 dvss.t1334 dvss 303.449
R14197 dvss.t1960 dvss 303.449
R14198 dvss.t2048 dvss.t322 303.449
R14199 dvss.t1255 dvss.t1530 303.449
R14200 dvss.t1209 dvss 303.449
R14201 dvss.t1968 dvss 303.449
R14202 dvss.t1195 dvss 303.449
R14203 dvss.t2111 dvss.t794 303.449
R14204 dvss.n6927 dvss.t1227 302.05
R14205 dvss.n682 dvss.t363 302.05
R14206 dvss.n6186 dvss.t782 302.05
R14207 dvss.n1027 dvss.t8 302.05
R14208 dvss.n2083 dvss.t1344 302.05
R14209 dvss.n1929 dvss.t977 302.05
R14210 dvss.n1814 dvss.t2218 302.05
R14211 dvss.n217 dvss.t1126 302.05
R14212 dvss.t1291 dvss.n5653 302.05
R14213 dvss.n6336 dvss.t1446 300.943
R14214 dvss.n6252 dvss.t675 300.943
R14215 dvss.t1066 dvss.n24 297.485
R14216 dvss.n6648 dvss.t909 297.485
R14217 dvss.n690 dvss.t1559 297.485
R14218 dvss.t1368 dvss.n526 297.485
R14219 dvss.n5612 dvss.t484 297.485
R14220 dvss.n1035 dvss.t2159 297.485
R14221 dvss.t607 dvss.n1349 297.485
R14222 dvss.n1984 dvss.t277 297.485
R14223 dvss.n1834 dvss.t109 297.485
R14224 dvss.n3265 dvss.n3160 295.522
R14225 dvss.t1404 dvss 295.019
R14226 dvss.t567 dvss.t1018 295.019
R14227 dvss dvss.t864 295.019
R14228 dvss.t929 dvss 295.019
R14229 dvss.n4192 dvss.t923 295.019
R14230 dvss.t201 dvss.t316 295.019
R14231 dvss.t1981 dvss.t2038 295.019
R14232 dvss.n6913 dvss.t1229 293.034
R14233 dvss.t359 dvss.n674 293.034
R14234 dvss.n6172 dvss.t784 293.034
R14235 dvss.t12 dvss.n1019 293.034
R14236 dvss.n2069 dvss.t1346 293.034
R14237 dvss.n1902 dvss.t979 293.034
R14238 dvss.t2220 dvss.n1795 293.034
R14239 dvss.n208 dvss.t1124 293.034
R14240 dvss.t1299 dvss.n1068 293.034
R14241 dvss.n6309 dvss.t1475 292.384
R14242 dvss.t1374 dvss.n6222 292.384
R14243 dvss.n5495 dvss.n1153 291.445
R14244 dvss.n3587 dvss.t1389 290.289
R14245 dvss.n4053 dvss.t1440 290.289
R14246 dvss.t451 dvss.t453 286.591
R14247 dvss.t944 dvss.t1938 286.591
R14248 dvss.t838 dvss.t741 286.591
R14249 dvss.t547 dvss 286.591
R14250 dvss.t2042 dvss.t931 286.591
R14251 dvss dvss.t315 286.591
R14252 dvss.t695 dvss.t1422 286.591
R14253 dvss.t1869 dvss.t964 286.591
R14254 dvss.t191 dvss.t0 286.591
R14255 dvss dvss.t4 286.591
R14256 dvss.t374 dvss 286.591
R14257 dvss.t1674 dvss.t2099 284.077
R14258 dvss.n6479 dvss.t1062 283.649
R14259 dvss.n6659 dvss.t903 283.649
R14260 dvss.n702 dvss.t1555 283.649
R14261 dvss.n648 dvss.t1362 283.649
R14262 dvss.n5622 dvss.t482 283.649
R14263 dvss.n1048 dvss.t2167 283.649
R14264 dvss.n1396 dvss.t615 283.649
R14265 dvss.n1962 dvss.t279 283.649
R14266 dvss.t107 dvss.n1852 283.649
R14267 dvss.n379 dvss.t814 283.474
R14268 dvss.n314 dvss.t1184 282.327
R14269 dvss.n455 dvss.t826 282.327
R14270 dvss.n6630 dvss.t810 282.327
R14271 dvss.n375 dvss.t222 282.327
R14272 dvss.t334 dvss.t330 281.707
R14273 dvss.t330 dvss.t324 281.707
R14274 dvss.t324 dvss.t336 281.707
R14275 dvss.t336 dvss.t326 281.707
R14276 dvss.t326 dvss.t338 281.707
R14277 dvss.t338 dvss.t348 281.707
R14278 dvss.t348 dvss.t328 281.707
R14279 dvss.t328 dvss.t340 281.707
R14280 dvss.t340 dvss.t332 281.707
R14281 dvss.t332 dvss.t344 281.707
R14282 dvss.t344 dvss.t354 281.707
R14283 dvss.t354 dvss.t350 281.707
R14284 dvss.t342 dvss.t346 281.707
R14285 dvss.t352 dvss.t342 281.707
R14286 dvss.t219 dvss.t223 281.707
R14287 dvss.t225 dvss.t219 281.707
R14288 dvss.t221 dvss.t225 281.707
R14289 dvss.t805 dvss.t815 281.707
R14290 dvss.t807 dvss.t805 281.707
R14291 dvss.t813 dvss.t807 281.707
R14292 dvss.n2533 dvss.t1405 281.25
R14293 dvss.n2678 dvss.t457 281.25
R14294 dvss.n3652 dvss.t1552 281.25
R14295 dvss.n311 dvss.t1182 281.13
R14296 dvss.n448 dvss.t828 281.13
R14297 dvss.n6623 dvss.t812 281.13
R14298 dvss.n372 dvss.t224 281.13
R14299 dvss.n376 dvss.t816 281.13
R14300 dvss.n2923 dvss.t560 280.822
R14301 dvss.n3483 dvss.t2188 280.259
R14302 dvss.n3502 dvss.t867 278.589
R14303 dvss.t1211 dvss.t1395 278.161
R14304 dvss.t577 dvss.t1020 278.161
R14305 dvss.t205 dvss 278.161
R14306 dvss.n3533 dvss.t1043 277.952
R14307 dvss.n3993 dvss.t1995 277.724
R14308 dvss.n6900 dvss.n6899 276.731
R14309 dvss.n189 dvss.n124 276.731
R14310 dvss.n662 dvss.n661 276.731
R14311 dvss.n6159 dvss.n6158 276.731
R14312 dvss.n1055 dvss.n972 276.731
R14313 dvss.n1007 dvss.n890 276.731
R14314 dvss.n2056 dvss.n2055 276.731
R14315 dvss.n1874 dvss.n1503 276.731
R14316 dvss.n6569 dvss.n6568 275.899
R14317 dvss.n6568 dvss.n6567 275.899
R14318 dvss.n6646 dvss.n227 275.899
R14319 dvss.n6552 dvss.n6362 275.899
R14320 dvss.n6552 dvss.n6551 275.899
R14321 dvss.n6551 dvss.n6550 275.899
R14322 dvss.n6550 dvss.n6363 275.899
R14323 dvss.n6544 dvss.n6363 275.899
R14324 dvss.n6543 dvss.n6542 275.899
R14325 dvss.n6536 dvss.n6383 275.899
R14326 dvss.n6536 dvss.n6535 275.899
R14327 dvss.n6535 dvss.n6534 275.899
R14328 dvss.n6534 dvss.n6384 275.899
R14329 dvss.n6528 dvss.n6384 275.899
R14330 dvss.n6528 dvss.n6527 275.899
R14331 dvss.n6527 dvss.n6526 275.899
R14332 dvss.n6520 dvss.n6519 275.899
R14333 dvss.n6511 dvss.n6510 275.899
R14334 dvss.n6510 dvss.n6509 275.899
R14335 dvss.n6509 dvss.n6409 275.899
R14336 dvss.n6503 dvss.n6409 275.899
R14337 dvss.n4302 dvss.t371 275.293
R14338 dvss.n4390 dvss.t1049 275.293
R14339 dvss.n4725 dvss.t860 275.293
R14340 dvss.t350 dvss.n6605 271.647
R14341 dvss.n3970 dvss.t1512 270.545
R14342 dvss.n420 dvss.n418 270.307
R14343 dvss.n431 dvss.n418 270.307
R14344 dvss.n430 dvss.n420 270.307
R14345 dvss.n431 dvss.n430 270.307
R14346 dvss.t2173 dvss.t436 269.733
R14347 dvss.t2072 dvss 269.733
R14348 dvss.t692 dvss.t1304 269.733
R14349 dvss.t2130 dvss 269.733
R14350 dvss.n4517 dvss.t2297 265.512
R14351 dvss.t1473 dvss.n6309 263.858
R14352 dvss.n6222 dvss.t1380 263.858
R14353 dvss.n2455 dvss.t2269 262.784
R14354 dvss.n2456 dvss.t2279 262.784
R14355 dvss.n2578 dvss.t2298 262.784
R14356 dvss.n2586 dvss.t2277 262.784
R14357 dvss.n2587 dvss.t2286 262.784
R14358 dvss.n2879 dvss.t2318 262.784
R14359 dvss.n2880 dvss.t2240 262.784
R14360 dvss.n3073 dvss.t2323 262.784
R14361 dvss.n3074 dvss.t2248 262.784
R14362 dvss.n2715 dvss.t2294 262.784
R14363 dvss.n2717 dvss.t2316 262.784
R14364 dvss.n3361 dvss.t2301 262.784
R14365 dvss.n3362 dvss.t2321 262.784
R14366 dvss.n3666 dvss.t2254 262.784
R14367 dvss.n3668 dvss.t2258 262.784
R14368 dvss.n3860 dvss.t2266 262.784
R14369 dvss.n3861 dvss.t2272 262.784
R14370 dvss.n3924 dvss.t2267 262.784
R14371 dvss.n3926 dvss.t2273 262.784
R14372 dvss.n3537 dvss.t2256 262.784
R14373 dvss.n3538 dvss.t2263 262.784
R14374 dvss.n4337 dvss.t2314 262.784
R14375 dvss.n4339 dvss.t2255 262.784
R14376 dvss.n2335 dvss.t2308 262.784
R14377 dvss.n2336 dvss.t2246 262.784
R14378 dvss.n4500 dvss.t2322 262.784
R14379 dvss.n4501 dvss.t2328 262.784
R14380 dvss.n4625 dvss.t2331 262.784
R14381 dvss.n4627 dvss.t2333 262.784
R14382 dvss.n4059 dvss.t2335 262.784
R14383 dvss.n4060 dvss.t2338 262.784
R14384 dvss.n4218 dvss.t2342 262.784
R14385 dvss.n4219 dvss.t2238 262.784
R14386 dvss.n2450 dvss.t2239 262.719
R14387 dvss.n2450 dvss.t2341 262.719
R14388 dvss.n2435 dvss.t2336 262.719
R14389 dvss.n2435 dvss.t2327 262.719
R14390 dvss.n2442 dvss.t2280 262.719
R14391 dvss.n2416 dvss.t2249 262.719
R14392 dvss.n2576 dvss.t2289 262.719
R14393 dvss.n2583 dvss.t2325 262.719
R14394 dvss.n2583 dvss.t2317 262.719
R14395 dvss.n2970 dvss.t2332 262.719
R14396 dvss.n2916 dvss.t2295 262.719
R14397 dvss.n2873 dvss.t2290 262.719
R14398 dvss.n3070 dvss.t2303 262.719
R14399 dvss.n3070 dvss.t2260 262.719
R14400 dvss.n2698 dvss.t2340 262.719
R14401 dvss.n3395 dvss.t2307 262.719
R14402 dvss.n3372 dvss.t2337 262.719
R14403 dvss.n3598 dvss.t2251 262.719
R14404 dvss.n2352 dvss.t2324 262.719
R14405 dvss.n2352 dvss.t2276 262.719
R14406 dvss.n4476 dvss.t2247 262.719
R14407 dvss.n2378 dvss.t2313 262.719
R14408 dvss.n4363 dvss.t2312 262.719
R14409 dvss.n4325 dvss.t2320 262.719
R14410 dvss.n4528 dvss.t2284 262.719
R14411 dvss.n4766 dvss.t2330 262.719
R14412 dvss.n4536 dvss.t2315 262.719
R14413 dvss.n4743 dvss.t2250 262.719
R14414 dvss.n4618 dvss.t2334 262.719
R14415 dvss.n4859 dvss.t2259 262.719
R14416 dvss dvss.t352 261.586
R14417 dvss.n6902 dvss.t1429 261.476
R14418 dvss.t1973 dvss.n670 261.476
R14419 dvss.n6161 dvss.t1986 261.476
R14420 dvss.t311 dvss.n1015 261.476
R14421 dvss.n2058 dvss.t357 261.476
R14422 dvss.n1502 dvss.t132 261.476
R14423 dvss.n1577 dvss.t297 261.476
R14424 dvss.t2058 dvss.n206 261.476
R14425 dvss.n971 dvss.t478 261.476
R14426 dvss dvss.t1110 261.303
R14427 dvss.t388 dvss.t603 261.303
R14428 dvss.t698 dvss 261.303
R14429 dvss.t1548 dvss.t888 261.303
R14430 dvss.t700 dvss 261.303
R14431 dvss dvss.t1388 261.303
R14432 dvss.t1547 dvss 261.303
R14433 dvss dvss.t1201 261.303
R14434 dvss dvss.t934 261.303
R14435 dvss.t171 dvss.t1195 261.303
R14436 dvss dvss.t504 261.303
R14437 dvss.t746 dvss 261.303
R14438 dvss dvss.t473 261.303
R14439 dvss dvss.t622 261.303
R14440 dvss.n4236 dvss.t1421 259.51
R14441 dvss.n2486 dvss.t2237 259.082
R14442 dvss.n3099 dvss.t2265 259.082
R14443 dvss.n4319 dvss.t2281 259.082
R14444 dvss.n4783 dvss.t2302 259.082
R14445 dvss.n4718 dvss.t2270 259.082
R14446 dvss.n4697 dvss.t2234 259.082
R14447 dvss.n4866 dvss.t2300 259.082
R14448 dvss.n4991 dvss.t2282 259.082
R14449 dvss.n4978 dvss.t2245 259.082
R14450 dvss.n4965 dvss.t2339 259.082
R14451 dvss.n4940 dvss.t2329 259.082
R14452 dvss.n5027 dvss.t2304 259.082
R14453 dvss.n2538 dvss.t2305 258.176
R14454 dvss.n6310 dvss.n121 256.726
R14455 dvss.n6239 dvss.n6238 256.726
R14456 dvss.t1060 dvss.n6479 255.976
R14457 dvss.n6659 dvss.t901 255.976
R14458 dvss.n702 dvss.t1553 255.976
R14459 dvss.n648 dvss.t1370 255.976
R14460 dvss.n5622 dvss.t490 255.976
R14461 dvss.n1048 dvss.t2161 255.976
R14462 dvss.n1396 dvss.t611 255.976
R14463 dvss.n1962 dvss.t275 255.976
R14464 dvss.n1852 dvss.t111 255.976
R14465 dvss.n2294 dvss.n2292 255.845
R14466 dvss.n2292 dvss.n2291 255.845
R14467 dvss.n2291 dvss.n2290 255.845
R14468 dvss.n2290 dvss.n1240 255.845
R14469 dvss.n1628 dvss.n1240 255.845
R14470 dvss.n1629 dvss.n1628 255.845
R14471 dvss.n1630 dvss.n1629 255.845
R14472 dvss.n1683 dvss.n1682 255.845
R14473 dvss.n1682 dvss.n1681 255.845
R14474 dvss.n1678 dvss.n1677 255.845
R14475 dvss.n1677 dvss.n1675 255.845
R14476 dvss.n1673 dvss.n1671 255.845
R14477 dvss.n4749 dvss.t793 255.326
R14478 dvss.n4723 dvss.t851 255.326
R14479 dvss.n4575 dvss.t2112 255.326
R14480 dvss.n3222 dvss.t531 253.702
R14481 dvss.n1674 dvss.n1673 253.18
R14482 dvss.n4597 dvss.t2235 253.029
R14483 dvss.t1401 dvss 252.875
R14484 dvss.t2046 dvss 252.875
R14485 dvss.t1336 dvss.t95 252.875
R14486 dvss.t768 dvss 252.875
R14487 dvss.t872 dvss 252.875
R14488 dvss dvss.t1328 252.875
R14489 dvss.t2189 dvss 252.875
R14490 dvss.t472 dvss.t2091 252.875
R14491 dvss.t470 dvss.t2090 252.875
R14492 dvss.t1439 dvss 252.875
R14493 dvss.t377 dvss.t2140 252.875
R14494 dvss dvss.t98 252.875
R14495 dvss dvss.t2226 252.875
R14496 dvss dvss.t177 252.875
R14497 dvss.n1671 dvss.n1670 252.209
R14498 dvss.t2021 dvss.t1617 252.159
R14499 dvss.t1617 dvss.t529 252.159
R14500 dvss.t529 dvss.t1677 252.159
R14501 dvss.n6813 dvss.n6812 251.879
R14502 dvss.n6817 dvss.n6806 251.879
R14503 dvss.n6820 dvss.n23 251.879
R14504 dvss.n6951 dvss.n6950 251.879
R14505 dvss.n6951 dvss.n18 251.879
R14506 dvss.n6967 dvss.n18 251.879
R14507 dvss.n6969 dvss.n12 251.879
R14508 dvss.n6980 dvss.n12 251.879
R14509 dvss.n6983 dvss.n6982 251.879
R14510 dvss.n6740 dvss.n6739 251.879
R14511 dvss.n6754 dvss.n103 251.879
R14512 dvss.n6757 dvss.n6756 251.879
R14513 dvss.n6770 dvss.n6769 251.879
R14514 dvss.n6772 dvss.n6770 251.879
R14515 dvss.n6772 dvss.n6771 251.879
R14516 dvss.n6786 dvss.n6785 251.879
R14517 dvss.n6786 dvss.n78 251.879
R14518 dvss.n6859 dvss.n79 251.879
R14519 dvss.n5925 dvss.n5924 251.879
R14520 dvss.n5930 dvss.n5929 251.879
R14521 dvss.n5933 dvss.n5932 251.879
R14522 dvss.n5979 dvss.n5978 251.879
R14523 dvss.n5980 dvss.n5979 251.879
R14524 dvss.n5981 dvss.n5980 251.879
R14525 dvss.n5986 dvss.n5985 251.879
R14526 dvss.n5988 dvss.n5986 251.879
R14527 dvss.n5991 dvss.n5990 251.879
R14528 dvss.n5999 dvss.n5998 251.879
R14529 dvss.n6003 dvss.n6002 251.879
R14530 dvss.n6006 dvss.n6005 251.879
R14531 dvss.n6009 dvss.n6008 251.879
R14532 dvss.n6010 dvss.n6009 251.879
R14533 dvss.n6011 dvss.n6010 251.879
R14534 dvss.n6016 dvss.n6015 251.879
R14535 dvss.n6016 dvss.n120 251.879
R14536 dvss.n6718 dvss.n6717 251.879
R14537 dvss.n5846 dvss.n5845 251.879
R14538 dvss.n5860 dvss.n832 251.879
R14539 dvss.n5863 dvss.n5862 251.879
R14540 dvss.n5876 dvss.n5875 251.879
R14541 dvss.n5878 dvss.n5876 251.879
R14542 dvss.n5878 dvss.n5877 251.879
R14543 dvss.n5892 dvss.n5891 251.879
R14544 dvss.n5892 dvss.n807 251.879
R14545 dvss.n6118 dvss.n808 251.879
R14546 dvss.n5754 dvss.n5753 251.879
R14547 dvss.n5769 dvss.n868 251.879
R14548 dvss.n5786 dvss.n5785 251.879
R14549 dvss.n5787 dvss.n857 251.879
R14550 dvss.n5799 dvss.n857 251.879
R14551 dvss.n5800 dvss.n5799 251.879
R14552 dvss.n5820 dvss.n850 251.879
R14553 dvss.n5821 dvss.n5820 251.879
R14554 dvss.n5824 dvss.n5823 251.879
R14555 dvss.n2012 dvss.n2011 251.879
R14556 dvss.n2006 dvss.n2005 251.879
R14557 dvss.n1348 dvss.n1347 251.879
R14558 dvss.n2108 dvss.n2107 251.879
R14559 dvss.n2109 dvss.n2108 251.879
R14560 dvss.n2111 dvss.n2109 251.879
R14561 dvss.n2113 dvss.n887 251.879
R14562 dvss.n5733 dvss.n887 251.879
R14563 dvss.n5751 dvss.n875 251.879
R14564 dvss.n1643 dvss.n1642 251.879
R14565 dvss.n1639 dvss.n1638 251.879
R14566 dvss.n1987 dvss.n1986 251.879
R14567 dvss.n1990 dvss.n1989 251.879
R14568 dvss.n1991 dvss.n1990 251.879
R14569 dvss.n1992 dvss.n1991 251.879
R14570 dvss.n1997 dvss.n1996 251.879
R14571 dvss.n1999 dvss.n1997 251.879
R14572 dvss.n2015 dvss.n2014 251.879
R14573 dvss.n1670 dvss.n1669 251.879
R14574 dvss.n1632 dvss.n1631 251.879
R14575 dvss.n1635 dvss.n1634 251.879
R14576 dvss.n1664 dvss.n1662 251.879
R14577 dvss.n1662 dvss.n1661 251.879
R14578 dvss.n1661 dvss.n1660 251.879
R14579 dvss.n1656 dvss.n1655 251.879
R14580 dvss.n1655 dvss.n1654 251.879
R14581 dvss.n1651 dvss.n1650 251.879
R14582 dvss dvss.t221 251.524
R14583 dvss dvss.t813 251.524
R14584 dvss.n6480 dvss.n11 249.058
R14585 dvss.n6862 dvss.n6861 249.058
R14586 dvss.n6715 dvss.n122 249.058
R14587 dvss.n651 dvss.n507 249.058
R14588 dvss.n6121 dvss.n6120 249.058
R14589 dvss.n1051 dvss.n849 249.058
R14590 dvss.n5731 dvss.n888 249.058
R14591 dvss.n2018 dvss.n2017 249.058
R14592 dvss.n1851 dvss.n1506 249.058
R14593 dvss.n1679 dvss.t128 247.851
R14594 dvss.t1519 dvss.n226 247.16
R14595 dvss.n6392 dvss.t1078 247.16
R14596 dvss.n3670 dvss.t1329 246.506
R14597 dvss.n4054 dvss.t90 246.506
R14598 dvss.n3208 dvss.t533 246.127
R14599 dvss.n1762 dvss.t397 245.276
R14600 dvss.n5125 dvss.t755 245.276
R14601 dvss.t454 dvss.t1267 244.445
R14602 dvss dvss.t1107 244.445
R14603 dvss dvss.t1941 244.445
R14604 dvss.t598 dvss 244.445
R14605 dvss.t492 dvss.t1209 244.445
R14606 dvss.t2171 dvss.t215 244.445
R14607 dvss.n6544 dvss.t1305 244.286
R14608 dvss.t56 dvss.n334 243.903
R14609 dvss.n3239 dvss.t1466 242.165
R14610 dvss.n2778 dvss.t590 242.067
R14611 dvss.n3765 dvss.t147 242.067
R14612 dvss.n2830 dvss.t2135 240.948
R14613 dvss.n3822 dvss.t887 240.948
R14614 dvss.n4142 dvss.t2131 240.948
R14615 dvss.n6611 dvss.t1164 240.701
R14616 dvss.t1035 dvss.n1683 239.856
R14617 dvss.n3484 dvss.t1244 239.4
R14618 dvss.n4274 dvss.t194 238.44
R14619 dvss.t402 dvss.n1674 237.19
R14620 dvss.n7007 dvss.t1616 236.975
R14621 dvss.n7009 dvss.t1676 236.975
R14622 dvss.n424 dvss.t1583 236.149
R14623 dvss.n2566 dvss.t1441 236.016
R14624 dvss.n3124 dvss.t1223 236.016
R14625 dvss.t1208 dvss.t840 236.016
R14626 dvss.t1245 dvss.t319 236.016
R14627 dvss.t410 dvss.t30 236.016
R14628 dvss.t508 dvss.t2089 236.016
R14629 dvss.t422 dvss.t22 236.016
R14630 dvss.t936 dvss.t1426 236.016
R14631 dvss.t1948 dvss 236.016
R14632 dvss.t2117 dvss.t724 236.016
R14633 dvss.n2302 dvss.t1598 236.011
R14634 dvss.n2301 dvss.t1637 236.011
R14635 dvss.n4847 dvss.t1658 236.011
R14636 dvss.n4844 dvss.t1643 236.011
R14637 dvss.n4843 dvss.t1604 236.011
R14638 dvss.n4842 dvss.t1625 236.011
R14639 dvss.n4838 dvss.t1619 236.011
R14640 dvss.n4839 dvss.t1640 236.011
R14641 dvss.n4834 dvss.t1634 236.011
R14642 dvss.n4835 dvss.t1667 236.011
R14643 dvss.n4830 dvss.t1664 236.011
R14644 dvss.n4831 dvss.t1646 236.011
R14645 dvss.n2321 dvss.t1670 236.011
R14646 dvss.n2319 dvss.t1622 236.011
R14647 dvss.n2318 dvss.t1592 236.011
R14648 dvss.n2316 dvss.t1661 236.011
R14649 dvss.n2315 dvss.t1652 236.011
R14650 dvss.n2309 dvss.t1679 236.011
R14651 dvss.n2310 dvss.t1628 236.011
R14652 dvss.n2312 dvss.t1595 236.011
R14653 dvss.n2799 dvss.t1021 235.607
R14654 dvss.n2381 dvss.t1984 235.607
R14655 dvss.n3823 dvss.t734 234.239
R14656 dvss.n4065 dvss.t1969 234.239
R14657 dvss.n2918 dvss.t1013 233.732
R14658 dvss.n2557 dvss.t880 233.459
R14659 dvss.n3423 dvss.t2180 233.459
R14660 dvss.n3707 dvss.t869 233.459
R14661 dvss.n4799 dvss.t1653 232.499
R14662 dvss.n4805 dvss.t1680 232.499
R14663 dvss.n3621 dvss.t691 231.529
R14664 dvss.n6812 dvss.n6811 230.888
R14665 dvss.n6739 dvss.n111 230.888
R14666 dvss.n5924 dvss.n5923 230.888
R14667 dvss.n5998 dvss.n5997 230.888
R14668 dvss.n5845 dvss.n840 230.888
R14669 dvss.n5754 dvss.n5752 230.888
R14670 dvss.n2013 dvss.n2012 230.888
R14671 dvss.n1649 dvss.n1643 230.888
R14672 dvss.n3119 dvss.t1396 230.488
R14673 dvss.n3057 dvss.t1054 230.488
R14674 dvss.n3343 dvss.t1964 230.488
R14675 dvss.n3534 dvss.t1333 229.833
R14676 dvss.n2546 dvss.t1573 227.68
R14677 dvss.n3800 dvss.t2082 227.68
R14678 dvss.n3461 dvss.t1095 227.68
R14679 dvss.t428 dvss.t37 227.587
R14680 dvss.t563 dvss.t995 227.587
R14681 dvss dvss.t1579 227.587
R14682 dvss.t593 dvss.t1171 227.587
R14683 dvss.t462 dvss 227.587
R14684 dvss dvss.t418 227.587
R14685 dvss.t690 dvss.t862 227.587
R14686 dvss.t122 dvss.t89 227.587
R14687 dvss.t1286 dvss.t189 227.587
R14688 dvss.n3350 dvss.t1942 227.256
R14689 dvss.n2854 dvss.t1266 226.882
R14690 dvss.n3753 dvss.t284 226.882
R14691 dvss.n3753 dvss.t1248 226.882
R14692 dvss.n3632 dvss.t743 226.882
R14693 dvss.n3859 dvss.t2011 226.882
R14694 dvss.n4124 dvss.t1508 226.882
R14695 dvss.n4044 dvss.t1453 226.882
R14696 dvss.n4024 dvss.t380 226.882
R14697 dvss.n4217 dvss.t2005 226.882
R14698 dvss.n5847 dvss.t667 226.6
R14699 dvss.n6741 dvss.t1406 226.6
R14700 dvss.n6816 dvss.t1097 226.6
R14701 dvss.n5928 dvss.t2199 226.6
R14702 dvss.n6001 dvss.t997 226.6
R14703 dvss.n5767 dvss.t1119 226.6
R14704 dvss.t1494 dvss.n2010 226.6
R14705 dvss.t1315 dvss.n1641 226.6
R14706 dvss.n1666 dvss.t267 226.6
R14707 dvss.n2706 dvss.t830 223.748
R14708 dvss.n3586 dvss.t1695 223.662
R14709 dvss.n6999 dvss.t1673 223.559
R14710 dvss.n3238 dvss.n3237 223.409
R14711 dvss.n2421 dvss.t1571 223.315
R14712 dvss.n2972 dvss.t1015 223.315
R14713 dvss.n3642 dvss.t395 223.315
R14714 dvss.n3963 dvss.t466 223.315
R14715 dvss.n3972 dvss.t1236 223.315
R14716 dvss.n2328 dvss.t308 223.315
R14717 dvss.n2392 dvss.t544 223.315
R14718 dvss.n2541 dvss.t2268 221.972
R14719 dvss.n2713 dvss.t2293 221.958
R14720 dvss.n4380 dvss.t1895 221.793
R14721 dvss.n6818 dvss.t1101 221.619
R14722 dvss.t1410 dvss.n6755 221.619
R14723 dvss.t2197 dvss.n5931 221.619
R14724 dvss.t999 dvss.n6004 221.619
R14725 dvss.t669 dvss.n5861 221.619
R14726 dvss.n5768 dvss.t1115 221.619
R14727 dvss.n2008 dvss.t1488 221.619
R14728 dvss.n1637 dvss.t1309 221.619
R14729 dvss.n1665 dvss.t261 221.619
R14730 dvss.n6518 dvss.n6517 220.345
R14731 dvss.n4507 dvss.t1845 220.222
R14732 dvss.n2483 dvss.t1927 220.082
R14733 dvss.n2540 dvss.t1952 219.972
R14734 dvss.t1749 dvss.t914 219.157
R14735 dvss.t1338 dvss.t2189 219.157
R14736 dvss.n3760 dvss.t1978 219.157
R14737 dvss.t1979 dvss.t160 219.157
R14738 dvss.t416 dvss.t1450 219.157
R14739 dvss.t1189 dvss 219.157
R14740 dvss.t545 dvss 219.157
R14741 dvss.t2144 dvss 219.157
R14742 dvss dvss.t924 219.157
R14743 dvss.t203 dvss.t2070 219.157
R14744 dvss dvss.t776 219.157
R14745 dvss.t1058 dvss.t962 219.157
R14746 dvss.t2098 dvss.t1674 218.643
R14747 dvss.n4312 dvss.t2278 218.607
R14748 dvss.n4385 dvss.t1892 218.428
R14749 dvss.n2427 dvss.t2343 218.308
R14750 dvss.n2683 dvss.t2253 218.308
R14751 dvss.n2676 dvss.t2319 218.308
R14752 dvss.n2749 dvss.t2310 218.308
R14753 dvss.n2790 dvss.t2275 218.308
R14754 dvss.n2390 dvss.t2285 218.308
R14755 dvss.n4134 dvss.t2274 218.308
R14756 dvss.n4185 dvss.t2264 218.308
R14757 dvss.n2714 dvss.t1879 217.934
R14758 dvss.n218 dvss.n183 217.099
R14759 dvss.n1120 dvss.n1118 217.099
R14760 dvss.n45 dvss.n44 217.097
R14761 dvss.n684 dvss.n683 217.097
R14762 dvss.n769 dvss.n768 217.097
R14763 dvss.n1029 dvss.n1028 217.097
R14764 dvss.n1419 dvss.n1418 217.097
R14765 dvss.n1930 dvss.n1471 217.097
R14766 dvss.n1819 dvss.n1818 217.097
R14767 dvss.n2885 dvss.t1698 216.933
R14768 dvss.n2544 dvss.t1761 216.632
R14769 dvss.n4320 dvss.t1816 216.632
R14770 dvss.n2611 dvss.t1958 216.624
R14771 dvss.n4319 dvss.t1896 215.905
R14772 dvss.n2723 dvss.t2309 215.754
R14773 dvss.n3196 dvss.t1037 214.554
R14774 dvss.n2477 dvss.t1809 214.456
R14775 dvss.n2454 dvss.t1808 214.456
R14776 dvss.n2477 dvss.t1739 214.456
R14777 dvss.n2454 dvss.t1738 214.456
R14778 dvss.n2455 dvss.t1722 214.456
R14779 dvss.n2455 dvss.t1721 214.456
R14780 dvss.n2456 dvss.t1930 214.456
R14781 dvss.n2456 dvss.t1929 214.456
R14782 dvss.n2585 dvss.t1857 214.456
R14783 dvss.n2579 dvss.t1856 214.456
R14784 dvss.n2585 dvss.t1796 214.456
R14785 dvss.n2579 dvss.t1795 214.456
R14786 dvss.n2578 dvss.t1877 214.456
R14787 dvss.n2578 dvss.t1876 214.456
R14788 dvss.n2569 dvss.t1957 214.456
R14789 dvss.n2428 dvss.t1807 214.456
R14790 dvss.n2636 dvss.t1806 214.456
R14791 dvss.n2420 dvss.t1762 214.456
R14792 dvss.n2541 dvss.t1953 214.456
R14793 dvss.n2539 dvss.t1906 214.456
R14794 dvss.n2537 dvss.t1905 214.456
R14795 dvss.n2445 dvss.t1802 214.456
R14796 dvss.n2485 dvss.t1801 214.456
R14797 dvss.n2440 dvss.t1719 214.456
R14798 dvss.n2444 dvss.t1718 214.456
R14799 dvss.n2440 dvss.t1928 214.456
R14800 dvss.n2522 dvss.t1832 214.456
R14801 dvss.n2439 dvss.t1831 214.456
R14802 dvss.n2522 dvss.t1786 214.456
R14803 dvss.n2439 dvss.t1785 214.456
R14804 dvss.n2586 dvss.t1702 214.456
R14805 dvss.n2586 dvss.t1701 214.456
R14806 dvss.n2587 dvss.t1903 214.456
R14807 dvss.n2587 dvss.t1902 214.456
R14808 dvss.n2879 dvss.t1804 214.456
R14809 dvss.n2879 dvss.t1803 214.456
R14810 dvss.n2880 dvss.t1731 214.456
R14811 dvss.n2880 dvss.t1730 214.456
R14812 dvss.n3072 dvss.t1947 214.456
R14813 dvss.n3067 dvss.t1946 214.456
R14814 dvss.n3072 dvss.t1862 214.456
R14815 dvss.n3067 dvss.t1861 214.456
R14816 dvss.n3098 dvss.t1693 214.456
R14817 dvss.n3101 dvss.t1692 214.456
R14818 dvss.n2915 dvss.t1771 214.456
R14819 dvss.n2917 dvss.t1890 214.456
R14820 dvss.n2963 dvss.t1772 214.456
R14821 dvss.n2908 dvss.t1883 214.456
R14822 dvss.n2902 dvss.t1889 214.456
R14823 dvss.n2874 dvss.t1699 214.456
R14824 dvss.n2887 dvss.t1882 214.456
R14825 dvss.n3073 dvss.t1791 214.456
R14826 dvss.n3073 dvss.t1790 214.456
R14827 dvss.n3074 dvss.t1708 214.456
R14828 dvss.n3074 dvss.t1707 214.456
R14829 dvss.n2715 dvss.t1799 214.456
R14830 dvss.n2715 dvss.t1798 214.456
R14831 dvss.n2717 dvss.t1811 214.456
R14832 dvss.n2717 dvss.t1810 214.456
R14833 dvss.n3366 dvss.t1943 214.456
R14834 dvss.n3379 dvss.t1899 214.456
R14835 dvss.n3389 dvss.t1759 214.456
R14836 dvss.n3348 dvss.t1898 214.456
R14837 dvss.n3342 dvss.t1758 214.456
R14838 dvss.n2677 dvss.t1713 214.456
R14839 dvss.n2819 dvss.t1712 214.456
R14840 dvss.n2685 dvss.t1868 214.456
R14841 dvss.n3418 dvss.t1867 214.456
R14842 dvss.n2788 dvss.t1933 214.456
R14843 dvss.n2785 dvss.t1932 214.456
R14844 dvss.n2696 dvss.t1940 214.456
R14845 dvss.n2756 dvss.t1939 214.456
R14846 dvss.n2704 dvss.t1751 214.456
R14847 dvss.n2747 dvss.t1750 214.456
R14848 dvss.n2724 dvss.t1756 214.456
R14849 dvss.n2712 dvss.t1755 214.456
R14850 dvss.n2713 dvss.t1880 214.456
R14851 dvss.n3361 dvss.t1789 214.456
R14852 dvss.n3361 dvss.t1788 214.456
R14853 dvss.n3362 dvss.t1793 214.456
R14854 dvss.n3362 dvss.t1792 214.456
R14855 dvss.n3666 dvss.t1865 214.456
R14856 dvss.n3666 dvss.t1864 214.456
R14857 dvss.n3668 dvss.t1885 214.456
R14858 dvss.n3668 dvss.t1884 214.456
R14859 dvss.n3860 dvss.t1849 214.456
R14860 dvss.n3860 dvss.t1848 214.456
R14861 dvss.n3861 dvss.t1859 214.456
R14862 dvss.n3861 dvss.t1858 214.456
R14863 dvss.n3924 dvss.t1937 214.456
R14864 dvss.n3924 dvss.t1936 214.456
R14865 dvss.n3926 dvss.t1855 214.456
R14866 dvss.n3926 dvss.t1854 214.456
R14867 dvss.n3607 dvss.t1696 214.456
R14868 dvss.n3599 dvss.t1777 214.456
R14869 dvss.n3521 dvss.t1920 214.456
R14870 dvss.n3526 dvss.t1919 214.456
R14871 dvss.n3537 dvss.t1955 214.456
R14872 dvss.n3537 dvss.t1954 214.456
R14873 dvss.n3538 dvss.t1874 214.456
R14874 dvss.n3538 dvss.t1873 214.456
R14875 dvss.n3514 dvss.t1778 214.456
R14876 dvss.n4326 dvss.t1817 214.456
R14877 dvss.n4370 dvss.t1747 214.456
R14878 dvss.n4329 dvss.t1748 214.456
R14879 dvss.n4337 dvss.t1814 214.456
R14880 dvss.n4337 dvss.t1813 214.456
R14881 dvss.n4339 dvss.t1901 214.456
R14882 dvss.n4339 dvss.t1900 214.456
R14883 dvss.n4376 dvss.t1893 214.456
R14884 dvss.n4313 dvss.t1909 214.456
R14885 dvss.n4392 dvss.t1908 214.456
R14886 dvss.n2391 dvss.t1835 214.456
R14887 dvss.n4438 dvss.t1834 214.456
R14888 dvss.n2380 dvss.t1783 214.456
R14889 dvss.n2371 dvss.t1782 214.456
R14890 dvss.n4469 dvss.t1923 214.456
R14891 dvss.n4488 dvss.t1922 214.456
R14892 dvss.n2359 dvss.t1914 214.456
R14893 dvss.n2334 dvss.t1913 214.456
R14894 dvss.n2359 dvss.t1736 214.456
R14895 dvss.n2334 dvss.t1735 214.456
R14896 dvss.n2335 dvss.t1827 214.456
R14897 dvss.n2335 dvss.t1826 214.456
R14898 dvss.n2336 dvss.t1925 214.456
R14899 dvss.n2336 dvss.t1924 214.456
R14900 dvss.n4500 dvss.t1780 214.456
R14901 dvss.n4500 dvss.t1779 214.456
R14902 dvss.n4501 dvss.t1725 214.456
R14903 dvss.n4501 dvss.t1724 214.456
R14904 dvss.n4625 dvss.t1753 214.456
R14905 dvss.n4625 dvss.t1752 214.456
R14906 dvss.n4627 dvss.t1705 214.456
R14907 dvss.n4627 dvss.t1704 214.456
R14908 dvss.n4638 dvss.t1745 214.456
R14909 dvss.n4619 dvss.t1819 214.456
R14910 dvss.n4616 dvss.t1818 214.456
R14911 dvss.n4656 dvss.t1744 214.456
R14912 dvss.n4661 dvss.t1822 214.456
R14913 dvss.n4603 dvss.t1821 214.456
R14914 dvss.n4598 dvss.t1687 214.456
R14915 dvss.n4596 dvss.t1686 214.456
R14916 dvss.n4592 dvss.t1840 214.456
R14917 dvss.n4583 dvss.t1839 214.456
R14918 dvss.n4696 dvss.t1716 214.456
R14919 dvss.n4580 dvss.t1715 214.456
R14920 dvss.n4717 dvss.t1912 214.456
R14921 dvss.n4554 dvss.t1911 214.456
R14922 dvss.n4543 dvss.t1950 214.456
R14923 dvss.n4534 dvss.t1949 214.456
R14924 dvss.n4537 dvss.t1775 214.456
R14925 dvss.n4760 dvss.t1767 214.456
R14926 dvss.n4530 dvss.t1774 214.456
R14927 dvss.n4526 dvss.t1766 214.456
R14928 dvss.n4529 dvss.t1843 214.456
R14929 dvss.n4782 dvss.t1830 214.456
R14930 dvss.n4525 dvss.t1829 214.456
R14931 dvss.n4520 dvss.t1846 214.456
R14932 dvss.n4519 dvss.t1842 214.456
R14933 dvss.n4495 dvss.t1728 214.456
R14934 dvss.n4498 dvss.t1727 214.456
R14935 dvss.n5026 dvss.t1824 214.456
R14936 dvss.n5024 dvss.t1823 214.456
R14937 dvss.n5022 dvss.t1710 214.456
R14938 dvss.n5021 dvss.t1709 214.456
R14939 dvss.n4939 dvss.t1769 214.456
R14940 dvss.n4916 dvss.t1768 214.456
R14941 dvss.n4964 dvss.t1733 214.456
R14942 dvss.n4907 dvss.t1732 214.456
R14943 dvss.n4977 dvss.t1684 214.456
R14944 dvss.n4902 dvss.t1683 214.456
R14945 dvss.n4990 dvss.t1887 214.456
R14946 dvss.n4897 dvss.t1886 214.456
R14947 dvss.n4889 dvss.t1935 214.456
R14948 dvss.n4863 dvss.t1934 214.456
R14949 dvss.n4867 dvss.t1837 214.456
R14950 dvss.n4865 dvss.t1836 214.456
R14951 dvss.n4133 dvss.t1852 214.456
R14952 dvss.n4130 dvss.t1851 214.456
R14953 dvss.n4081 dvss.t1916 214.456
R14954 dvss.n4083 dvss.t1917 214.456
R14955 dvss.n4059 dvss.t1764 214.456
R14956 dvss.n4059 dvss.t1763 214.456
R14957 dvss.n4060 dvss.t1690 214.456
R14958 dvss.n4060 dvss.t1689 214.456
R14959 dvss.n4184 dvss.t1871 214.456
R14960 dvss.n4140 dvss.t1870 214.456
R14961 dvss.n4218 dvss.t1742 214.456
R14962 dvss.n4218 dvss.t1741 214.456
R14963 dvss.n4219 dvss.t1945 214.456
R14964 dvss.n4219 dvss.t1944 214.456
R14965 dvss.n4809 dvss.n2299 213.835
R14966 dvss.n4820 dvss.n2299 213.835
R14967 dvss.n4809 dvss.n2300 213.835
R14968 dvss.n1755 dvss.n1594 212.969
R14969 dvss.n1730 dvss.n1594 212.969
R14970 dvss.t579 dvss.t877 210.728
R14971 dvss dvss.t587 210.728
R14972 dvss.t581 dvss.t97 210.728
R14973 dvss.t1468 dvss 210.728
R14974 dvss.t138 dvss 210.728
R14975 dvss dvss.t313 210.728
R14976 dvss.t502 dvss.t195 210.728
R14977 dvss.n3676 dvss.n3664 210.601
R14978 dvss.n6291 dvss.n487 210.374
R14979 dvss.n6208 dvss.n525 210.374
R14980 dvss.n2755 dvss.n2754 209.989
R14981 dvss.n6983 dvss.n8 209.899
R14982 dvss.n6811 dvss.n79 209.899
R14983 dvss.n5997 dvss.n5991 209.899
R14984 dvss.n6717 dvss.n111 209.899
R14985 dvss.n5923 dvss.n808 209.899
R14986 dvss.n5823 dvss.n840 209.899
R14987 dvss.n5752 dvss.n5751 209.899
R14988 dvss.n2014 dvss.n2013 209.899
R14989 dvss.n1650 dvss.n1649 209.899
R14990 dvss.n2932 dvss.n2931 209.254
R14991 dvss.n2852 dvss.n2851 209.254
R14992 dvss.n3747 dvss.n3745 209.254
R14993 dvss.n3747 dvss.n3746 209.254
R14994 dvss.n3834 dvss.n3833 209.254
R14995 dvss.n3871 dvss.n3856 209.254
R14996 dvss.n3956 dvss.n3955 209.254
R14997 dvss.n4427 dvss.n2396 209.254
R14998 dvss.n4100 dvss.n4099 209.254
R14999 dvss.n2558 dvss.n2535 208.553
R15000 dvss.n3496 dvss.n3471 208.553
R15001 dvss.n3466 dvss.n3465 208.553
R15002 dvss.n4950 dvss.n4914 208.553
R15003 dvss.n2426 dvss.n2425 208.025
R15004 dvss.n2956 dvss.n2925 207.965
R15005 dvss.n2856 dvss.n2855 207.213
R15006 dvss.n3518 dvss.n3517 207.213
R15007 dvss.n4050 dvss.n4048 207.213
R15008 dvss.n6584 dvss.n378 207.213
R15009 dvss.n6593 dvss.n374 207.213
R15010 dvss.n318 dvss.n313 207.213
R15011 dvss.n288 dvss.n287 207.213
R15012 dvss.n292 dvss.n286 207.213
R15013 dvss.n295 dvss.n294 207.213
R15014 dvss.n301 dvss.n283 207.213
R15015 dvss.n304 dvss.n303 207.213
R15016 dvss.n281 dvss.n280 207.213
R15017 dvss.n328 dvss.n309 207.213
R15018 dvss.n453 dvss.n382 207.213
R15019 dvss.n397 dvss.n396 207.213
R15020 dvss.n399 dvss.n398 207.213
R15021 dvss.n405 dvss.n393 207.213
R15022 dvss.n408 dvss.n407 207.213
R15023 dvss.n414 dvss.n390 207.213
R15024 dvss.n388 dvss.n387 207.213
R15025 dvss.n442 dvss.n386 207.213
R15026 dvss.n6628 dvss.n244 207.213
R15027 dvss.n259 dvss.n258 207.213
R15028 dvss.n261 dvss.n260 207.213
R15029 dvss.n267 dvss.n255 207.213
R15030 dvss.n270 dvss.n269 207.213
R15031 dvss.n276 dvss.n252 207.213
R15032 dvss.n250 dvss.n249 207.213
R15033 dvss.n6617 dvss.n248 207.213
R15034 dvss.n347 dvss.n346 207.213
R15035 dvss.n349 dvss.n348 207.213
R15036 dvss.n355 dvss.n343 207.213
R15037 dvss.n358 dvss.n357 207.213
R15038 dvss.n364 dvss.n340 207.213
R15039 dvss.n367 dvss.n366 207.213
R15040 dvss.n6603 dvss.n337 207.213
R15041 dvss.n3815 dvss.n3814 206.909
R15042 dvss.n3818 dvss.n3817 206.909
R15043 dvss.n4178 dvss.n4144 206.909
R15044 dvss.n4176 dvss.n4147 206.909
R15045 dvss.n2813 dvss.n2811 206.02
R15046 dvss.n3785 dvss.n3784 205.899
R15047 dvss.n4161 dvss.n4160 205.899
R15048 dvss.n4287 dvss.n4014 205.899
R15049 dvss.n4070 dvss.n4057 205.541
R15050 dvss.n3775 dvss.n3774 205.481
R15051 dvss.n4280 dvss.n4019 205.481
R15052 dvss.n3487 dvss.n3486 205.078
R15053 dvss.n2809 dvss.n2808 204.692
R15054 dvss.n2694 dvss.n2693 204.692
R15055 dvss.n3798 dvss.n3797 204.692
R15056 dvss.n4174 dvss.n4150 204.692
R15057 dvss.n4157 dvss.n4156 204.692
R15058 dvss.n4021 dvss.n4020 204.692
R15059 dvss.n3561 dvss.n3560 204.457
R15060 dvss.n6357 dvss.n236 204.279
R15061 dvss.n2675 dvss.n2674 204.201
R15062 dvss.n3571 dvss.n3525 204.201
R15063 dvss.n6949 dvss.n24 204.089
R15064 dvss.n6648 dvss.n6647 204.089
R15065 dvss.n690 dvss.n487 204.089
R15066 dvss.n6208 dvss.n526 204.089
R15067 dvss.n5612 dvss.n5610 204.089
R15068 dvss.n1035 dvss.n862 204.089
R15069 dvss.n2105 dvss.n1349 204.089
R15070 dvss.n1985 dvss.n1984 204.089
R15071 dvss.n1834 dvss.n1530 204.089
R15072 dvss.n3046 dvss.n3045 203.619
R15073 dvss.n3491 dvss.n3473 203.619
R15074 dvss.n4443 dvss.n2385 203.619
R15075 dvss.n2964 dvss.n2922 203.526
R15076 dvss.n3779 dvss.n3778 203.526
R15077 dvss.n3964 dvss.n3912 203.526
R15078 dvss.n2367 dvss.n2366 203.526
R15079 dvss.n4131 dvss.n4028 203.526
R15080 dvss.n4196 dvss.n4195 203.526
R15081 dvss.n4229 dvss.n4214 203.526
R15082 dvss.n3869 dvss.n3858 203.016
R15083 dvss.n2394 dvss.n2393 203.016
R15084 dvss.n4091 dvss.n4046 203.016
R15085 dvss.n2836 dvss.n2810 202.724
R15086 dvss.t295 dvss.t1650 202.685
R15087 dvss.n3616 dvss.n3508 202.564
R15088 dvss dvss.t1392 202.299
R15089 dvss.t913 dvss.t1437 202.299
R15090 dvss.n3981 dvss.n3980 202.282
R15091 dvss.n4273 dvss.n4023 201.782
R15092 dvss.n2795 dvss.n2689 201.458
R15093 dvss.n2800 dvss.n2798 201.458
R15094 dvss.n3787 dvss.n3644 201.458
R15095 dvss.n3470 dvss.n3469 201.332
R15096 dvss.n226 dvss.t1521 201.177
R15097 dvss.n6392 dvss.t1082 201.177
R15098 dvss.n2786 dvss.n2692 201.129
R15099 dvss.n2789 dvss.n2787 201.129
R15100 dvss.n3777 dvss.n3647 201.129
R15101 dvss.n4017 dvss.n4016 201.129
R15102 dvss.t817 dvss.n3252 201.119
R15103 dvss.n2897 dvss.n2896 200.692
R15104 dvss.n3381 dvss.n3380 200.692
R15105 dvss.n3581 dvss.n3580 200.692
R15106 dvss.n4663 dvss.n4662 200.692
R15107 dvss.n4683 dvss.n4591 200.692
R15108 dvss.n3223 dvss.t537 200.689
R15109 dvss.n3634 dvss.n3633 200.516
R15110 dvss.n3981 dvss.n3979 200.516
R15111 dvss.n2844 dvss.n2805 200.508
R15112 dvss.n3769 dvss.n3768 200.508
R15113 dvss.n3801 dvss.n3799 200.508
R15114 dvss.n3336 dvss.t1037 200.25
R15115 dvss.n1593 dvss.n1578 200.215
R15116 dvss.n1593 dvss.n1592 200.215
R15117 dvss.n1878 dvss.n1877 200.215
R15118 dvss.n1879 dvss.n1878 200.215
R15119 dvss.n2030 dvss.n1439 200.215
R15120 dvss.n2033 dvss.n1439 200.215
R15121 dvss.n1006 dvss.n1005 200.215
R15122 dvss.n1006 dvss.n1001 200.215
R15123 dvss.n6133 dvss.n789 200.215
R15124 dvss.n6136 dvss.n789 200.215
R15125 dvss.n658 dvss.n608 200.215
R15126 dvss.n655 dvss.n608 200.215
R15127 dvss.n6874 dvss.n65 200.215
R15128 dvss.n6877 dvss.n65 200.215
R15129 dvss.n201 dvss.n200 200.215
R15130 dvss.n202 dvss.n201 200.215
R15131 dvss.n1772 dvss.n1771 200.215
R15132 dvss.n1773 dvss.n1772 200.215
R15133 dvss.n1888 dvss.n1887 200.215
R15134 dvss.n1889 dvss.n1888 200.215
R15135 dvss.n2043 dvss.n2042 200.215
R15136 dvss.n2044 dvss.n2043 200.215
R15137 dvss.n1011 dvss.n1010 200.215
R15138 dvss.n1012 dvss.n1011 200.215
R15139 dvss.n6146 dvss.n6145 200.215
R15140 dvss.n6147 dvss.n6146 200.215
R15141 dvss.n666 dvss.n665 200.215
R15142 dvss.n667 dvss.n666 200.215
R15143 dvss.n193 dvss.n192 200.215
R15144 dvss.n194 dvss.n193 200.215
R15145 dvss.n6887 dvss.n6886 200.215
R15146 dvss.n6888 dvss.n6887 200.215
R15147 dvss.n5670 dvss.n5668 200.215
R15148 dvss.n5668 dvss.n5667 200.215
R15149 dvss.n1059 dvss.n1058 200.215
R15150 dvss.n1060 dvss.n1059 200.215
R15151 dvss.n3336 dvss.n3335 200.215
R15152 dvss.n5495 dvss.n5494 200.215
R15153 dvss.n5495 dvss.n1154 200.215
R15154 dvss.n5495 dvss.n1155 200.215
R15155 dvss.n5495 dvss.n1156 200.215
R15156 dvss.n5495 dvss.n1157 200.215
R15157 dvss.n5495 dvss.n1158 200.215
R15158 dvss.n5495 dvss.n1159 200.215
R15159 dvss.n5495 dvss.n1160 200.215
R15160 dvss.n5495 dvss.n1161 200.215
R15161 dvss.n5495 dvss.n1162 200.215
R15162 dvss.n5495 dvss.n1163 200.215
R15163 dvss.n5495 dvss.n1164 200.215
R15164 dvss.n5495 dvss.n1165 200.215
R15165 dvss.n5495 dvss.n1166 200.215
R15166 dvss.n5495 dvss.n1167 200.215
R15167 dvss.n5495 dvss.n1168 200.215
R15168 dvss.n5495 dvss.n1169 200.215
R15169 dvss.n5495 dvss.n1170 200.215
R15170 dvss.n5495 dvss.n1171 200.215
R15171 dvss.n5495 dvss.n1172 200.215
R15172 dvss.n5495 dvss.n1173 200.215
R15173 dvss.n5495 dvss.n1174 200.215
R15174 dvss.n5495 dvss.n1175 200.215
R15175 dvss.n5495 dvss.n1176 200.215
R15176 dvss.n5495 dvss.n1177 200.215
R15177 dvss.n5495 dvss.n1178 200.215
R15178 dvss.n5495 dvss.n1179 200.215
R15179 dvss.n5495 dvss.n1180 200.215
R15180 dvss.n5495 dvss.n1181 200.215
R15181 dvss.n5495 dvss.n1182 200.215
R15182 dvss.n5495 dvss.n1183 200.215
R15183 dvss.n5495 dvss.n1184 200.215
R15184 dvss.n5495 dvss.n1185 200.215
R15185 dvss.n5495 dvss.n1186 200.215
R15186 dvss.n5495 dvss.n1187 200.215
R15187 dvss.n5495 dvss.n1188 200.215
R15188 dvss.n5495 dvss.n1189 200.215
R15189 dvss.n5495 dvss.n1190 200.215
R15190 dvss.n5495 dvss.n1191 200.215
R15191 dvss.n5495 dvss.n1192 200.215
R15192 dvss.n5495 dvss.n1193 200.215
R15193 dvss.n5495 dvss.n1194 200.215
R15194 dvss.n5495 dvss.n1195 200.215
R15195 dvss.n5495 dvss.n1196 200.215
R15196 dvss.n5495 dvss.n1197 200.215
R15197 dvss.n5495 dvss.n1198 200.215
R15198 dvss.n5495 dvss.n1199 200.215
R15199 dvss.n5495 dvss.n1200 200.215
R15200 dvss.n5495 dvss.n1201 200.215
R15201 dvss.n5495 dvss.n1202 200.215
R15202 dvss.n5495 dvss.n1203 200.215
R15203 dvss.n5495 dvss.n1204 200.215
R15204 dvss.n5496 dvss.n5495 200.215
R15205 dvss.n5495 dvss.n1205 200.215
R15206 dvss.n1730 dvss.n1729 200.215
R15207 dvss.n1730 dvss.n1625 200.215
R15208 dvss.n1730 dvss.n1626 200.215
R15209 dvss.n1730 dvss.n1627 200.215
R15210 dvss.n1731 dvss.n1730 200.215
R15211 dvss.n1755 dvss.n1754 200.215
R15212 dvss.n1755 dvss.n1573 200.215
R15213 dvss.n1755 dvss.n1574 200.215
R15214 dvss.n1755 dvss.n1575 200.215
R15215 dvss.n1755 dvss.n1576 200.215
R15216 dvss.n1648 dvss.n1647 200.215
R15217 dvss.n1648 dvss.n1645 200.215
R15218 dvss.n2004 dvss.n2003 200.215
R15219 dvss.n2004 dvss.n2001 200.215
R15220 dvss.n5738 dvss.n874 200.215
R15221 dvss.n5740 dvss.n874 200.215
R15222 dvss.n5834 dvss.n5833 200.215
R15223 dvss.n5835 dvss.n5834 200.215
R15224 dvss.n5922 dvss.n5921 200.215
R15225 dvss.n5922 dvss.n5920 200.215
R15226 dvss.n5996 dvss.n5995 200.215
R15227 dvss.n5996 dvss.n5993 200.215
R15228 dvss.n6728 dvss.n6727 200.215
R15229 dvss.n6729 dvss.n6728 200.215
R15230 dvss.n6810 dvss.n6809 200.215
R15231 dvss.n6810 dvss.n6808 200.215
R15232 dvss.n3468 dvss.n3467 200.127
R15233 dvss.n4405 dvss.n4300 200.127
R15234 dvss.n4552 dvss.n4551 200.127
R15235 dvss.n5010 dvss.n5009 200.127
R15236 dvss.n2684 dvss.n2682 200.105
R15237 dvss.n2708 dvss.n2707 199.966
R15238 dvss.n3682 dvss.n3661 199.966
R15239 dvss.n3877 dvss.n3853 199.966
R15240 dvss.n4421 dvss.n2399 199.966
R15241 dvss.n4098 dvss.n4043 199.966
R15242 dvss.n4159 dvss.n4158 199.966
R15243 dvss.n4542 dvss.n4541 199.923
R15244 dvss.n4550 dvss.n4549 199.917
R15245 dvss.n4557 dvss.n4556 199.917
R15246 dvss.n2528 dvss.n2432 199.739
R15247 dvss.n2927 dvss.n2926 199.739
R15248 dvss.n2995 dvss.n2994 199.739
R15249 dvss.n3106 dvss.n3059 199.739
R15250 dvss.n2780 dvss.n2779 199.739
R15251 dvss.n3716 dvss.n3708 199.739
R15252 dvss.n3722 dvss.n3706 199.739
R15253 dvss.n3722 dvss.n3721 199.739
R15254 dvss.n3737 dvss.n3735 199.739
R15255 dvss.n3737 dvss.n3736 199.739
R15256 dvss.n3899 dvss.n3841 199.739
R15257 dvss.n3844 dvss.n3843 199.739
R15258 dvss.n3884 dvss.n3848 199.739
R15259 dvss.n3852 dvss.n3851 199.739
R15260 dvss.n3922 dvss.n3921 199.739
R15261 dvss.n3932 dvss.n3923 199.739
R15262 dvss.n3937 dvss.n3920 199.739
R15263 dvss.n3945 dvss.n3944 199.739
R15264 dvss.n3953 dvss.n3952 199.739
R15265 dvss.n4335 dvss.n4334 199.739
R15266 dvss.n4399 dvss.n4304 199.739
R15267 dvss.n4623 dvss.n4622 199.739
R15268 dvss.n4631 dvss.n4630 199.739
R15269 dvss.n4896 dvss.n4895 199.739
R15270 dvss.n4901 dvss.n4900 199.739
R15271 dvss.n4906 dvss.n4905 199.739
R15272 dvss.n4911 dvss.n4910 199.739
R15273 dvss.n1223 dvss.n1222 199.739
R15274 dvss.n5075 dvss.n1227 199.739
R15275 dvss.n4125 dvss.n4031 199.739
R15276 dvss.n4175 dvss.n4148 199.739
R15277 dvss.n2797 dvss.n2688 199.662
R15278 dvss.n4037 dvss.n4036 199.417
R15279 dvss.n2389 dvss.n2388 199.131
R15280 dvss.n2824 dvss.n2817 199.052
R15281 dvss.n4333 dvss.n4332 199.052
R15282 dvss.n2731 dvss.n2710 198.986
R15283 dvss.n3657 dvss.n3656 198.986
R15284 dvss.n2384 dvss.n2383 198.986
R15285 dvss.n4285 dvss.n4015 198.986
R15286 dvss.n2529 dvss.n2431 198.964
R15287 dvss.n2813 dvss.n2812 198.964
R15288 dvss.n3683 dvss.n3660 198.964
R15289 dvss.n3677 dvss.n3663 198.964
R15290 dvss.n4227 dvss.n4216 198.654
R15291 dvss.n3004 dvss.n3002 198.577
R15292 dvss.n4611 dvss.n4610 197.535
R15293 dvss.n3616 dvss.n3510 197.288
R15294 dvss.n2419 dvss.n2418 197.219
R15295 dvss.n4230 dvss.n4213 197.219
R15296 dvss.n6339 dvss.t1446 197.171
R15297 dvss.n6266 dvss.t675 197.171
R15298 dvss.n4576 dvss.n4565 196.831
R15299 dvss.n4604 dvss.n4602 196.831
R15300 dvss.n3460 dvss.n3459 196.619
R15301 dvss.n2568 dvss.n2567 196.442
R15302 dvss.n2575 dvss.n2574 196.442
R15303 dvss.n2937 dvss.n2936 196.442
R15304 dvss.n2938 dvss.n2935 196.442
R15305 dvss.n2849 dvss.n2848 196.442
R15306 dvss.n3367 dvss.n3360 196.442
R15307 dvss.n2701 dvss.n2700 196.442
R15308 dvss.n3767 dvss.n3650 196.442
R15309 dvss.n3544 dvss.n3535 196.442
R15310 dvss.n3553 dvss.n3532 196.442
R15311 dvss.n4331 dvss.n4330 196.442
R15312 dvss.n4328 dvss.n4327 196.442
R15313 dvss.n4470 dvss.n2370 196.442
R15314 dvss.n2377 dvss.n2376 196.442
R15315 dvss.n4419 dvss.n2400 196.442
R15316 dvss.n4547 dvss.n4546 196.442
R15317 dvss.n4141 dvss.n4139 196.442
R15318 dvss.n4253 dvss.n4201 196.442
R15319 dvss.n4254 dvss.n4200 196.442
R15320 dvss.n4209 dvss.n4208 196.442
R15321 dvss.n4207 dvss.n4206 196.442
R15322 dvss.n4588 dvss.n4587 195.851
R15323 dvss.n2823 dvss.n2818 195.667
R15324 dvss.n4261 dvss.n4198 195.667
R15325 dvss.n4586 dvss.n4585 194.809
R15326 dvss.n7019 dvss.t295 194.704
R15327 dvss.t1403 dvss.t426 193.87
R15328 dvss.t95 dvss 193.87
R15329 dvss.t1581 dvss 193.87
R15330 dvss.t1042 dvss 193.87
R15331 dvss.t732 dvss 193.87
R15332 dvss.n3253 dvss.t817 192.911
R15333 dvss.n2895 dvss.n2894 190.399
R15334 dvss.n3355 dvss.n3351 190.399
R15335 dvss.n3579 dvss.n3578 190.399
R15336 dvss.n4609 dvss.n4607 190.399
R15337 dvss.n4685 dvss.n4684 190.399
R15338 dvss.n3064 dvss.n3063 190.237
R15339 dvss.n4310 dvss.n4309 189.4
R15340 dvss.n6981 dvss.n6980 188.91
R15341 dvss.n6860 dvss.n78 188.91
R15342 dvss.n5989 dvss.n5988 188.91
R15343 dvss.n6716 dvss.n120 188.91
R15344 dvss.n6119 dvss.n807 188.91
R15345 dvss.n5822 dvss.n5821 188.91
R15346 dvss.n5733 dvss.n5732 188.91
R15347 dvss.n2016 dvss.n1999 188.91
R15348 dvss.n1654 dvss.n1652 188.91
R15349 dvss.n4579 dvss.n4578 188.425
R15350 dvss.n6408 dvss.t1074 188.212
R15351 dvss.n6358 dvss.t1515 188.212
R15352 dvss.n2163 dvss.t2261 186.374
R15353 dvss.n880 dvss.t2291 186.374
R15354 dvss.n5812 dvss.t2287 186.374
R15355 dvss.n5896 dvss.t2243 186.374
R15356 dvss.n1400 dvss.t2292 186.374
R15357 dvss.n1449 dvss.t2262 186.374
R15358 dvss.n982 dvss.t2288 186.374
R15359 dvss.n799 dvss.t2244 186.374
R15360 dvss dvss.t120 185.441
R15361 dvss.t934 dvss.t1528 185.441
R15362 dvss.n3056 dvss.n3055 185
R15363 dvss.n3054 dvss.n3053 185
R15364 dvss.n3062 dvss.n3060 185
R15365 dvss.n3692 dvss.n3691 185
R15366 dvss.n3690 dvss.n3689 185
R15367 dvss.n3832 dvss.n3831 185
R15368 dvss.n3830 dvss.n3829 185
R15369 dvss.n4921 dvss.n4920 185
R15370 dvss.n4923 dvss.n4922 185
R15371 dvss.n1220 dvss.n1219 185
R15372 dvss.n5055 dvss.n5054 185
R15373 dvss.n5048 dvss.n5047 185
R15374 dvss.n5018 dvss.n5017 185
R15375 dvss.n4115 dvss.n4114 185
R15376 dvss.n4113 dvss.n4112 185
R15377 dvss.n1761 dvss.n1760 185
R15378 dvss.n5124 dvss.n5123 185
R15379 dvss.n5489 dvss.n1154 184.572
R15380 dvss.n5486 dvss.n1155 184.572
R15381 dvss.n5482 dvss.n1156 184.572
R15382 dvss.n5478 dvss.n1157 184.572
R15383 dvss.n5474 dvss.n1158 184.572
R15384 dvss.n5470 dvss.n1159 184.572
R15385 dvss.n5466 dvss.n1160 184.572
R15386 dvss.n5462 dvss.n1161 184.572
R15387 dvss.n5458 dvss.n1162 184.572
R15388 dvss.n5454 dvss.n1163 184.572
R15389 dvss.n5450 dvss.n1164 184.572
R15390 dvss.n5446 dvss.n1165 184.572
R15391 dvss.n5442 dvss.n1166 184.572
R15392 dvss.n5438 dvss.n1167 184.572
R15393 dvss.n5434 dvss.n1168 184.572
R15394 dvss.n5430 dvss.n1169 184.572
R15395 dvss.n5426 dvss.n1170 184.572
R15396 dvss.n5422 dvss.n1171 184.572
R15397 dvss.n5418 dvss.n1172 184.572
R15398 dvss.n5414 dvss.n1173 184.572
R15399 dvss.n5410 dvss.n1174 184.572
R15400 dvss.n5406 dvss.n1175 184.572
R15401 dvss.n5402 dvss.n1176 184.572
R15402 dvss.n5398 dvss.n1177 184.572
R15403 dvss.n5394 dvss.n1178 184.572
R15404 dvss.n5390 dvss.n1179 184.572
R15405 dvss.n5386 dvss.n1180 184.572
R15406 dvss.n5382 dvss.n1181 184.572
R15407 dvss.n5378 dvss.n1182 184.572
R15408 dvss.n5374 dvss.n1183 184.572
R15409 dvss.n5370 dvss.n1184 184.572
R15410 dvss.n5366 dvss.n1185 184.572
R15411 dvss.n5362 dvss.n1186 184.572
R15412 dvss.n5358 dvss.n1187 184.572
R15413 dvss.n5354 dvss.n1188 184.572
R15414 dvss.n5350 dvss.n1189 184.572
R15415 dvss.n5346 dvss.n1190 184.572
R15416 dvss.n5342 dvss.n1191 184.572
R15417 dvss.n5338 dvss.n1192 184.572
R15418 dvss.n5334 dvss.n1193 184.572
R15419 dvss.n5330 dvss.n1194 184.572
R15420 dvss.n5326 dvss.n1195 184.572
R15421 dvss.n5322 dvss.n1196 184.572
R15422 dvss.n5318 dvss.n1197 184.572
R15423 dvss.n5314 dvss.n1198 184.572
R15424 dvss.n5310 dvss.n1199 184.572
R15425 dvss.n5306 dvss.n1200 184.572
R15426 dvss.n5302 dvss.n1201 184.572
R15427 dvss.n5298 dvss.n1202 184.572
R15428 dvss.n5294 dvss.n1203 184.572
R15429 dvss.n5290 dvss.n1204 184.572
R15430 dvss.n5496 dvss.n1152 184.572
R15431 dvss.n1205 dvss.n1151 184.572
R15432 dvss.n1754 dvss.n1753 184.572
R15433 dvss.n1748 dvss.n1573 184.572
R15434 dvss.n1745 dvss.n1574 184.572
R15435 dvss.n1741 dvss.n1575 184.572
R15436 dvss.n1737 dvss.n1576 184.572
R15437 dvss.n1581 dvss.n1578 184.572
R15438 dvss.n1592 dvss.n1590 184.572
R15439 dvss.n1877 dvss.n1876 184.572
R15440 dvss.n1879 dvss.n1499 184.572
R15441 dvss.n2030 dvss.n1443 184.572
R15442 dvss.n2033 dvss.n2032 184.572
R15443 dvss.n1005 dvss.n1004 184.572
R15444 dvss.n1001 dvss.n1000 184.572
R15445 dvss.n1058 dvss.n1057 184.572
R15446 dvss.n1061 dvss.n1060 184.572
R15447 dvss.n6133 dvss.n793 184.572
R15448 dvss.n6136 dvss.n6135 184.572
R15449 dvss.n659 dvss.n658 184.572
R15450 dvss.n655 dvss.n654 184.572
R15451 dvss.n200 dvss.n199 184.572
R15452 dvss.n203 dvss.n202 184.572
R15453 dvss.n6874 dvss.n69 184.572
R15454 dvss.n6877 dvss.n6876 184.572
R15455 dvss.n1579 dvss.n1578 184.572
R15456 dvss.n1592 dvss.n1591 184.572
R15457 dvss.n1877 dvss.n1498 184.572
R15458 dvss.n1880 dvss.n1879 184.572
R15459 dvss.n2031 dvss.n2030 184.572
R15460 dvss.n2034 dvss.n2033 184.572
R15461 dvss.n1005 dvss.n1003 184.572
R15462 dvss.n1002 dvss.n1001 184.572
R15463 dvss.n6134 dvss.n6133 184.572
R15464 dvss.n6137 dvss.n6136 184.572
R15465 dvss.n658 dvss.n657 184.572
R15466 dvss.n656 dvss.n655 184.572
R15467 dvss.n6875 dvss.n6874 184.572
R15468 dvss.n6878 dvss.n6877 184.572
R15469 dvss.n200 dvss.n198 184.572
R15470 dvss.n202 dvss.n197 184.572
R15471 dvss.n1729 dvss.n1728 184.572
R15472 dvss.n1723 dvss.n1625 184.572
R15473 dvss.n1720 dvss.n1626 184.572
R15474 dvss.n1716 dvss.n1627 184.572
R15475 dvss.n1732 dvss.n1731 184.572
R15476 dvss.n1771 dvss.n1770 184.572
R15477 dvss.n1773 dvss.n1556 184.572
R15478 dvss.n1887 dvss.n1886 184.572
R15479 dvss.n1890 dvss.n1889 184.572
R15480 dvss.n2042 dvss.n2027 184.572
R15481 dvss.n2044 dvss.n1437 184.572
R15482 dvss.n1010 dvss.n1009 184.572
R15483 dvss.n1013 dvss.n1012 184.572
R15484 dvss.n5670 dvss.n5669 184.572
R15485 dvss.n5667 dvss.n5666 184.572
R15486 dvss.n6145 dvss.n6130 184.572
R15487 dvss.n6147 dvss.n787 184.572
R15488 dvss.n665 dvss.n664 184.572
R15489 dvss.n668 dvss.n667 184.572
R15490 dvss.n192 dvss.n191 184.572
R15491 dvss.n195 dvss.n194 184.572
R15492 dvss.n6886 dvss.n6871 184.572
R15493 dvss.n6888 dvss.n63 184.572
R15494 dvss.n1771 dvss.n1559 184.572
R15495 dvss.n1774 dvss.n1773 184.572
R15496 dvss.n1887 dvss.n1492 184.572
R15497 dvss.n1889 dvss.n1490 184.572
R15498 dvss.n2042 dvss.n2041 184.572
R15499 dvss.n2045 dvss.n2044 184.572
R15500 dvss.n1010 dvss.n901 184.572
R15501 dvss.n1012 dvss.n902 184.572
R15502 dvss.n6145 dvss.n6144 184.572
R15503 dvss.n6148 dvss.n6147 184.572
R15504 dvss.n665 dvss.n547 184.572
R15505 dvss.n667 dvss.n548 184.572
R15506 dvss.n192 dvss.n135 184.572
R15507 dvss.n194 dvss.n136 184.572
R15508 dvss.n6886 dvss.n6885 184.572
R15509 dvss.n6889 dvss.n6888 184.572
R15510 dvss.n5671 dvss.n5670 184.572
R15511 dvss.n5667 dvss.n952 184.572
R15512 dvss.n1058 dvss.n973 184.572
R15513 dvss.n1060 dvss.n970 184.572
R15514 dvss.n3335 dvss.n3127 184.572
R15515 dvss.n5494 dvss.n1207 184.572
R15516 dvss.n5487 dvss.n1154 184.572
R15517 dvss.n5483 dvss.n1155 184.572
R15518 dvss.n5479 dvss.n1156 184.572
R15519 dvss.n5475 dvss.n1157 184.572
R15520 dvss.n5471 dvss.n1158 184.572
R15521 dvss.n5467 dvss.n1159 184.572
R15522 dvss.n5463 dvss.n1160 184.572
R15523 dvss.n5459 dvss.n1161 184.572
R15524 dvss.n5455 dvss.n1162 184.572
R15525 dvss.n5451 dvss.n1163 184.572
R15526 dvss.n5447 dvss.n1164 184.572
R15527 dvss.n5443 dvss.n1165 184.572
R15528 dvss.n5439 dvss.n1166 184.572
R15529 dvss.n5435 dvss.n1167 184.572
R15530 dvss.n5431 dvss.n1168 184.572
R15531 dvss.n5427 dvss.n1169 184.572
R15532 dvss.n5423 dvss.n1170 184.572
R15533 dvss.n5419 dvss.n1171 184.572
R15534 dvss.n5415 dvss.n1172 184.572
R15535 dvss.n5411 dvss.n1173 184.572
R15536 dvss.n5407 dvss.n1174 184.572
R15537 dvss.n5403 dvss.n1175 184.572
R15538 dvss.n5399 dvss.n1176 184.572
R15539 dvss.n5395 dvss.n1177 184.572
R15540 dvss.n5391 dvss.n1178 184.572
R15541 dvss.n5387 dvss.n1179 184.572
R15542 dvss.n5383 dvss.n1180 184.572
R15543 dvss.n5379 dvss.n1181 184.572
R15544 dvss.n5375 dvss.n1182 184.572
R15545 dvss.n5371 dvss.n1183 184.572
R15546 dvss.n5367 dvss.n1184 184.572
R15547 dvss.n5363 dvss.n1185 184.572
R15548 dvss.n5359 dvss.n1186 184.572
R15549 dvss.n5355 dvss.n1187 184.572
R15550 dvss.n5351 dvss.n1188 184.572
R15551 dvss.n5347 dvss.n1189 184.572
R15552 dvss.n5343 dvss.n1190 184.572
R15553 dvss.n5339 dvss.n1191 184.572
R15554 dvss.n5335 dvss.n1192 184.572
R15555 dvss.n5331 dvss.n1193 184.572
R15556 dvss.n5327 dvss.n1194 184.572
R15557 dvss.n5323 dvss.n1195 184.572
R15558 dvss.n5319 dvss.n1196 184.572
R15559 dvss.n5315 dvss.n1197 184.572
R15560 dvss.n5311 dvss.n1198 184.572
R15561 dvss.n5307 dvss.n1199 184.572
R15562 dvss.n5303 dvss.n1200 184.572
R15563 dvss.n5299 dvss.n1201 184.572
R15564 dvss.n5295 dvss.n1202 184.572
R15565 dvss.n5291 dvss.n1203 184.572
R15566 dvss.n5287 dvss.n1204 184.572
R15567 dvss.n5497 dvss.n5496 184.572
R15568 dvss.n1205 dvss.n1146 184.572
R15569 dvss.n1729 dvss.n1689 184.572
R15570 dvss.n1721 dvss.n1625 184.572
R15571 dvss.n1717 dvss.n1626 184.572
R15572 dvss.n1627 dvss.n1623 184.572
R15573 dvss.n1731 dvss.n1624 184.572
R15574 dvss.n1754 dvss.n1596 184.572
R15575 dvss.n1746 dvss.n1573 184.572
R15576 dvss.n1742 dvss.n1574 184.572
R15577 dvss.n1738 dvss.n1575 184.572
R15578 dvss.n1576 dvss.n1568 184.572
R15579 dvss.n1647 dvss.n1646 184.572
R15580 dvss.n1645 dvss.n1290 184.572
R15581 dvss.n2003 dvss.n2002 184.572
R15582 dvss.n2001 dvss.n1321 184.572
R15583 dvss.n5738 dvss.n877 184.572
R15584 dvss.n5741 dvss.n5740 184.572
R15585 dvss.n5833 dvss.n5832 184.572
R15586 dvss.n5836 dvss.n5835 184.572
R15587 dvss.n5921 dvss.n5902 184.572
R15588 dvss.n5920 dvss.n5919 184.572
R15589 dvss.n5995 dvss.n5994 184.572
R15590 dvss.n5993 dvss.n5951 184.572
R15591 dvss.n6727 dvss.n6726 184.572
R15592 dvss.n6730 dvss.n6729 184.572
R15593 dvss.n6809 dvss.n6791 184.572
R15594 dvss.n6808 dvss.n6807 184.572
R15595 dvss.n6986 dvss.n6985 184.572
R15596 dvss.n1647 dvss.n1289 184.572
R15597 dvss.n1645 dvss.n1644 184.572
R15598 dvss.n2003 dvss.n1320 184.572
R15599 dvss.n2001 dvss.n2000 184.572
R15600 dvss.n5739 dvss.n5738 184.572
R15601 dvss.n5740 dvss.n873 184.572
R15602 dvss.n5833 dvss.n844 184.572
R15603 dvss.n5835 dvss.n841 184.572
R15604 dvss.n5921 dvss.n5903 184.572
R15605 dvss.n5920 dvss.n5905 184.572
R15606 dvss.n5995 dvss.n5950 184.572
R15607 dvss.n5993 dvss.n5992 184.572
R15608 dvss.n6727 dvss.n115 184.572
R15609 dvss.n6729 dvss.n112 184.572
R15610 dvss.n6809 dvss.n6792 184.572
R15611 dvss.n6808 dvss.n6794 184.572
R15612 dvss.n6293 dvss.t1481 178.282
R15613 dvss.t1376 dvss.n6221 178.282
R15614 dvss.t2060 dvss.t2028 177.012
R15615 dvss.t1551 dvss.t617 177.012
R15616 dvss.t36 dvss.t892 177.012
R15617 dvss.t1046 dvss.t317 177.012
R15618 dvss.t1288 dvss.t2130 177.012
R15619 dvss.t183 dvss.t1176 177.012
R15620 dvss.t1283 dvss.t919 177.012
R15621 dvss.n6460 dvss.t1064 172.957
R15622 dvss.n6652 dvss.t907 172.957
R15623 dvss.n694 dvss.t1563 172.957
R15624 dvss.n633 dvss.t1364 172.957
R15625 dvss.t486 dvss.n5616 172.957
R15626 dvss.t2163 dvss.n1039 172.957
R15627 dvss.n1381 dvss.t613 172.957
R15628 dvss.n1955 dvss.t281 172.957
R15629 dvss.t113 dvss.n1848 172.957
R15630 dvss.t1653 dvss.t1662 172.464
R15631 dvss.t1662 dvss.t1593 172.464
R15632 dvss.t1593 dvss.t1623 172.464
R15633 dvss.t1671 dvss.t1596 172.464
R15634 dvss.t1596 dvss.t1629 172.464
R15635 dvss.t1629 dvss.t1680 172.464
R15636 dvss.t1429 dvss.n6901 171.311
R15637 dvss.n671 dvss.t1973 171.311
R15638 dvss.t1986 dvss.n6160 171.311
R15639 dvss.n1016 dvss.t311 171.311
R15640 dvss.t357 dvss.n2057 171.311
R15641 dvss.n1901 dvss.t132 171.311
R15642 dvss.n1792 dvss.t297 171.311
R15643 dvss.n207 dvss.t2058 171.311
R15644 dvss.n5661 dvss.t478 171.311
R15645 dvss.n2163 dvss.t1631 170.308
R15646 dvss.n880 dvss.t1607 170.308
R15647 dvss.n5812 dvss.t1610 170.308
R15648 dvss.n5896 dvss.t1655 170.308
R15649 dvss.n1400 dvss.t1586 170.308
R15650 dvss.n1449 dvss.t1601 170.308
R15651 dvss.n982 dvss.t1589 170.308
R15652 dvss.n799 dvss.t1613 170.308
R15653 dvss.n6358 dvss.t1513 169.85
R15654 dvss.t1072 dvss.n6408 169.85
R15655 dvss.t217 dvss.n6471 169.498
R15656 dvss.n6655 dvss.t1301 169.498
R15657 dvss.t2109 dvss.n698 169.498
R15658 dvss.n632 dvss.t2096 169.498
R15659 dvss.n5618 dvss.t1614 169.498
R15660 dvss.n1040 dvss.t1590 169.498
R15661 dvss.t1587 dvss.n1392 169.498
R15662 dvss.n1958 dvss.t1602 169.498
R15663 dvss.t2142 dvss.n1849 169.498
R15664 dvss.t444 dvss.t2103 168.583
R15665 dvss.t140 dvss.t392 168.583
R15666 dvss.t1549 dvss.t384 168.583
R15667 dvss.t1052 dvss 168.583
R15668 dvss.t2191 dvss.t1966 168.583
R15669 dvss.t173 dvss.t1261 168.583
R15670 dvss.n4193 dvss.t1051 168.583
R15671 dvss.t130 dvss.n1679 167.899
R15672 dvss.n5861 dvss.t663 166.838
R15673 dvss.n6755 dvss.t1414 166.838
R15674 dvss.n6818 dvss.t1103 166.838
R15675 dvss.n5931 dvss.t2203 166.838
R15676 dvss.n6004 dvss.t1005 166.838
R15677 dvss.t1113 dvss.n5768 166.838
R15678 dvss.t1490 dvss.n2008 166.838
R15679 dvss.t1311 dvss.n1637 166.838
R15680 dvss.t263 dvss.n1665 166.838
R15681 dvss.n6542 dvss.t660 166.689
R15682 dvss.t1481 dvss.n477 164.019
R15683 dvss.n6224 dvss.t1376 164.019
R15684 dvss.n3236 dvss.t537 162.823
R15685 dvss.n6472 dvss.t217 162.579
R15686 dvss.n6658 dvss.t1301 162.579
R15687 dvss.n699 dvss.t2109 162.579
R15688 dvss.n647 dvss.t2096 162.579
R15689 dvss.n5621 dvss.t1614 162.579
R15690 dvss.n1047 dvss.t1590 162.579
R15691 dvss.n1393 dvss.t1587 162.579
R15692 dvss.n1961 dvss.t1602 162.579
R15693 dvss.n1853 dvss.t2142 162.579
R15694 dvss.n4034 dvss.t174 162.471
R15695 dvss.n3215 dvss 161.882
R15696 dvss.n6920 dvss 161.882
R15697 dvss.n6692 dvss 161.882
R15698 dvss.n736 dvss 161.882
R15699 dvss.n6179 dvss 161.882
R15700 dvss.n1087 dvss 161.882
R15701 dvss.n5708 dvss 161.882
R15702 dvss.n2076 dvss 161.882
R15703 dvss.n1478 dvss 161.882
R15704 dvss.n1544 dvss 161.882
R15705 dvss.n6803 dvss 161.882
R15706 dvss.n6748 dvss 161.882
R15707 dvss.n5961 dvss 161.882
R15708 dvss.n5914 dvss 161.882
R15709 dvss.n5854 dvss 161.882
R15710 dvss.n865 dvss 161.882
R15711 dvss.n1331 dvss 161.882
R15712 dvss.n1300 dvss 161.882
R15713 dvss.n1269 dvss 161.882
R15714 dvss.t1105 dvss.n6816 161.857
R15715 dvss.n6741 dvss.t1412 161.857
R15716 dvss.t2205 dvss.n5928 161.857
R15717 dvss.t1001 dvss.n6001 161.857
R15718 dvss.n5847 dvss.t671 161.857
R15719 dvss.t1117 dvss.n5767 161.857
R15720 dvss.n2010 dvss.t1492 161.857
R15721 dvss.n1641 dvss.t1313 161.857
R15722 dvss.n1666 dvss.t265 161.857
R15723 dvss.n289 dvss.t63 161.522
R15724 dvss.n257 dvss.t1139 161.522
R15725 dvss.n4819 dvss.n2300 161.506
R15726 dvss.n395 dvss.t228 161.47
R15727 dvss.n3326 dvss.n3325 161.345
R15728 dvss.n3325 dvss.n3324 161.345
R15729 dvss.n3324 dvss.n3137 161.345
R15730 dvss.n3318 dvss.n3137 161.345
R15731 dvss.n3318 dvss.n3317 161.345
R15732 dvss.n3317 dvss.n3316 161.345
R15733 dvss.n3316 dvss.n3145 161.345
R15734 dvss.n3309 dvss.n3308 161.345
R15735 dvss.n3299 dvss.n3266 161.345
R15736 dvss.n3293 dvss.n3266 161.345
R15737 dvss.n3293 dvss.n3292 161.345
R15738 dvss.n3292 dvss.n3291 161.345
R15739 dvss.n345 dvss.t335 161.143
R15740 dvss.n2951 dvss.t556 160.8
R15741 dvss.t1016 dvss 160.154
R15742 dvss.t645 dvss 160.154
R15743 dvss.t970 dvss.t968 160.154
R15744 dvss dvss.t744 160.154
R15745 dvss dvss.t1454 160.154
R15746 dvss.t990 dvss.t1263 160.154
R15747 dvss.t463 dvss.t197 160.154
R15748 dvss.n1614 dvss.t1026 160.064
R15749 dvss.n1250 dvss.t125 160.064
R15750 dvss.n4122 dvss.t172 160.017
R15751 dvss.n4620 dvss.t1357 157.291
R15752 dvss.n1686 dvss.n1630 157.238
R15753 dvss.n3511 dvss.t2068 156.915
R15754 dvss.n5571 dvss.n5564 155.566
R15755 dvss.n4637 dvss.t1355 155.286
R15756 dvss.t1070 dvss.n6967 154.8
R15757 dvss.n6771 dvss.t905 154.8
R15758 dvss.n5981 dvss.t1366 154.8
R15759 dvss.n6011 dvss.t1557 154.8
R15760 dvss.n5877 dvss.t480 154.8
R15761 dvss.t2157 dvss.n5800 154.8
R15762 dvss.t605 dvss.n2111 154.8
R15763 dvss.n1992 dvss.t271 154.8
R15764 dvss.n1660 dvss.t115 154.8
R15765 dvss.n2726 dvss.t2047 154.746
R15766 dvss.n4024 dvss.t103 154.725
R15767 dvss.n2429 dvss.t2148 154.561
R15768 dvss.n3928 dvss.t835 154.561
R15769 dvss.n3536 dvss.t1192 154.561
R15770 dvss.n3531 dvss.t546 154.561
R15771 dvss.n4341 dvss.t2077 154.561
R15772 dvss.n4629 dvss.t2229 154.561
R15773 dvss.n5001 dvss.t1976 154.561
R15774 dvss.n4988 dvss.t1486 154.561
R15775 dvss.n4975 dvss.t753 154.561
R15776 dvss.n4962 dvss.t2088 154.561
R15777 dvss.n5081 dvss.t1360 154.561
R15778 dvss.n1225 dvss.t967 154.561
R15779 dvss.n2164 dvss 154.56
R15780 dvss.n881 dvss 154.56
R15781 dvss.n5813 dvss 154.56
R15782 dvss.n5897 dvss 154.56
R15783 dvss.n1401 dvss 154.56
R15784 dvss.n1450 dvss 154.56
R15785 dvss.n983 dvss 154.56
R15786 dvss.n800 dvss 154.56
R15787 dvss.n1710 dvss.t1258 154.305
R15788 dvss.n2279 dvss.t1036 154.305
R15789 dvss.n4736 dvss.t1499 154.129
R15790 dvss.n2165 dvss.n2164 153.462
R15791 dvss.n882 dvss.n881 153.462
R15792 dvss.n5814 dvss.n5813 153.462
R15793 dvss.n5898 dvss.n5897 153.462
R15794 dvss.n1402 dvss.n1401 153.462
R15795 dvss.n1451 dvss.n1450 153.462
R15796 dvss.n984 dvss.n983 153.462
R15797 dvss.n801 dvss.n800 153.462
R15798 dvss.t1650 dvss.t2098 153.21
R15799 dvss.n310 dvss.t61 152.838
R15800 dvss.n384 dvss.t258 152.838
R15801 dvss.n246 dvss.t1137 152.838
R15802 dvss.n371 dvss.t353 152.838
R15803 dvss.n3611 dvss.t865 152.466
R15804 dvss.n2896 dvss.n2876 152
R15805 dvss.n3382 dvss.n3381 152
R15806 dvss.n3580 dvss.n3522 152
R15807 dvss.n4683 dvss.n4682 152
R15808 dvss.n4664 dvss.n4663 152
R15809 dvss.n3252 dvss.t1466 151.867
R15810 dvss.t1444 dvss.t619 151.725
R15811 dvss.t984 dvss.t700 151.725
R15812 dvss.t494 dvss.t476 151.725
R15813 dvss.t1918 dvss.t1330 151.725
R15814 dvss.t693 dvss.t31 151.725
R15815 dvss.t168 dvss.t181 151.725
R15816 dvss dvss.t20 151.725
R15817 dvss.t1279 dvss.t213 151.725
R15818 dvss.n2642 dvss.t2104 150.922
R15819 dvss.n2732 dvss.t1335 150.922
R15820 dvss.n2737 dvss.t1961 150.922
R15821 dvss.n4092 dvss.t86 150.922
R15822 dvss.n4654 dvss.t3 150.376
R15823 dvss.n2730 dvss.t96 150.101
R15824 dvss.n3992 dvss.t461 149.493
R15825 dvss.n3429 dvss.t873 149.493
R15826 dvss.n3897 dvss.t2174 149.493
R15827 dvss.n3035 dvss.t2106 149.395
R15828 dvss.n6948 dvss.t1233 148.743
R15829 dvss.t1130 dvss.n225 148.743
R15830 dvss.n688 dvss.t361 148.743
R15831 dvss.n6207 dvss.t780 148.743
R15832 dvss.t1293 dvss.n1121 148.743
R15833 dvss.n1033 dvss.t6 148.743
R15834 dvss.n2104 dvss.t1340 148.743
R15835 dvss.n1469 dvss.t973 148.743
R15836 dvss.t2214 dvss.n1538 148.743
R15837 dvss.n2838 dvss.t1172 147.411
R15838 dvss.n3406 dvss.t2182 147.411
R15839 dvss.n432 dvss.n431 146.25
R15840 dvss.n433 dvss.n432 146.25
R15841 dvss.n420 dvss.n419 146.25
R15842 dvss.n419 dvss.n335 146.25
R15843 dvss.n4400 dvss.t2170 144.886
R15844 dvss.n3310 dvss.t1462 144.538
R15845 dvss.n227 dvss.t1517 143.697
R15846 dvss.n6519 dvss.t1076 143.697
R15847 dvss dvss.t1904 143.296
R15848 dvss dvss.t1691 143.296
R15849 dvss.n4049 dvss 143.296
R15850 dvss dvss.t1685 143.296
R15851 dvss.n4593 dvss 143.296
R15852 dvss.n4418 dvss.t1438 141.135
R15853 dvss.n3302 dvss.n3301 140.614
R15854 dvss.n3237 dvss.n3236 140.103
R15855 dvss.t1229 dvss.n48 139.755
R15856 dvss.n675 dvss.t359 139.755
R15857 dvss.t784 dvss.n772 139.755
R15858 dvss.n1020 dvss.t12 139.755
R15859 dvss.t1346 dvss.n1422 139.755
R15860 dvss.n1914 dvss.t979 139.755
R15861 dvss.n1797 dvss.t2220 139.755
R15862 dvss.t1124 dvss.n185 139.755
R15863 dvss.n5655 dvss.t1299 139.755
R15864 dvss.n1609 dvss.t401 139.52
R15865 dvss.n5113 dvss.t760 139.52
R15866 dvss.t1099 dvss.n23 139.059
R15867 dvss.n6756 dvss.t1408 139.059
R15868 dvss.n5933 dvss.t2201 139.059
R15869 dvss.t1003 dvss.n6006 139.059
R15870 dvss.n5862 dvss.t665 139.059
R15871 dvss.t1121 dvss.n5786 139.059
R15872 dvss.t1496 dvss.n1347 139.059
R15873 dvss.t1307 dvss.n1987 139.059
R15874 dvss.t259 dvss.n1635 139.059
R15875 dvss.n1614 dvss.t1028 137.442
R15876 dvss.n1615 dvss.t1031 137.442
R15877 dvss.n1250 dvss.t127 137.442
R15878 dvss.n1251 dvss.t131 137.442
R15879 dvss.t1760 dvss.t1399 134.867
R15880 dvss.t1213 dvss.t639 134.867
R15881 dvss.t637 dvss.t738 134.867
R15882 dvss.t704 dvss.t595 134.867
R15883 dvss.t118 dvss.t34 134.867
R15884 dvss.t381 dvss.t2013 134.867
R15885 dvss dvss.t2119 134.867
R15886 dvss.n44 dvss.t1233 134.488
R15887 dvss.t1130 dvss.n183 134.488
R15888 dvss.n684 dvss.t361 134.488
R15889 dvss.n768 dvss.t780 134.488
R15890 dvss.t1293 dvss.n1120 134.488
R15891 dvss.n1029 dvss.t6 134.488
R15892 dvss.n1418 dvss.t1340 134.488
R15893 dvss.n1471 dvss.t973 134.488
R15894 dvss.n1819 dvss.t2214 134.488
R15895 dvss.n6640 dvss.t1517 132.202
R15896 dvss.t1227 dvss.n6926 130.738
R15897 dvss.n678 dvss.t363 130.738
R15898 dvss.t782 dvss.n6185 130.738
R15899 dvss.n1023 dvss.t8 130.738
R15900 dvss.t1344 dvss.n2082 130.738
R15901 dvss.n1915 dvss.t977 130.738
R15902 dvss.n1796 dvss.t2218 130.738
R15903 dvss.t1126 dvss.n216 130.738
R15904 dvss.n5654 dvss.t1291 130.738
R15905 dvss.n4850 dvss.n1232 129.882
R15906 dvss.t1326 dvss.n6968 128.564
R15907 dvss.t2023 dvss.n6784 128.564
R15908 dvss.t2107 dvss.n5984 128.564
R15909 dvss.t1533 dvss.n6014 128.564
R15910 dvss.t1656 dvss.n5890 128.564
R15911 dvss.n5801 dvss.t1611 128.564
R15912 dvss.t1608 dvss.n2112 128.564
R15913 dvss.t1632 dvss.n1995 128.564
R15914 dvss.n1657 dvss.t1023 128.564
R15915 dvss.n6471 dvss.t1080 127.987
R15916 dvss.n6655 dvss.t1523 127.987
R15917 dvss.n698 dvss.t1483 127.987
R15918 dvss.t1384 dvss.n632 127.987
R15919 dvss.n5618 dvss.t1541 127.987
R15920 dvss.n1040 dvss.t2053 127.987
R15921 dvss.n1392 dvss.t514 127.987
R15922 dvss.n1958 dvss.t682 127.987
R15923 dvss.n1849 dvss.t44 127.987
R15924 dvss.t1390 dvss.t1262 126.438
R15925 dvss.t1424 dvss.t2155 126.438
R15926 dvss.n6949 dvss.t1082 125.389
R15927 dvss.n6647 dvss.t1521 125.389
R15928 dvss.n3153 dvss.t1458 125.389
R15929 dvss.n5610 dvss.t1543 125.389
R15930 dvss.n6969 dvss.t1326 123.316
R15931 dvss.n6785 dvss.t2023 123.316
R15932 dvss.n5985 dvss.t2107 123.316
R15933 dvss.n6015 dvss.t1533 123.316
R15934 dvss.n5891 dvss.t1656 123.316
R15935 dvss.t1611 dvss.n850 123.316
R15936 dvss.n2113 dvss.t1608 123.316
R15937 dvss.n1996 dvss.t1632 123.316
R15938 dvss.t1023 dvss.n1656 123.316
R15939 dvss.n5022 dvss.t2236 121.927
R15940 dvss.n4083 dvss.t2242 121.927
R15941 dvss.n4702 dvss.n4579 121.6
R15942 dvss.n3998 dvss.n3454 121.451
R15943 dvss.t1460 dvss.n3300 120.108
R15944 dvss.t1269 dvss.t589 118.008
R15945 dvss.t1526 dvss.t636 118.008
R15946 dvss.t146 dvss.t430 118.008
R15947 dvss.t1971 dvss.t1418 118.008
R15948 dvss.n4106 dvss.n4039 117.889
R15949 dvss.n3310 dvss.t1458 117.647
R15950 dvss.t533 dvss.n3185 117.385
R15951 dvss.n3281 dvss.t1457 116.939
R15952 dvss.n6485 dvss.t1061 116.939
R15953 dvss.n6867 dvss.t902 116.939
R15954 dvss.n708 dvss.t1554 116.939
R15955 dvss.n757 dvss.t1371 116.939
R15956 dvss.n6126 dvss.t491 116.939
R15957 dvss.n5680 dvss.t2162 116.939
R15958 dvss.n1407 dvss.t612 116.939
R15959 dvss.n2023 dvss.t276 116.939
R15960 dvss.n1864 dvss.t112 116.939
R15961 dvss.n6423 dvss.t1073 116.939
R15962 dvss.n6557 dvss.t1514 116.939
R15963 dvss.n6301 dvss.t1474 116.939
R15964 dvss.n6233 dvss.t1381 116.939
R15965 dvss.n5537 dvss.t1546 116.939
R15966 dvss.n5280 dvss.t2051 116.939
R15967 dvss.n5241 dvss.t512 116.939
R15968 dvss.n5202 dvss.t680 116.939
R15969 dvss.n5163 dvss.t46 116.939
R15970 dvss.n3231 dvss.t538 116.938
R15971 dvss.n6937 dvss.t1234 116.938
R15972 dvss.n6683 dvss.t1131 116.938
R15973 dvss.n727 dvss.t362 116.938
R15974 dvss.n6196 dvss.t781 116.938
R15975 dvss.n1099 dvss.t1294 116.938
R15976 dvss.n5699 dvss.t7 116.938
R15977 dvss.n2093 dvss.t1341 116.938
R15978 dvss.n1940 dvss.t974 116.938
R15979 dvss.n1828 dvss.t2215 116.938
R15980 dvss.n6826 dvss.t1100 116.938
R15981 dvss.n6764 dvss.t1409 116.938
R15982 dvss.n6035 dvss.t1004 116.938
R15983 dvss.n6085 dvss.t2202 116.938
R15984 dvss.n5870 dvss.t666 116.938
R15985 dvss.n5792 dvss.t1122 116.938
R15986 dvss.n2129 dvss.t1497 116.938
R15987 dvss.n2184 dvss.t1308 116.938
R15988 dvss.n2234 dvss.t260 116.938
R15989 dvss.n4617 dvss.t2296 116.734
R15990 dvss.t40 dvss.n862 116.547
R15991 dvss.n2105 dvss.t40 116.547
R15992 dvss.n1985 dvss.t40 116.547
R15993 dvss.n1530 dvss.t40 116.547
R15994 dvss.n3013 dvss.n3011 114.377
R15995 dvss.n3529 dvss.n3528 114.376
R15996 dvss dvss.n3170 113.316
R15997 dvss dvss.n6449 113.316
R15998 dvss dvss.n174 113.316
R15999 dvss dvss.n583 113.316
R16000 dvss dvss.n622 113.316
R16001 dvss dvss.n1107 113.316
R16002 dvss dvss.n937 113.316
R16003 dvss dvss.n1371 113.316
R16004 dvss dvss.n1947 113.316
R16005 dvss dvss.n1841 113.316
R16006 dvss dvss.n6957 113.316
R16007 dvss dvss.n88 113.316
R16008 dvss dvss.n5972 113.316
R16009 dvss dvss.n5941 113.316
R16010 dvss dvss.n817 113.316
R16011 dvss dvss.n854 113.316
R16012 dvss dvss.n1342 113.316
R16013 dvss dvss.n1311 113.316
R16014 dvss dvss.n1280 113.316
R16015 dvss.n6950 dvss.t1099 112.822
R16016 dvss.n6769 dvss.t1408 112.822
R16017 dvss.n5978 dvss.t2201 112.822
R16018 dvss.n6008 dvss.t1003 112.822
R16019 dvss.n5875 dvss.t665 112.822
R16020 dvss.n5787 dvss.t1121 112.822
R16021 dvss.n2107 dvss.t1496 112.822
R16022 dvss.n1989 dvss.t1307 112.822
R16023 dvss.t259 dvss.n1664 112.822
R16024 dvss.n3515 dvss.t2311 112.349
R16025 dvss.n4567 dvss.n4566 111.15
R16026 dvss.n5068 dvss.n5006 111.15
R16027 dvss.t531 dvss.n3221 109.811
R16028 dvss dvss.t569 109.579
R16029 dvss.t1977 dvss.t144 109.579
R16030 dvss.t1174 dvss.t890 109.579
R16031 dvss.t1094 dvss.t1091 109.579
R16032 dvss.t915 dvss 109.579
R16033 dvss.t20 dvss.t1420 109.579
R16034 dvss.n4315 dvss.t2040 109.579
R16035 dvss.n6383 dvss.t660 109.21
R16036 dvss.n3011 dvss.t1575 108.505
R16037 dvss.n3528 dvss.t2033 108.505
R16038 dvss.n3300 dvss.t1456 108.389
R16039 dvss.n4670 dvss.n4605 107.853
R16040 dvss.n1766 dvss.n1565 105.862
R16041 dvss.n2264 dvss.n1255 105.862
R16042 dvss.t1076 dvss.n6518 105.582
R16043 dvss.n4495 dvss.t2326 102.353
R16044 dvss.n2164 dvss.n2163 101.513
R16045 dvss.n881 dvss.n880 101.513
R16046 dvss.n5813 dvss.n5812 101.513
R16047 dvss.n5897 dvss.n5896 101.513
R16048 dvss.n1401 dvss.n1400 101.513
R16049 dvss.n1450 dvss.n1449 101.513
R16050 dvss.n983 dvss.n982 101.513
R16051 dvss.n800 dvss.n799 101.513
R16052 dvss.n2535 dvss.t871 101.43
R16053 dvss.n2674 dvss.t2176 101.43
R16054 dvss.n3471 dvss.t884 101.43
R16055 dvss.n3465 dvss.t39 101.43
R16056 dvss.n3525 dvss.t2031 101.43
R16057 dvss.n4914 dvss.t2125 101.43
R16058 dvss.t561 dvss.t748 101.15
R16059 dvss.t941 dvss.t993 101.15
R16060 dvss.t642 dvss.t452 101.15
R16061 dvss.t456 dvss.t1581 101.15
R16062 dvss dvss.t170 101.15
R16063 dvss.t850 dvss.t859 101.15
R16064 dvss.n2425 dvss.t429 100.001
R16065 dvss.n2931 dvss.t415 100.001
R16066 dvss.n2922 dvss.t413 100.001
R16067 dvss.n2851 dvss.t427 100.001
R16068 dvss.n2754 dvss.t959 100.001
R16069 dvss.n3745 dvss.t961 100.001
R16070 dvss.n3746 dvss.t409 100.001
R16071 dvss.n3778 dvss.t443 100.001
R16072 dvss.n3833 dvss.t421 100.001
R16073 dvss.n3856 dvss.t417 100.001
R16074 dvss.n3955 dvss.t1419 100.001
R16075 dvss.n3912 dvss.t405 100.001
R16076 dvss.n2366 dvss.t947 100.001
R16077 dvss.n2396 dvss.t963 100.001
R16078 dvss.n4028 dvss.t951 100.001
R16079 dvss.n4099 dvss.t955 100.001
R16080 dvss.n4195 dvss.t433 100.001
R16081 dvss.n4214 dvss.t1425 100.001
R16082 dvss.n3003 dvss.t727 99.9005
R16083 dvss.n2501 dvss.t2271 99.7825
R16084 dvss.n1686 dvss.n1685 98.6074
R16085 dvss.n3265 dvss.n3264 98.508
R16086 dvss.n2299 dvss.n2297 97.5005
R16087 dvss.n4808 dvss.n2297 97.5005
R16088 dvss.n4810 dvss.n4809 97.5005
R16089 dvss.n4811 dvss.n4810 97.5005
R16090 dvss.n4821 dvss.n4820 97.5005
R16091 dvss.n4822 dvss.n4821 97.5005
R16092 dvss.n2300 dvss.n2298 97.5005
R16093 dvss.n4808 dvss.n2298 97.5005
R16094 dvss.n4801 dvss.n4800 97.5005
R16095 dvss.n4800 dvss.n4799 97.5005
R16096 dvss.n4804 dvss.n4803 97.5005
R16097 dvss.n4805 dvss.n4804 97.5005
R16098 dvss.n4855 dvss.n4854 97.5005
R16099 dvss.n4856 dvss.n4855 97.5005
R16100 dvss.n4852 dvss.n4851 97.5005
R16101 dvss.n4851 dvss.n1153 97.5005
R16102 dvss.t2224 dvss.n3136 97.4795
R16103 dvss.n4377 dvss.t2257 97.4077
R16104 dvss.n6968 dvss.t1070 97.0786
R16105 dvss.n6784 dvss.t905 97.0786
R16106 dvss.n5984 dvss.t1366 97.0786
R16107 dvss.n6014 dvss.t1557 97.0786
R16108 dvss.n5890 dvss.t480 97.0786
R16109 dvss.n5801 dvss.t2157 97.0786
R16110 dvss.n2112 dvss.t605 97.0786
R16111 dvss.n1995 dvss.t271 97.0786
R16112 dvss.n1657 dvss.t115 97.0786
R16113 dvss.n3136 dvss.n3126 95.7988
R16114 dvss.t1009 dvss.t2149 92.7208
R16115 dvss dvss.t718 92.7208
R16116 dvss.t1239 dvss.t2186 92.7208
R16117 dvss.t1435 dvss.t2211 92.7208
R16118 dvss.t2015 dvss.t193 92.7208
R16119 dvss dvss.t211 92.7208
R16120 dvss.n6279 dvss.t1479 92.7071
R16121 dvss.n6209 dvss.t1382 92.7071
R16122 dvss.n3130 dvss.n3129 90.0716
R16123 dvss.n6881 dvss.n6880 90.0716
R16124 dvss.n141 dvss.n140 90.0716
R16125 dvss.n553 dvss.n552 90.0716
R16126 dvss.n6140 dvss.n6139 90.0716
R16127 dvss.n960 dvss.n959 90.0716
R16128 dvss.n907 dvss.n906 90.0716
R16129 dvss.n2037 dvss.n2036 90.0716
R16130 dvss.n1895 dvss.n1894 90.0716
R16131 dvss.n1780 dvss.n1779 90.0716
R16132 dvss.n1611 dvss.n1610 90.0716
R16133 dvss.n6376 dvss.n6375 90.0716
R16134 dvss.n6325 dvss.n6324 90.0716
R16135 dvss.n6259 dvss.n6258 90.0716
R16136 dvss.n5556 dvss.n5555 90.0716
R16137 dvss.n5502 dvss.n5501 90.0716
R16138 dvss.n5252 dvss.n5251 90.0716
R16139 dvss.n5213 dvss.n5212 90.0716
R16140 dvss.n5174 dvss.n5173 90.0716
R16141 dvss.n5135 dvss.n5134 90.0716
R16142 dvss.n5115 dvss.n5114 90.0716
R16143 dvss.t1068 dvss.n6948 89.9376
R16144 dvss.n225 dvss.t911 89.9376
R16145 dvss.n688 dvss.t1561 89.9376
R16146 dvss.t1372 dvss.n6207 89.9376
R16147 dvss.n1121 dvss.t488 89.9376
R16148 dvss.n1033 dvss.t2165 89.9376
R16149 dvss.t609 dvss.n2104 89.9376
R16150 dvss.n1469 dvss.t273 89.9376
R16151 dvss.n1538 dvss.t105 89.9376
R16152 dvss.n1681 dvss.t130 87.9472
R16153 dvss.t1623 dvss.n4798 86.2322
R16154 dvss.n4798 dvss.t1671 86.2322
R16155 dvss.n6315 dvss.n121 85.5759
R16156 dvss.n6240 dvss.n6239 85.5759
R16157 dvss.n3004 dvss.n3003 84.6851
R16158 dvss.t1012 dvss.t1770 84.2917
R16159 dvss.t158 dvss.t1470 84.2917
R16160 dvss.t120 dvss.t2101 84.2917
R16161 dvss dvss.t1550 84.2917
R16162 dvss.t1505 dvss.t1850 84.2917
R16163 dvss.t1907 dvss.t1048 84.2917
R16164 dvss.n427 dvss.t651 84.171
R16165 dvss.n3308 dvss.t1464 84.0341
R16166 dvss.n4549 dvss.t2118 83.899
R16167 dvss.n4556 dvss.t853 83.899
R16168 dvss.n4541 dvss.t849 83.8933
R16169 dvss.n2301 dvss.t1639 83.4205
R16170 dvss.n4843 dvss.t1606 83.4205
R16171 dvss.n4830 dvss.t1666 83.4205
R16172 dvss.n2315 dvss.t1654 83.4205
R16173 dvss.n2309 dvss.t1681 83.4205
R16174 dvss.n2303 dvss.t1600 83.1135
R16175 dvss.n6437 dvss.n11 83.0194
R16176 dvss.n6861 dvss.n66 83.0194
R16177 dvss.n6715 dvss.n6714 83.0194
R16178 dvss.n609 dvss.n507 83.0194
R16179 dvss.n6120 dvss.n790 83.0194
R16180 dvss.n1054 dvss.n849 83.0194
R16181 dvss.n5731 dvss.n5730 83.0194
R16182 dvss.n2017 dvss.n1440 83.0194
R16183 dvss.n1873 dvss.n1506 83.0194
R16184 dvss.n3346 dvss.n3345 81.965
R16185 dvss.n4072 dvss.n4056 81.965
R16186 dvss.t1105 dvss.n6817 81.3362
R16187 dvss.n103 dvss.t1412 81.3362
R16188 dvss.n5929 dvss.t2205 81.3362
R16189 dvss.n6002 dvss.t1001 81.3362
R16190 dvss.n832 dvss.t671 81.3362
R16191 dvss.t1117 dvss.n868 81.3362
R16192 dvss.t1492 dvss.n2005 81.3362
R16193 dvss.t1313 dvss.n1639 81.3362
R16194 dvss.t265 dvss.n1631 81.3362
R16195 dvss.n7022 dvss.n7021 79.7974
R16196 dvss.n6310 dvss.t1473 78.4446
R16197 dvss.n6238 dvss.t1380 78.4446
R16198 dvss.n3003 dvss.t646 77.0434
R16199 dvss.n3279 dvss.n3274 76.7239
R16200 dvss.n3281 dvss.n3279 76.7239
R16201 dvss.n6940 dvss.n34 76.7239
R16202 dvss.n6485 dvss.n34 76.7239
R16203 dvss.n169 dvss.n74 76.7239
R16204 dvss.n6867 dvss.n74 76.7239
R16205 dvss.n709 dvss.n588 76.7239
R16206 dvss.n709 dvss.n708 76.7239
R16207 dvss.n6199 dvss.n758 76.7239
R16208 dvss.n758 dvss.n757 76.7239
R16209 dvss.n5643 dvss.n798 76.7239
R16210 dvss.n6126 dvss.n798 76.7239
R16211 dvss.n5681 dvss.n942 76.7239
R16212 dvss.n5681 dvss.n5680 76.7239
R16213 dvss.n2096 dvss.n1408 76.7239
R16214 dvss.n1408 dvss.n1407 76.7239
R16215 dvss.n1943 dvss.n1448 76.7239
R16216 dvss.n2023 dvss.n1448 76.7239
R16217 dvss.n1863 dvss.n1513 76.7239
R16218 dvss.n1864 dvss.n1863 76.7239
R16219 dvss.n6421 dvss.n6414 76.7239
R16220 dvss.n6423 dvss.n6421 76.7239
R16221 dvss.n6562 dvss.n6558 76.7239
R16222 dvss.n6558 dvss.n6557 76.7239
R16223 dvss.n6300 dvss.n482 76.7239
R16224 dvss.n6301 dvss.n6300 76.7239
R16225 dvss.n6230 dvss.n511 76.7239
R16226 dvss.n6233 dvss.n6230 76.7239
R16227 dvss.n5535 dvss.n5529 76.7239
R16228 dvss.n5537 dvss.n5535 76.7239
R16229 dvss.n5278 dvss.n5273 76.7239
R16230 dvss.n5280 dvss.n5278 76.7239
R16231 dvss.n5239 dvss.n5234 76.7239
R16232 dvss.n5241 dvss.n5239 76.7239
R16233 dvss.n5200 dvss.n5195 76.7239
R16234 dvss.n5202 dvss.n5200 76.7239
R16235 dvss.n5161 dvss.n5156 76.7239
R16236 dvss.n5163 dvss.n5161 76.7239
R16237 dvss.n4856 dvss.t1665 76.357
R16238 dvss.n1153 dvss.t1605 76.357
R16239 dvss.n6480 dvss.t1060 76.1011
R16240 dvss.n6862 dvss.t901 76.1011
R16241 dvss.t1553 dvss.n122 76.1011
R16242 dvss.n651 dvss.t1370 76.1011
R16243 dvss.n6121 dvss.t490 76.1011
R16244 dvss.n1051 dvss.t2161 76.1011
R16245 dvss.t611 dvss.n888 76.1011
R16246 dvss.n2018 dvss.t275 76.1011
R16247 dvss.t111 dvss.n1851 76.1011
R16248 dvss.t1103 dvss.n6806 76.0887
R16249 dvss.t1414 dvss.n6754 76.0887
R16250 dvss.t2203 dvss.n5930 76.0887
R16251 dvss.t1005 dvss.n6003 76.0887
R16252 dvss.t663 dvss.n5860 76.0887
R16253 dvss.n5769 dvss.t1113 76.0887
R16254 dvss.t1490 dvss.n2006 76.0887
R16255 dvss.n1638 dvss.t1311 76.0887
R16256 dvss.t263 dvss.n1632 76.0887
R16257 dvss.t688 dvss.t2065 75.8626
R16258 dvss.t1215 dvss.t921 75.8626
R16259 dvss.n6567 dvss.t1521 74.7229
R16260 dvss.n6526 dvss.t1082 74.7229
R16261 dvss.n2994 dvss.t644 74.2862
R16262 dvss.n7044 dvss.n7043 73.1255
R16263 dvss.n7043 dvss.n7042 73.1255
R16264 dvss.n7020 dvss.n7001 73.1255
R16265 dvss.n7021 dvss.n7020 73.1255
R16266 dvss.n3215 dvss 73.0358
R16267 dvss.n3230 dvss 73.0358
R16268 dvss.n6920 dvss 73.0358
R16269 dvss.n6936 dvss 73.0358
R16270 dvss dvss.n6692 73.0358
R16271 dvss.n6682 dvss 73.0358
R16272 dvss dvss.n736 73.0358
R16273 dvss.n726 dvss 73.0358
R16274 dvss.n6179 dvss 73.0358
R16275 dvss.n6195 dvss 73.0358
R16276 dvss.n1087 dvss 73.0358
R16277 dvss.n1098 dvss 73.0358
R16278 dvss dvss.n5708 73.0358
R16279 dvss.n5698 dvss 73.0358
R16280 dvss.n2076 dvss 73.0358
R16281 dvss.n2092 dvss 73.0358
R16282 dvss dvss.n1478 73.0358
R16283 dvss dvss.n1923 73.0358
R16284 dvss dvss.n1544 73.0358
R16285 dvss dvss.n1808 73.0358
R16286 dvss.n6803 dvss 73.0358
R16287 dvss.n6825 dvss 73.0358
R16288 dvss.n6748 dvss 73.0358
R16289 dvss.n6763 dvss 73.0358
R16290 dvss.n5961 dvss 73.0358
R16291 dvss.n6034 dvss 73.0358
R16292 dvss.n5914 dvss 73.0358
R16293 dvss.n6084 dvss 73.0358
R16294 dvss.n5854 dvss 73.0358
R16295 dvss.n5869 dvss 73.0358
R16296 dvss dvss.n865 73.0358
R16297 dvss dvss.n5778 73.0358
R16298 dvss.n1331 dvss 73.0358
R16299 dvss.n2128 dvss 73.0358
R16300 dvss.n1300 dvss 73.0358
R16301 dvss.n2183 dvss 73.0358
R16302 dvss.n1269 dvss 73.0358
R16303 dvss.n2233 dvss 73.0358
R16304 dvss.n2567 dvss.t441 72.8576
R16305 dvss.n2936 dvss.t435 72.8576
R16306 dvss.n2926 dvss.t425 72.8576
R16307 dvss.n2848 dvss.t439 72.8576
R16308 dvss.n2682 dvss.t716 72.8576
R16309 dvss.n2700 dvss.t945 72.8576
R16310 dvss.n3735 dvss.t960 72.8576
R16311 dvss.n3736 dvss.t407 72.8576
R16312 dvss.n3650 dvss.t431 72.8576
R16313 dvss.n3841 dvss.t437 72.8576
R16314 dvss.n3851 dvss.t419 72.8576
R16315 dvss.n3944 dvss.t1423 72.8576
R16316 dvss.n3952 dvss.t411 72.8576
R16317 dvss.n3560 dvss.t176 72.8576
R16318 dvss.n2370 dvss.t953 72.8576
R16319 dvss.n2400 dvss.t949 72.8576
R16320 dvss.n4036 dvss.t957 72.8576
R16321 dvss.n4139 dvss.t965 72.8576
R16322 dvss.n4200 dvss.t423 72.8576
R16323 dvss.n4208 dvss.t1427 72.8576
R16324 dvss.t2025 dvss.t1177 70.8111
R16325 dvss.t1177 dvss.t1057 70.8111
R16326 dvss.t1057 dvss.t632 70.8111
R16327 dvss.t632 dvss.t2207 70.8111
R16328 dvss.t1443 dvss.t2062 70.8111
R16329 dvss.t2026 dvss.t895 70.8111
R16330 dvss.t1178 dvss.t2026 70.8111
R16331 dvss.n2425 dvss.t1569 70.0005
R16332 dvss.n2931 dvss.t558 70.0005
R16333 dvss.n2922 dvss.t1017 70.0005
R16334 dvss.n2851 dvss.t1268 70.0005
R16335 dvss.n2754 dvss.t832 70.0005
R16336 dvss.n3745 dvss.t286 70.0005
R16337 dvss.n3746 dvss.t1247 70.0005
R16338 dvss.n3778 dvss.t393 70.0005
R16339 dvss.n3833 dvss.t745 70.0005
R16340 dvss.n3856 dvss.t2009 70.0005
R16341 dvss.n3955 dvss.t468 70.0005
R16342 dvss.n3912 dvss.t1238 70.0005
R16343 dvss.n2366 dvss.t310 70.0005
R16344 dvss.n2396 dvss.t542 70.0005
R16345 dvss.n4028 dvss.t1506 70.0005
R16346 dvss.n4099 dvss.t1455 70.0005
R16347 dvss.n4195 dvss.t382 70.0005
R16348 dvss.n4214 dvss.t2003 70.0005
R16349 dvss.n3345 dvss.t843 68.4925
R16350 dvss.n3345 dvss.t554 68.4925
R16351 dvss.n4056 dvss.t2192 68.4925
R16352 dvss.n4056 dvss.t123 68.4925
R16353 dvss.n4039 dvss.t1391 68.1564
R16354 dvss.n2989 dvss.t1985 67.4335
R16355 dvss.t1397 dvss.t1577 67.4335
R16356 dvss.n3338 dvss.t84 67.4335
R16357 dvss.t842 dvss.t1757 67.4335
R16358 dvss.t846 dvss.t1042 67.4335
R16359 dvss.t38 dvss.n3629 67.4335
R16360 dvss dvss.t883 67.4335
R16361 dvss.t2083 dvss.t386 67.4335
R16362 dvss.t2169 dvss.t1281 67.4335
R16363 dvss.n3301 dvss.t1464 67.3778
R16364 dvss.n6999 dvss.n6998 66.9177
R16365 dvss.n7006 dvss.n7005 66.9014
R16366 dvss.n7008 dvss.n7004 66.9014
R16367 dvss.n7010 dvss.n7003 66.9014
R16368 dvss.n422 dvss.n421 66.771
R16369 dvss.n428 dvss.n423 66.771
R16370 dvss.n4846 dvss.n4845 66.7384
R16371 dvss.n4833 dvss.n4832 66.7384
R16372 dvss.n4837 dvss.n4836 66.7384
R16373 dvss.n4841 dvss.n4840 66.7384
R16374 dvss.n2320 dvss.n2313 66.6759
R16375 dvss.n2317 dvss.n2314 66.6759
R16376 dvss.n2311 dvss.n2308 66.6759
R16377 dvss.n7012 dvss.n7011 66.6759
R16378 dvss.n3691 dvss.n3690 66.462
R16379 dvss.n5495 dvss.t517 65.2441
R16380 dvss.n953 dvss.t2193 64.6673
R16381 dvss.n64 dvss.t739 64.6673
R16382 dvss.n663 dvss.t762 64.6673
R16383 dvss.n788 dvss.t1988 64.6673
R16384 dvss.n1008 dvss.t1253 64.6673
R16385 dvss.n1438 dvss.t2034 64.6673
R16386 dvss.n1491 dvss.t2085 64.6673
R16387 dvss.n190 dvss.t2195 64.6673
R16388 dvss.n4114 dvss.n4113 64.6159
R16389 dvss.t1040 dvss.n1557 63.9189
R16390 dvss.n3326 dvss.t2224 63.866
R16391 dvss.n4597 dvss.n4596 63.5738
R16392 dvss.n2325 dvss.n2324 63.2476
R16393 dvss.n6362 dvss.t1513 63.2272
R16394 dvss.n6511 dvss.t1072 63.2272
R16395 dvss.n6982 dvss.n6981 62.9701
R16396 dvss.n6860 dvss.n6859 62.9701
R16397 dvss.n5990 dvss.n5989 62.9701
R16398 dvss.n6718 dvss.n6716 62.9701
R16399 dvss.n6119 dvss.n6118 62.9701
R16400 dvss.n5824 dvss.n5822 62.9701
R16401 dvss.n5732 dvss.n875 62.9701
R16402 dvss.n2016 dvss.n2015 62.9701
R16403 dvss.n1652 dvss.n1651 62.9701
R16404 dvss.n3063 dvss.n3062 62.7697
R16405 dvss.n3055 dvss.n3054 62.7697
R16406 dvss.n3831 dvss.n3830 62.7697
R16407 dvss dvss.n4856 62.3763
R16408 dvss.n2567 dvss.t1442 60.5809
R16409 dvss.n2936 dvss.t942 60.5809
R16410 dvss.n2926 dvss.t749 60.5809
R16411 dvss.n2848 dvss.t1224 60.5809
R16412 dvss.n2700 dvss.t1274 60.5809
R16413 dvss.n3735 dvss.t1084 60.5809
R16414 dvss.n3736 dvss.t918 60.5809
R16415 dvss.n3650 dvss.t1980 60.5809
R16416 dvss.n3841 dvss.t627 60.5809
R16417 dvss.n3851 dvss.t1180 60.5809
R16418 dvss.n3944 dvss.t2210 60.5809
R16419 dvss.n3952 dvss.t1359 60.5809
R16420 dvss.n2370 dvss.t270 60.5809
R16421 dvss.n2400 dvss.t1353 60.5809
R16422 dvss.n4036 dvss.t1264 60.5809
R16423 dvss.n4139 dvss.t1290 60.5809
R16424 dvss.n4200 dvss.t940 60.5809
R16425 dvss.n4208 dvss.t212 60.5809
R16426 dvss.n5511 dvss.n5510 59.6531
R16427 dvss.n5512 dvss.n5511 59.6531
R16428 dvss.n5512 dvss.n1140 59.6531
R16429 dvss.n5521 dvss.n1140 59.6531
R16430 dvss.n5522 dvss.n5521 59.6531
R16431 dvss.n5523 dvss.n5522 59.6531
R16432 dvss.n5609 dvss.n1123 59.6531
R16433 dvss.n5595 dvss.n5542 59.6531
R16434 dvss.n5595 dvss.n5594 59.6531
R16435 dvss.n5594 dvss.n5593 59.6531
R16436 dvss.n5593 dvss.n5543 59.6531
R16437 dvss.n5587 dvss.n5543 59.6531
R16438 dvss.n5586 dvss.n5585 59.6531
R16439 dvss.n5579 dvss.n5563 59.6531
R16440 dvss.n5579 dvss.n5578 59.6531
R16441 dvss.n5578 dvss.n5577 59.6531
R16442 dvss.n5577 dvss.n5564 59.6531
R16443 dvss.n3619 dvss.t863 59.0774
R16444 dvss.t1219 dvss.t773 59.0043
R16445 dvss dvss.t579 59.0043
R16446 dvss.t2132 dvss.t768 59.0043
R16447 dvss.t2179 dvss.t1398 59.0043
R16448 dvss.t735 dvss.t1500 59.0043
R16449 dvss.t2123 dvss.t732 59.0043
R16450 dvss.n2817 dvss.t101 58.5719
R16451 dvss.n4332 dvss.t178 58.5719
R16452 dvss.n4566 dvss.t855 57.875
R16453 dvss.n4605 dvss.t791 57.875
R16454 dvss.n5006 dvss.t2122 57.875
R16455 dvss.t291 dvss.n7019 57.4543
R16456 dvss.n3274 dvss.n3272 57.0829
R16457 dvss.n3278 dvss.n3276 57.0829
R16458 dvss.n6940 dvss.n35 57.0829
R16459 dvss.n6451 dvss.n6450 57.0829
R16460 dvss.n169 dvss.n168 57.0829
R16461 dvss.n6668 dvss.n6666 57.0829
R16462 dvss.n588 dvss.n587 57.0829
R16463 dvss.n712 dvss.n710 57.0829
R16464 dvss.n6199 dvss.n759 57.0829
R16465 dvss.n537 dvss.n536 57.0829
R16466 dvss.n5643 dvss.n5642 57.0829
R16467 dvss.n5631 dvss.n5629 57.0829
R16468 dvss.n942 dvss.n941 57.0829
R16469 dvss.n5684 dvss.n5682 57.0829
R16470 dvss.n2096 dvss.n1409 57.0829
R16471 dvss.n1360 dvss.n1359 57.0829
R16472 dvss.n1943 dvss.n1465 57.0829
R16473 dvss.n1971 dvss.n1969 57.0829
R16474 dvss.n1513 dvss.n1512 57.0829
R16475 dvss.n1862 dvss.n1515 57.0829
R16476 dvss.n6414 dvss.n6412 57.0829
R16477 dvss.n6420 dvss.n6416 57.0829
R16478 dvss.n6562 dvss.n6561 57.0829
R16479 dvss.n6348 dvss.n6346 57.0829
R16480 dvss.n482 dvss.n481 57.0829
R16481 dvss.n6299 dvss.n484 57.0829
R16482 dvss.n511 dvss.n510 57.0829
R16483 dvss.n6229 dvss.n513 57.0829
R16484 dvss.n5529 dvss.n1137 57.0829
R16485 dvss.n5534 dvss.n5532 57.0829
R16486 dvss.n5273 dvss.n5271 57.0829
R16487 dvss.n5277 dvss.n5275 57.0829
R16488 dvss.n5234 dvss.n5232 57.0829
R16489 dvss.n5238 dvss.n5236 57.0829
R16490 dvss.n5195 dvss.n5193 57.0829
R16491 dvss.n5199 dvss.n5197 57.0829
R16492 dvss.n5156 dvss.n5154 57.0829
R16493 dvss.n5160 dvss.n5158 57.0829
R16494 dvss.n6335 dvss.t1085 57.076
R16495 dvss.n6253 dvss.t1319 57.076
R16496 dvss.t1647 dvss.t1665 56.6405
R16497 dvss.t1635 dvss.t1647 56.6405
R16498 dvss.t1668 dvss.t1635 56.6405
R16499 dvss.t1620 dvss.t1668 56.6405
R16500 dvss.t1641 dvss.t1626 56.6405
R16501 dvss.t1644 dvss.t1659 56.6405
R16502 dvss.t1605 dvss.t1644 56.6405
R16503 dvss.n5603 dvss.n5602 56.5704
R16504 dvss.n3619 dvss.t314 56.3082
R16505 dvss.n3664 dvss.t600 55.7148
R16506 dvss.n3473 dvss.t1242 55.7148
R16507 dvss.n4057 dvss.t933 55.7148
R16508 dvss.t1537 dvss.n1122 53.4393
R16509 dvss.n2688 dvss.t1019 52.8576
R16510 dvss.n3508 dvss.t689 52.8576
R16511 dvss.n2385 dvss.t1982 52.8576
R16512 dvss.n5587 dvss.t766 52.8179
R16513 dvss.n4820 dvss.n4819 52.3299
R16514 dvss.n3045 dvss.t455 51.6928
R16515 dvss.t895 dvss.n7022 51.5162
R16516 dvss.n2432 dvss.t2105 51.4291
R16517 dvss.n3923 dvss.t1202 51.4291
R16518 dvss.n3535 dvss.t2045 51.4291
R16519 dvss.n3532 dvss.t847 51.4291
R16520 dvss.n4334 dvss.t623 51.4291
R16521 dvss.n4610 dvss.t474 51.4291
R16522 dvss.n4546 dvss.t725 51.4291
R16523 dvss.n4622 dvss.t2227 51.4291
R16524 dvss.n4895 dvss.t678 51.4291
R16525 dvss.n4900 dvss.t737 51.4291
R16526 dvss.n4905 dvss.t770 51.4291
R16527 dvss.n4910 dvss.t2001 51.4291
R16528 dvss.n1222 dvss.t1022 51.4291
R16529 dvss.n1227 dvss.t2151 51.4291
R16530 dvss.n4216 dvss.t2156 51.4291
R16531 dvss.t1535 dvss.n5601 50.9538
R16532 dvss.t1805 dvss.t448 50.5752
R16533 dvss.t440 dvss 50.5752
R16534 dvss.t619 dvss 50.5752
R16535 dvss.t709 dvss.t844 50.5752
R16536 dvss.t313 dvss.t2080 50.5752
R16537 dvss.t300 dvss.t1915 50.5752
R16538 dvss.t1351 dvss.t369 50.5752
R16539 dvss.t1475 dvss.n6308 49.9195
R16540 dvss.n6223 dvss.t1374 49.9195
R16541 dvss.n4822 dvss.n1238 49.781
R16542 dvss.n7023 dvss.t1178 49.3028
R16543 dvss.n6472 dvss.t1062 48.4282
R16544 dvss.t903 dvss.n6658 48.4282
R16545 dvss.n699 dvss.t1555 48.4282
R16546 dvss.t1362 dvss.n647 48.4282
R16547 dvss.t482 dvss.n5621 48.4282
R16548 dvss.t2167 dvss.n1047 48.4282
R16549 dvss.n1393 dvss.t615 48.4282
R16550 dvss.t279 dvss.n1961 48.4282
R16551 dvss.n1853 dvss.t107 48.4282
R16552 dvss.t1626 dvss.n1145 47.32
R16553 dvss.n3620 dvss.n3619 46.2505
R16554 dvss.n3190 dvss.n3189 46.2505
R16555 dvss.n3181 dvss.n3180 46.2505
R16556 dvss.n54 dvss.n53 46.2505
R16557 dvss.n37 dvss.n36 46.2505
R16558 dvss.n151 dvss.n150 46.2505
R16559 dvss.n153 dvss.n152 46.2505
R16560 dvss.n563 dvss.n562 46.2505
R16561 dvss.n565 dvss.n564 46.2505
R16562 dvss.n778 dvss.n777 46.2505
R16563 dvss.n761 dvss.n760 46.2505
R16564 dvss.n1084 dvss.n1083 46.2505
R16565 dvss.n1095 dvss.n1094 46.2505
R16566 dvss.n917 dvss.n916 46.2505
R16567 dvss.n919 dvss.n918 46.2505
R16568 dvss.n1428 dvss.n1427 46.2505
R16569 dvss.n1411 dvss.n1410 46.2505
R16570 dvss.n1908 dvss.n1907 46.2505
R16571 dvss.n1922 dvss.n1921 46.2505
R16572 dvss.n1787 dvss.n1783 46.2505
R16573 dvss.n1807 dvss.n1806 46.2505
R16574 dvss.n6843 dvss.n6797 46.2505
R16575 dvss.n6834 dvss.n6804 46.2505
R16576 dvss.n108 dvss.n107 46.2505
R16577 dvss.n99 dvss.n98 46.2505
R16578 dvss.n6052 dvss.n5956 46.2505
R16579 dvss.n6043 dvss.n5962 46.2505
R16580 dvss.n6102 dvss.n5908 46.2505
R16581 dvss.n6093 dvss.n5915 46.2505
R16582 dvss.n837 dvss.n836 46.2505
R16583 dvss.n828 dvss.n827 46.2505
R16584 dvss.n5761 dvss.n5760 46.2505
R16585 dvss.n5777 dvss.n5776 46.2505
R16586 dvss.n2146 dvss.n1326 46.2505
R16587 dvss.n2137 dvss.n1332 46.2505
R16588 dvss.n2201 dvss.n1295 46.2505
R16589 dvss.n2192 dvss.n1301 46.2505
R16590 dvss.n2251 dvss.n1263 46.2505
R16591 dvss.n2242 dvss.n1270 46.2505
R16592 dvss.n2707 dvss.t1108 45.7148
R16593 dvss.n3661 dvss.t323 45.7148
R16594 dvss.n3853 dvss.t1432 45.7148
R16595 dvss.n3459 dvss.t1092 45.7148
R16596 dvss.n2388 dvss.t2041 45.7148
R16597 dvss.n2399 dvss.t391 45.7148
R16598 dvss.n4587 dvss.t2095 45.7148
R16599 dvss.n4578 dvss.t899 45.7148
R16600 dvss.n4585 dvss.t800 45.7148
R16601 dvss.n5017 dvss.t1325 45.7148
R16602 dvss.n5047 dvss.t2114 45.7148
R16603 dvss.n5054 dvss.t2213 45.7148
R16604 dvss.n1219 dvss.t1303 45.7148
R16605 dvss.n4922 dvss.t856 45.7148
R16606 dvss.n4920 dvss.t1033 45.7148
R16607 dvss.n4043 dvss.t1318 45.7148
R16608 dvss.n4158 dvss.t169 45.7148
R16609 dvss.n437 dvss.n436 45.0005
R16610 dvss.n430 dvss.n417 45.0005
R16611 dvss.n417 dvss.t819 45.0005
R16612 dvss.n418 dvss.n416 45.0005
R16613 dvss.t819 dvss.n416 45.0005
R16614 dvss.n334 dvss.n333 45.0005
R16615 dvss.n6612 dvss.n6611 45.0005
R16616 dvss.n7041 dvss.t2025 44.9596
R16617 dvss.n3230 dvss 44.424
R16618 dvss.n6936 dvss 44.424
R16619 dvss.n6682 dvss 44.424
R16620 dvss.n726 dvss 44.424
R16621 dvss.n6195 dvss 44.424
R16622 dvss.n1098 dvss 44.424
R16623 dvss.n5698 dvss 44.424
R16624 dvss.n2092 dvss 44.424
R16625 dvss.n1923 dvss 44.424
R16626 dvss.n1808 dvss 44.424
R16627 dvss.n6825 dvss 44.424
R16628 dvss.n6763 dvss 44.424
R16629 dvss.n6034 dvss 44.424
R16630 dvss.n6084 dvss 44.424
R16631 dvss.n5869 dvss 44.424
R16632 dvss.n5778 dvss 44.424
R16633 dvss.n2128 dvss 44.424
R16634 dvss.n2183 dvss 44.424
R16635 dvss.n2233 dvss 44.424
R16636 dvss.t1458 dvss.n3145 43.698
R16637 dvss.n1122 dvss.t1543 43.4972
R16638 dvss.t397 dvss.n1761 43.2419
R16639 dvss.t755 dvss.n5124 43.2419
R16640 dvss.t414 dvss.t996 42.1461
R16641 dvss dvss.t434 42.1461
R16642 dvss.t643 dvss.t525 42.1461
R16643 dvss.t1471 dvss 42.1461
R16644 dvss.t1332 dvss.t2044 42.1461
R16645 dvss.t601 dvss.t545 42.1461
R16646 dvss.t91 dvss.t1565 42.1461
R16647 dvss dvss.t952 42.1461
R16648 dvss.n4039 dvss.t1250 41.6479
R16649 dvss.n3062 dvss.t845 41.539
R16650 dvss.n3063 dvss.t321 41.539
R16651 dvss.n3054 dvss.t841 41.539
R16652 dvss.n3055 dvss.t604 41.539
R16653 dvss.n3830 dvss.t839 41.539
R16654 dvss.n3831 dvss.t1997 41.539
R16655 dvss.n4114 dvss.t1252 41.539
R16656 dvss.n3690 dvss.t1194 40.6159
R16657 dvss.n3691 dvss.t2061 40.6159
R16658 dvss.n4113 dvss.t306 40.6159
R16659 dvss.n5601 dvss.n1132 40.3903
R16660 dvss.n2692 dvss.t586 40.0005
R16661 dvss.n2692 dvss.t572 40.0005
R16662 dvss.n2811 dvss.t2133 40.0005
R16663 dvss.n2811 dvss.t2129 40.0005
R16664 dvss.n2810 dvss.t594 40.0005
R16665 dvss.n2810 dvss.t2139 40.0005
R16666 dvss.n2808 dvss.t566 40.0005
R16667 dvss.n2808 dvss.t582 40.0005
R16668 dvss.n2693 dvss.t596 40.0005
R16669 dvss.n2693 dvss.t576 40.0005
R16670 dvss.n2787 dvss.t584 40.0005
R16671 dvss.n2787 dvss.t570 40.0005
R16672 dvss.n2689 dvss.t568 40.0005
R16673 dvss.n2688 dvss.t878 40.0005
R16674 dvss.n2798 dvss.t578 40.0005
R16675 dvss.n2798 dvss.t592 40.0005
R16676 dvss.n2805 dvss.t574 40.0005
R16677 dvss.n2805 dvss.t588 40.0005
R16678 dvss.n3768 dvss.t149 40.0005
R16679 dvss.n3768 dvss.t161 40.0005
R16680 dvss.n3774 dvss.t145 40.0005
R16681 dvss.n3774 dvss.t159 40.0005
R16682 dvss.n3647 dvss.t141 40.0005
R16683 dvss.n3647 dvss.t155 40.0005
R16684 dvss.n3784 dvss.t153 40.0005
R16685 dvss.n3644 dvss.t165 40.0005
R16686 dvss.n3644 dvss.t151 40.0005
R16687 dvss.n3797 dvss.t163 40.0005
R16688 dvss.n3797 dvss.t139 40.0005
R16689 dvss.n3799 dvss.t157 40.0005
R16690 dvss.n3799 dvss.t137 40.0005
R16691 dvss.n3814 dvss.t143 40.0005
R16692 dvss.n3814 dvss.t889 40.0005
R16693 dvss.n3817 dvss.t893 40.0005
R16694 dvss.n3817 dvss.t891 40.0005
R16695 dvss.n3486 dvss.t1246 40.0005
R16696 dvss.n3486 dvss.t1240 40.0005
R16697 dvss.n3473 dvss.t2073 40.0005
R16698 dvss.n3508 dvss.t2102 40.0005
R16699 dvss.n2385 dvss.t2075 40.0005
R16700 dvss.n4144 dvss.t2141 40.0005
R16701 dvss.n4144 dvss.t2137 40.0005
R16702 dvss.n4147 dvss.t2127 40.0005
R16703 dvss.n4147 dvss.t190 40.0005
R16704 dvss.n4150 dvss.t196 40.0005
R16705 dvss.n4150 dvss.t208 40.0005
R16706 dvss.n4156 dvss.t188 40.0005
R16707 dvss.n4156 dvss.t204 40.0005
R16708 dvss.n4160 dvss.t182 40.0005
R16709 dvss.n4160 dvss.t200 40.0005
R16710 dvss.n4014 dvss.t180 40.0005
R16711 dvss.n4016 dvss.t210 40.0005
R16712 dvss.n4016 dvss.t192 40.0005
R16713 dvss.n4019 dvss.t206 40.0005
R16714 dvss.n4019 dvss.t186 40.0005
R16715 dvss.n4020 dvss.t202 40.0005
R16716 dvss.n4020 dvss.t184 40.0005
R16717 dvss.n3045 dvss.t1991 39.6928
R16718 dvss.t1479 dvss.n487 39.2225
R16719 dvss.t1382 dvss.n6208 39.2225
R16720 dvss.n2418 dvss.t926 38.7697
R16721 dvss.n3011 dvss.t1214 38.7697
R16722 dvss.n3633 dvss.t2084 38.7697
R16723 dvss.n3979 dvss.t1047 38.7697
R16724 dvss.n3510 dvss.t121 38.7697
R16725 dvss.n3510 dvss.t2066 38.7697
R16726 dvss.n3528 dvss.t1256 38.7697
R16727 dvss.n2574 dvss.t446 38.5719
R16728 dvss.n2574 dvss.t708 38.5719
R16729 dvss.n2935 dvss.t994 38.5719
R16730 dvss.n2935 dvss.t714 38.5719
R16731 dvss.n3002 dvss.t528 38.5719
R16732 dvss.n3002 dvss.t712 38.5719
R16733 dvss.n3059 dvss.t1220 38.5719
R16734 dvss.n3059 dvss.t710 38.5719
R16735 dvss.n2710 dvss.t1337 38.5719
R16736 dvss.n2710 dvss.t719 38.5719
R16737 dvss.n2779 dvss.t1270 38.5719
R16738 dvss.n2779 dvss.t705 38.5719
R16739 dvss.n2689 dvss.t580 38.5719
R16740 dvss.n3708 dvss.t699 38.5719
R16741 dvss.n3708 dvss.t1469 38.5719
R16742 dvss.n3706 dvss.t751 38.5719
R16743 dvss.n3706 dvss.t706 38.5719
R16744 dvss.n3721 dvss.t521 38.5719
R16745 dvss.n3721 dvss.t703 38.5719
R16746 dvss.n3656 dvss.t729 38.5719
R16747 dvss.n3656 dvss.t2029 38.5719
R16748 dvss.n3784 dvss.t135 38.5719
R16749 dvss.n3843 dvss.t701 38.5719
R16750 dvss.n3843 dvss.t2092 38.5719
R16751 dvss.n3848 dvss.t471 38.5719
R16752 dvss.n3848 dvss.t495 38.5719
R16753 dvss.n3858 dvss.t1451 38.5719
R16754 dvss.n3858 dvss.t2007 38.5719
R16755 dvss.n3921 dvss.t33 38.5719
R16756 dvss.n3921 dvss.t497 38.5719
R16757 dvss.n3920 dvss.t694 38.5719
R16758 dvss.n3920 dvss.t493 38.5719
R16759 dvss.n3980 dvss.t1090 38.5719
R16760 dvss.n3980 dvss.t318 38.5719
R16761 dvss.n2376 dvss.t28 38.5719
R16762 dvss.n2376 dvss.t501 38.5719
R16763 dvss.n2383 dvss.t1510 38.5719
R16764 dvss.n2383 dvss.t2039 38.5719
R16765 dvss.n2393 dvss.t2185 38.5719
R16766 dvss.n2393 dvss.t1059 38.5719
R16767 dvss.n4304 dvss.t1282 38.5719
R16768 dvss.n4304 dvss.t499 38.5719
R16769 dvss.n4031 dvss.t1260 38.5719
R16770 dvss.n4031 dvss.t509 38.5719
R16771 dvss.n4046 dvss.t1529 38.5719
R16772 dvss.n4046 dvss.t916 38.5719
R16773 dvss.n4148 dvss.t1287 38.5719
R16774 dvss.n4148 dvss.t503 38.5719
R16775 dvss.n4014 dvss.t198 38.5719
R16776 dvss.n4015 dvss.t464 38.5719
R16777 dvss.n4015 dvss.t1 38.5719
R16778 dvss.n4201 dvss.t505 38.5719
R16779 dvss.n4201 dvss.t23 38.5719
R16780 dvss.n4206 dvss.t937 38.5719
R16781 dvss.n4206 dvss.t507 38.5719
R16782 dvss.n4213 dvss.t1198 38.5719
R16783 dvss.n4213 dvss.t1200 38.5719
R16784 dvss.n6949 dvss.t1068 38.0508
R16785 dvss.n6647 dvss.t911 38.0508
R16786 dvss.t1561 dvss.n487 38.0508
R16787 dvss.n6208 dvss.t1372 38.0508
R16788 dvss.n5610 dvss.t488 38.0508
R16789 dvss.t2165 dvss.n862 38.0508
R16790 dvss.n2105 dvss.t609 38.0508
R16791 dvss.n1985 dvss.t273 38.0508
R16792 dvss.t105 dvss.n1530 38.0508
R16793 dvss.n4816 dvss.n1234 37.9094
R16794 dvss.n4828 dvss.n1234 37.9005
R16795 dvss.n1565 dvss.t758 37.7206
R16796 dvss.n1255 dvss.t403 37.7206
R16797 dvss.t1456 dvss.n3299 36.9753
R16798 dvss.n6605 dvss.n6604 36.563
R16799 dvss.t1029 dvss.t1257 36.1649
R16800 dvss.n3334 dvss.n3128 36.1417
R16801 dvss.n3132 dvss.n3128 36.1417
R16802 dvss.n3328 dvss.n3132 36.1417
R16803 dvss.n3328 dvss.n3133 36.1417
R16804 dvss.n3322 dvss.n3133 36.1417
R16805 dvss.n3322 dvss.n3321 36.1417
R16806 dvss.n3321 dvss.n3320 36.1417
R16807 dvss.n3320 dvss.n3143 36.1417
R16808 dvss.n3314 dvss.n3143 36.1417
R16809 dvss.n3314 dvss.n3313 36.1417
R16810 dvss.n3313 dvss.n3312 36.1417
R16811 dvss.n3312 dvss.n3151 36.1417
R16812 dvss.n3306 dvss.n3151 36.1417
R16813 dvss.n3306 dvss.n3305 36.1417
R16814 dvss.n3305 dvss.n3304 36.1417
R16815 dvss.n3304 dvss.n3158 36.1417
R16816 dvss.n3297 dvss.n3158 36.1417
R16817 dvss.n3297 dvss.n3296 36.1417
R16818 dvss.n3296 dvss.n3295 36.1417
R16819 dvss.n3295 dvss.n3285 36.1417
R16820 dvss.n3289 dvss.n3285 36.1417
R16821 dvss.n5493 dvss.n5492 36.1417
R16822 dvss.n5492 dvss.n5491 36.1417
R16823 dvss.n5491 dvss.n5490 36.1417
R16824 dvss.n5490 dvss.n5488 36.1417
R16825 dvss.n5488 dvss.n5485 36.1417
R16826 dvss.n5485 dvss.n5484 36.1417
R16827 dvss.n5484 dvss.n5481 36.1417
R16828 dvss.n5481 dvss.n5480 36.1417
R16829 dvss.n5480 dvss.n5477 36.1417
R16830 dvss.n5477 dvss.n5476 36.1417
R16831 dvss.n5476 dvss.n5473 36.1417
R16832 dvss.n5473 dvss.n5472 36.1417
R16833 dvss.n5472 dvss.n5469 36.1417
R16834 dvss.n5469 dvss.n5468 36.1417
R16835 dvss.n5468 dvss.n5465 36.1417
R16836 dvss.n5465 dvss.n5464 36.1417
R16837 dvss.n5461 dvss.n5460 36.1417
R16838 dvss.n5460 dvss.n5457 36.1417
R16839 dvss.n5457 dvss.n5456 36.1417
R16840 dvss.n5456 dvss.n5453 36.1417
R16841 dvss.n5453 dvss.n5452 36.1417
R16842 dvss.n5452 dvss.n5449 36.1417
R16843 dvss.n5449 dvss.n5448 36.1417
R16844 dvss.n5448 dvss.n5445 36.1417
R16845 dvss.n5445 dvss.n5444 36.1417
R16846 dvss.n5444 dvss.n5441 36.1417
R16847 dvss.n5441 dvss.n5440 36.1417
R16848 dvss.n5440 dvss.n5437 36.1417
R16849 dvss.n5437 dvss.n5436 36.1417
R16850 dvss.n5436 dvss.n5433 36.1417
R16851 dvss.n5433 dvss.n5432 36.1417
R16852 dvss.n5432 dvss.n5429 36.1417
R16853 dvss.n5429 dvss.n5428 36.1417
R16854 dvss.n5428 dvss.n5425 36.1417
R16855 dvss.n5425 dvss.n5424 36.1417
R16856 dvss.n5424 dvss.n5421 36.1417
R16857 dvss.n5421 dvss.n5420 36.1417
R16858 dvss.n5417 dvss.n5416 36.1417
R16859 dvss.n5416 dvss.n5413 36.1417
R16860 dvss.n5413 dvss.n5412 36.1417
R16861 dvss.n5412 dvss.n5409 36.1417
R16862 dvss.n5409 dvss.n5408 36.1417
R16863 dvss.n5408 dvss.n5405 36.1417
R16864 dvss.n5405 dvss.n5404 36.1417
R16865 dvss.n5404 dvss.n5401 36.1417
R16866 dvss.n5401 dvss.n5400 36.1417
R16867 dvss.n5400 dvss.n5397 36.1417
R16868 dvss.n5397 dvss.n5396 36.1417
R16869 dvss.n5396 dvss.n5393 36.1417
R16870 dvss.n5393 dvss.n5392 36.1417
R16871 dvss.n5392 dvss.n5389 36.1417
R16872 dvss.n5389 dvss.n5388 36.1417
R16873 dvss.n5388 dvss.n5385 36.1417
R16874 dvss.n5385 dvss.n5384 36.1417
R16875 dvss.n5384 dvss.n5381 36.1417
R16876 dvss.n5381 dvss.n5380 36.1417
R16877 dvss.n5380 dvss.n5377 36.1417
R16878 dvss.n5377 dvss.n5376 36.1417
R16879 dvss.n5373 dvss.n5372 36.1417
R16880 dvss.n5372 dvss.n5369 36.1417
R16881 dvss.n5369 dvss.n5368 36.1417
R16882 dvss.n5368 dvss.n5365 36.1417
R16883 dvss.n5365 dvss.n5364 36.1417
R16884 dvss.n5364 dvss.n5361 36.1417
R16885 dvss.n5361 dvss.n5360 36.1417
R16886 dvss.n5360 dvss.n5357 36.1417
R16887 dvss.n5357 dvss.n5356 36.1417
R16888 dvss.n5356 dvss.n5353 36.1417
R16889 dvss.n5353 dvss.n5352 36.1417
R16890 dvss.n5352 dvss.n5349 36.1417
R16891 dvss.n5349 dvss.n5348 36.1417
R16892 dvss.n5348 dvss.n5345 36.1417
R16893 dvss.n5345 dvss.n5344 36.1417
R16894 dvss.n5344 dvss.n5341 36.1417
R16895 dvss.n5341 dvss.n5340 36.1417
R16896 dvss.n5340 dvss.n5337 36.1417
R16897 dvss.n5337 dvss.n5336 36.1417
R16898 dvss.n5336 dvss.n5333 36.1417
R16899 dvss.n5333 dvss.n5332 36.1417
R16900 dvss.n5329 dvss.n5328 36.1417
R16901 dvss.n5328 dvss.n5325 36.1417
R16902 dvss.n5325 dvss.n5324 36.1417
R16903 dvss.n5324 dvss.n5321 36.1417
R16904 dvss.n5321 dvss.n5320 36.1417
R16905 dvss.n5320 dvss.n5317 36.1417
R16906 dvss.n5317 dvss.n5316 36.1417
R16907 dvss.n5316 dvss.n5313 36.1417
R16908 dvss.n5313 dvss.n5312 36.1417
R16909 dvss.n5312 dvss.n5309 36.1417
R16910 dvss.n5309 dvss.n5308 36.1417
R16911 dvss.n5308 dvss.n5305 36.1417
R16912 dvss.n5305 dvss.n5304 36.1417
R16913 dvss.n5304 dvss.n5301 36.1417
R16914 dvss.n5301 dvss.n5300 36.1417
R16915 dvss.n5300 dvss.n5297 36.1417
R16916 dvss.n5297 dvss.n5296 36.1417
R16917 dvss.n5296 dvss.n5293 36.1417
R16918 dvss.n5293 dvss.n5292 36.1417
R16919 dvss.n5292 dvss.n5289 36.1417
R16920 dvss.n5289 dvss.n5288 36.1417
R16921 dvss.n5498 dvss.n1149 36.1417
R16922 dvss.n5498 dvss.n1150 36.1417
R16923 dvss.n1150 dvss.n1147 36.1417
R16924 dvss.n5508 dvss.n1147 36.1417
R16925 dvss.n5508 dvss.n1143 36.1417
R16926 dvss.n5514 dvss.n1143 36.1417
R16927 dvss.n5514 dvss.n1142 36.1417
R16928 dvss.n5519 dvss.n1142 36.1417
R16929 dvss.n5519 dvss.n1138 36.1417
R16930 dvss.n5525 dvss.n1138 36.1417
R16931 dvss.n5525 dvss.n1126 36.1417
R16932 dvss.n5607 dvss.n1126 36.1417
R16933 dvss.n5607 dvss.n5606 36.1417
R16934 dvss.n5606 dvss.n5605 36.1417
R16935 dvss.n5605 dvss.n1130 36.1417
R16936 dvss.n5599 dvss.n1130 36.1417
R16937 dvss.n5599 dvss.n5598 36.1417
R16938 dvss.n5598 dvss.n5597 36.1417
R16939 dvss.n5597 dvss.n5540 36.1417
R16940 dvss.n5591 dvss.n5540 36.1417
R16941 dvss.n5591 dvss.n5590 36.1417
R16942 dvss.n5589 dvss.n5549 36.1417
R16943 dvss.n5583 dvss.n5549 36.1417
R16944 dvss.n5583 dvss.n5582 36.1417
R16945 dvss.n5582 dvss.n5581 36.1417
R16946 dvss.n5581 dvss.n5561 36.1417
R16947 dvss.n5575 dvss.n5561 36.1417
R16948 dvss.n5575 dvss.n5574 36.1417
R16949 dvss.n5574 dvss.n5573 36.1417
R16950 dvss.n5573 dvss.n522 36.1417
R16951 dvss.n6211 dvss.n522 36.1417
R16952 dvss.n6211 dvss.n521 36.1417
R16953 dvss.n6218 dvss.n521 36.1417
R16954 dvss.n6218 dvss.n514 36.1417
R16955 dvss.n6226 dvss.n514 36.1417
R16956 dvss.n6226 dvss.n517 36.1417
R16957 dvss.n517 dvss.n509 36.1417
R16958 dvss.n6236 dvss.n509 36.1417
R16959 dvss.n6236 dvss.n505 36.1417
R16960 dvss.n6243 dvss.n505 36.1417
R16961 dvss.n6243 dvss.n504 36.1417
R16962 dvss.n6248 dvss.n504 36.1417
R16963 dvss.n6255 dvss.n500 36.1417
R16964 dvss.n6255 dvss.n498 36.1417
R16965 dvss.n6264 dvss.n498 36.1417
R16966 dvss.n6264 dvss.n495 36.1417
R16967 dvss.n6270 dvss.n495 36.1417
R16968 dvss.n6270 dvss.n494 36.1417
R16969 dvss.n6275 dvss.n494 36.1417
R16970 dvss.n6275 dvss.n490 36.1417
R16971 dvss.n6282 dvss.n490 36.1417
R16972 dvss.n6282 dvss.n489 36.1417
R16973 dvss.n6289 dvss.n489 36.1417
R16974 dvss.n6289 dvss.n485 36.1417
R16975 dvss.n6295 dvss.n485 36.1417
R16976 dvss.n6295 dvss.n479 36.1417
R16977 dvss.n6306 dvss.n479 36.1417
R16978 dvss.n6306 dvss.n480 36.1417
R16979 dvss.n480 dvss.n475 36.1417
R16980 dvss.n6317 dvss.n475 36.1417
R16981 dvss.n6317 dvss.n472 36.1417
R16982 dvss.n6321 dvss.n472 36.1417
R16983 dvss.n6322 dvss.n6321 36.1417
R16984 dvss.n6332 dvss.n471 36.1417
R16985 dvss.n471 dvss.n468 36.1417
R16986 dvss.n468 dvss.n459 36.1417
R16987 dvss.n6577 dvss.n459 36.1417
R16988 dvss.n6577 dvss.n6576 36.1417
R16989 dvss.n6576 dvss.n462 36.1417
R16990 dvss.n6572 dvss.n462 36.1417
R16991 dvss.n6572 dvss.n6571 36.1417
R16992 dvss.n6571 dvss.n465 36.1417
R16993 dvss.n6565 dvss.n465 36.1417
R16994 dvss.n6565 dvss.n230 36.1417
R16995 dvss.n6644 dvss.n230 36.1417
R16996 dvss.n6644 dvss.n6643 36.1417
R16997 dvss.n6643 dvss.n6642 36.1417
R16998 dvss.n6642 dvss.n234 36.1417
R16999 dvss.n6356 dvss.n234 36.1417
R17000 dvss.n6356 dvss.n6350 36.1417
R17001 dvss.n6554 dvss.n6350 36.1417
R17002 dvss.n6554 dvss.n6351 36.1417
R17003 dvss.n6548 dvss.n6351 36.1417
R17004 dvss.n6548 dvss.n6547 36.1417
R17005 dvss.n6546 dvss.n6369 36.1417
R17006 dvss.n6540 dvss.n6369 36.1417
R17007 dvss.n6540 dvss.n6539 36.1417
R17008 dvss.n6539 dvss.n6538 36.1417
R17009 dvss.n6538 dvss.n6381 36.1417
R17010 dvss.n6532 dvss.n6381 36.1417
R17011 dvss.n6532 dvss.n6531 36.1417
R17012 dvss.n6531 dvss.n6530 36.1417
R17013 dvss.n6530 dvss.n6390 36.1417
R17014 dvss.n6524 dvss.n6390 36.1417
R17015 dvss.n6524 dvss.n6523 36.1417
R17016 dvss.n6523 dvss.n6522 36.1417
R17017 dvss.n6522 dvss.n6398 36.1417
R17018 dvss.n6402 dvss.n6398 36.1417
R17019 dvss.n6515 dvss.n6402 36.1417
R17020 dvss.n6515 dvss.n6514 36.1417
R17021 dvss.n6514 dvss.n6513 36.1417
R17022 dvss.n6513 dvss.n6406 36.1417
R17023 dvss.n6507 dvss.n6406 36.1417
R17024 dvss.n6507 dvss.n6506 36.1417
R17025 dvss.n6506 dvss.n6505 36.1417
R17026 dvss.n1698 dvss.n1598 36.1417
R17027 dvss.n1752 dvss.n1598 36.1417
R17028 dvss.n1752 dvss.n1751 36.1417
R17029 dvss.n1751 dvss.n1750 36.1417
R17030 dvss.n1750 dvss.n1749 36.1417
R17031 dvss.n1749 dvss.n1747 36.1417
R17032 dvss.n1747 dvss.n1744 36.1417
R17033 dvss.n1744 dvss.n1743 36.1417
R17034 dvss.n1743 dvss.n1740 36.1417
R17035 dvss.n1740 dvss.n1739 36.1417
R17036 dvss.n1739 dvss.n1736 36.1417
R17037 dvss.n1736 dvss.n1566 36.1417
R17038 dvss.n1757 dvss.n1566 36.1417
R17039 dvss.n1757 dvss.n1567 36.1417
R17040 dvss.n1582 dvss.n1567 36.1417
R17041 dvss.n1582 dvss.n1580 36.1417
R17042 dvss.n1589 dvss.n1580 36.1417
R17043 dvss.n1589 dvss.n1554 36.1417
R17044 dvss.n1554 dvss.n1552 36.1417
R17045 dvss.n1790 dvss.n1552 36.1417
R17046 dvss.n1790 dvss.n1547 36.1417
R17047 dvss.n1799 dvss.n1547 36.1417
R17048 dvss.n1799 dvss.n1542 36.1417
R17049 dvss.n1812 dvss.n1542 36.1417
R17050 dvss.n1812 dvss.n1536 36.1417
R17051 dvss.n1822 dvss.n1536 36.1417
R17052 dvss.n1822 dvss.n1532 36.1417
R17053 dvss.n1832 dvss.n1532 36.1417
R17054 dvss.n1832 dvss.n1527 36.1417
R17055 dvss.n1846 dvss.n1527 36.1417
R17056 dvss.n1846 dvss.n1516 36.1417
R17057 dvss.n1855 dvss.n1516 36.1417
R17058 dvss.n1855 dvss.n1510 36.1417
R17059 dvss.n1867 dvss.n1510 36.1417
R17060 dvss.n1868 dvss.n1867 36.1417
R17061 dvss.n1868 dvss.n1505 36.1417
R17062 dvss.n1505 dvss.n1496 36.1417
R17063 dvss.n1497 dvss.n1496 36.1417
R17064 dvss.n1881 dvss.n1497 36.1417
R17065 dvss.n1881 dvss.n1488 36.1417
R17066 dvss.n1500 dvss.n1488 36.1417
R17067 dvss.n1500 dvss.n1483 36.1417
R17068 dvss.n1904 dvss.n1483 36.1417
R17069 dvss.n1904 dvss.n1479 36.1417
R17070 dvss.n1917 dvss.n1479 36.1417
R17071 dvss.n1917 dvss.n1476 36.1417
R17072 dvss.n1476 dvss.n1473 36.1417
R17073 dvss.n1473 dvss.n1466 36.1417
R17074 dvss.n1466 dvss.n1460 36.1417
R17075 dvss.n1982 dvss.n1460 36.1417
R17076 dvss.n1982 dvss.n1461 36.1417
R17077 dvss.n1945 dvss.n1461 36.1417
R17078 dvss.n1953 dvss.n1945 36.1417
R17079 dvss.n1953 dvss.n1949 36.1417
R17080 dvss.n1949 dvss.n1454 36.1417
R17081 dvss.n2020 dvss.n1454 36.1417
R17082 dvss.n2020 dvss.n1444 36.1417
R17083 dvss.n2053 dvss.n1444 36.1417
R17084 dvss.n2053 dvss.n1445 36.1417
R17085 dvss.n2029 dvss.n1445 36.1417
R17086 dvss.n2035 dvss.n2029 36.1417
R17087 dvss.n2035 dvss.n1433 36.1417
R17088 dvss.n2062 dvss.n1433 36.1417
R17089 dvss.n2063 dvss.n2062 36.1417
R17090 dvss.n2063 dvss.n1429 36.1417
R17091 dvss.n2072 dvss.n1429 36.1417
R17092 dvss.n2072 dvss.n1425 36.1417
R17093 dvss.n1425 dvss.n1421 36.1417
R17094 dvss.n1421 dvss.n1412 36.1417
R17095 dvss.n1412 dvss.n1353 36.1417
R17096 dvss.n2102 dvss.n1353 36.1417
R17097 dvss.n2102 dvss.n1354 36.1417
R17098 dvss.n1377 dvss.n1354 36.1417
R17099 dvss.n1383 dvss.n1377 36.1417
R17100 dvss.n1383 dvss.n1370 36.1417
R17101 dvss.n1370 dvss.n1366 36.1417
R17102 dvss.n1366 dvss.n1361 36.1417
R17103 dvss.n1361 dvss.n893 36.1417
R17104 dvss.n5728 dvss.n893 36.1417
R17105 dvss.n5728 dvss.n894 36.1417
R17106 dvss.n899 dvss.n894 36.1417
R17107 dvss.n900 dvss.n899 36.1417
R17108 dvss.n904 dvss.n900 36.1417
R17109 dvss.n905 dvss.n904 36.1417
R17110 dvss.n998 dvss.n905 36.1417
R17111 dvss.n998 dvss.n909 36.1417
R17112 dvss.n914 dvss.n909 36.1417
R17113 dvss.n994 dvss.n914 36.1417
R17114 dvss.n997 dvss.n994 36.1417
R17115 dvss.n997 dvss.n920 36.1417
R17116 dvss.n925 dvss.n920 36.1417
R17117 dvss.n926 dvss.n925 36.1417
R17118 dvss.n991 dvss.n926 36.1417
R17119 dvss.n991 dvss.n929 36.1417
R17120 dvss.n934 dvss.n929 36.1417
R17121 dvss.n935 dvss.n934 36.1417
R17122 dvss.n979 dvss.n935 36.1417
R17123 dvss.n1045 dvss.n979 36.1417
R17124 dvss.n1045 dvss.n980 36.1417
R17125 dvss.n980 dvss.n975 36.1417
R17126 dvss.n975 dvss.n944 36.1417
R17127 dvss.n949 dvss.n944 36.1417
R17128 dvss.n950 dvss.n949 36.1417
R17129 dvss.n951 dvss.n950 36.1417
R17130 dvss.n969 dvss.n951 36.1417
R17131 dvss.n1062 dvss.n969 36.1417
R17132 dvss.n1063 dvss.n1062 36.1417
R17133 dvss.n5659 dvss.n1063 36.1417
R17134 dvss.n5659 dvss.n5658 36.1417
R17135 dvss.n5658 dvss.n5657 36.1417
R17136 dvss.n5657 dvss.n1066 36.1417
R17137 dvss.n5651 dvss.n1066 36.1417
R17138 dvss.n5651 dvss.n5650 36.1417
R17139 dvss.n5650 dvss.n5649 36.1417
R17140 dvss.n5649 dvss.n1076 36.1417
R17141 dvss.n1115 dvss.n1076 36.1417
R17142 dvss.n1115 dvss.n1101 36.1417
R17143 dvss.n1105 dvss.n1101 36.1417
R17144 dvss.n1112 dvss.n1105 36.1417
R17145 dvss.n1112 dvss.n1109 36.1417
R17146 dvss.n1109 dvss.n804 36.1417
R17147 dvss.n6123 dvss.n804 36.1417
R17148 dvss.n6123 dvss.n794 36.1417
R17149 dvss.n6156 dvss.n794 36.1417
R17150 dvss.n6156 dvss.n795 36.1417
R17151 dvss.n6132 dvss.n795 36.1417
R17152 dvss.n6138 dvss.n6132 36.1417
R17153 dvss.n6138 dvss.n783 36.1417
R17154 dvss.n6165 dvss.n783 36.1417
R17155 dvss.n6166 dvss.n6165 36.1417
R17156 dvss.n6166 dvss.n779 36.1417
R17157 dvss.n6175 dvss.n779 36.1417
R17158 dvss.n6175 dvss.n775 36.1417
R17159 dvss.n775 dvss.n771 36.1417
R17160 dvss.n771 dvss.n762 36.1417
R17161 dvss.n762 dvss.n530 36.1417
R17162 dvss.n6205 dvss.n530 36.1417
R17163 dvss.n6205 dvss.n531 36.1417
R17164 dvss.n627 dvss.n531 36.1417
R17165 dvss.n635 dvss.n627 36.1417
R17166 dvss.n635 dvss.n615 36.1417
R17167 dvss.n645 dvss.n615 36.1417
R17168 dvss.n645 dvss.n616 36.1417
R17169 dvss.n616 dvss.n611 36.1417
R17170 dvss.n611 dvss.n539 36.1417
R17171 dvss.n544 dvss.n539 36.1417
R17172 dvss.n545 dvss.n544 36.1417
R17173 dvss.n546 dvss.n545 36.1417
R17174 dvss.n550 dvss.n546 36.1417
R17175 dvss.n551 dvss.n550 36.1417
R17176 dvss.n606 dvss.n551 36.1417
R17177 dvss.n606 dvss.n555 36.1417
R17178 dvss.n560 dvss.n555 36.1417
R17179 dvss.n602 dvss.n560 36.1417
R17180 dvss.n605 dvss.n602 36.1417
R17181 dvss.n605 dvss.n566 36.1417
R17182 dvss.n571 dvss.n566 36.1417
R17183 dvss.n572 dvss.n571 36.1417
R17184 dvss.n599 dvss.n572 36.1417
R17185 dvss.n599 dvss.n575 36.1417
R17186 dvss.n580 dvss.n575 36.1417
R17187 dvss.n581 dvss.n580 36.1417
R17188 dvss.n594 dvss.n581 36.1417
R17189 dvss.n596 dvss.n594 36.1417
R17190 dvss.n596 dvss.n589 36.1417
R17191 dvss.n589 dvss.n127 36.1417
R17192 dvss.n6712 dvss.n127 36.1417
R17193 dvss.n6712 dvss.n128 36.1417
R17194 dvss.n133 dvss.n128 36.1417
R17195 dvss.n134 dvss.n133 36.1417
R17196 dvss.n138 dvss.n134 36.1417
R17197 dvss.n139 dvss.n138 36.1417
R17198 dvss.n204 dvss.n139 36.1417
R17199 dvss.n204 dvss.n143 36.1417
R17200 dvss.n148 dvss.n143 36.1417
R17201 dvss.n211 dvss.n148 36.1417
R17202 dvss.n214 dvss.n211 36.1417
R17203 dvss.n214 dvss.n154 36.1417
R17204 dvss.n159 dvss.n154 36.1417
R17205 dvss.n160 dvss.n159 36.1417
R17206 dvss.n181 dvss.n160 36.1417
R17207 dvss.n181 dvss.n163 36.1417
R17208 dvss.n171 dvss.n163 36.1417
R17209 dvss.n172 dvss.n171 36.1417
R17210 dvss.n180 dvss.n172 36.1417
R17211 dvss.n180 dvss.n176 36.1417
R17212 dvss.n176 dvss.n75 36.1417
R17213 dvss.n6864 dvss.n75 36.1417
R17214 dvss.n6864 dvss.n70 36.1417
R17215 dvss.n6897 dvss.n70 36.1417
R17216 dvss.n6897 dvss.n71 36.1417
R17217 dvss.n6873 dvss.n71 36.1417
R17218 dvss.n6879 dvss.n6873 36.1417
R17219 dvss.n6879 dvss.n59 36.1417
R17220 dvss.n6906 dvss.n59 36.1417
R17221 dvss.n6907 dvss.n6906 36.1417
R17222 dvss.n6907 dvss.n55 36.1417
R17223 dvss.n6916 dvss.n55 36.1417
R17224 dvss.n6916 dvss.n51 36.1417
R17225 dvss.n51 dvss.n47 36.1417
R17226 dvss.n47 dvss.n38 36.1417
R17227 dvss.n38 dvss.n28 36.1417
R17228 dvss.n6946 dvss.n28 36.1417
R17229 dvss.n6946 dvss.n29 36.1417
R17230 dvss.n6457 dvss.n29 36.1417
R17231 dvss.n6457 dvss.n6447 36.1417
R17232 dvss.n6469 dvss.n6447 36.1417
R17233 dvss.n6469 dvss.n6443 36.1417
R17234 dvss.n6477 dvss.n6443 36.1417
R17235 dvss.n6477 dvss.n6439 36.1417
R17236 dvss.n6488 dvss.n6439 36.1417
R17237 dvss.n6488 dvss.n6433 36.1417
R17238 dvss.n6496 dvss.n6433 36.1417
R17239 dvss.n6497 dvss.n6496 36.1417
R17240 dvss.n3199 dvss.n3195 36.1417
R17241 dvss.n3204 dvss.n3195 36.1417
R17242 dvss.n3204 dvss.n3191 36.1417
R17243 dvss.n3210 dvss.n3191 36.1417
R17244 dvss.n3210 dvss.n3187 36.1417
R17245 dvss.n3219 dvss.n3187 36.1417
R17246 dvss.n3219 dvss.n3183 36.1417
R17247 dvss.n3226 dvss.n3183 36.1417
R17248 dvss.n3226 dvss.n3177 36.1417
R17249 dvss.n3234 dvss.n3177 36.1417
R17250 dvss.n3234 dvss.n3174 36.1417
R17251 dvss.n3242 dvss.n3174 36.1417
R17252 dvss.n3242 dvss.n3169 36.1417
R17253 dvss.n3250 dvss.n3169 36.1417
R17254 dvss.n3250 dvss.n3166 36.1417
R17255 dvss.n3256 dvss.n3166 36.1417
R17256 dvss.n3256 dvss.n3164 36.1417
R17257 dvss.n3262 dvss.n3164 36.1417
R17258 dvss.n3262 dvss.n3165 36.1417
R17259 dvss.n3165 dvss.n240 36.1417
R17260 dvss.n6635 dvss.n240 36.1417
R17261 dvss.n1703 dvss.n1691 36.1417
R17262 dvss.n1727 dvss.n1703 36.1417
R17263 dvss.n1727 dvss.n1726 36.1417
R17264 dvss.n1726 dvss.n1725 36.1417
R17265 dvss.n1725 dvss.n1724 36.1417
R17266 dvss.n1724 dvss.n1722 36.1417
R17267 dvss.n1722 dvss.n1719 36.1417
R17268 dvss.n1719 dvss.n1718 36.1417
R17269 dvss.n1718 dvss.n1715 36.1417
R17270 dvss.n1715 dvss.n1619 36.1417
R17271 dvss.n1733 dvss.n1619 36.1417
R17272 dvss.n1733 dvss.n1622 36.1417
R17273 dvss.n1622 dvss.n1561 36.1417
R17274 dvss.n1769 dvss.n1561 36.1417
R17275 dvss.n1769 dvss.n1562 36.1417
R17276 dvss.n1586 dvss.n1562 36.1417
R17277 dvss.n1776 dvss.n1555 36.1417
R17278 dvss.n1776 dvss.n1775 36.1417
R17279 dvss.n1775 dvss.n1550 36.1417
R17280 dvss.n1550 dvss.n1545 36.1417
R17281 dvss.n1801 dvss.n1545 36.1417
R17282 dvss.n1802 dvss.n1801 36.1417
R17283 dvss.n1802 dvss.n1540 36.1417
R17284 dvss.n1540 dvss.n1534 36.1417
R17285 dvss.n1824 dvss.n1534 36.1417
R17286 dvss.n1825 dvss.n1824 36.1417
R17287 dvss.n1825 dvss.n1528 36.1417
R17288 dvss.n1837 dvss.n1528 36.1417
R17289 dvss.n1837 dvss.n1518 36.1417
R17290 dvss.n1859 dvss.n1518 36.1417
R17291 dvss.n1859 dvss.n1858 36.1417
R17292 dvss.n1858 dvss.n1521 36.1417
R17293 dvss.n1521 dvss.n1508 36.1417
R17294 dvss.n1871 dvss.n1508 36.1417
R17295 dvss.n1871 dvss.n1494 36.1417
R17296 dvss.n1885 dvss.n1494 36.1417
R17297 dvss.n1885 dvss.n1495 36.1417
R17298 dvss.n1891 dvss.n1489 36.1417
R17299 dvss.n1891 dvss.n1486 36.1417
R17300 dvss.n1899 dvss.n1486 36.1417
R17301 dvss.n1899 dvss.n1482 36.1417
R17302 dvss.n1912 dvss.n1482 36.1417
R17303 dvss.n1912 dvss.n1475 36.1417
R17304 dvss.n1927 dvss.n1475 36.1417
R17305 dvss.n1927 dvss.n1467 36.1417
R17306 dvss.n1936 dvss.n1467 36.1417
R17307 dvss.n1936 dvss.n1462 36.1417
R17308 dvss.n1980 dvss.n1462 36.1417
R17309 dvss.n1980 dvss.n1979 36.1417
R17310 dvss.n1979 dvss.n1464 36.1417
R17311 dvss.n1950 dvss.n1464 36.1417
R17312 dvss.n1966 dvss.n1950 36.1417
R17313 dvss.n1966 dvss.n1965 36.1417
R17314 dvss.n1965 dvss.n1446 36.1417
R17315 dvss.n2026 dvss.n1446 36.1417
R17316 dvss.n2051 dvss.n2026 36.1417
R17317 dvss.n2051 dvss.n2050 36.1417
R17318 dvss.n2050 dvss.n2028 36.1417
R17319 dvss.n2046 dvss.n1436 36.1417
R17320 dvss.n2060 dvss.n1436 36.1417
R17321 dvss.n2060 dvss.n1432 36.1417
R17322 dvss.n2067 dvss.n1432 36.1417
R17323 dvss.n2067 dvss.n1424 36.1417
R17324 dvss.n2080 dvss.n1424 36.1417
R17325 dvss.n2080 dvss.n1414 36.1417
R17326 dvss.n2088 dvss.n1414 36.1417
R17327 dvss.n2088 dvss.n1356 36.1417
R17328 dvss.n2100 dvss.n1356 36.1417
R17329 dvss.n2100 dvss.n2099 36.1417
R17330 dvss.n2099 dvss.n1358 36.1417
R17331 dvss.n1368 dvss.n1358 36.1417
R17332 dvss.n1390 dvss.n1368 36.1417
R17333 dvss.n1390 dvss.n1362 36.1417
R17334 dvss.n1398 dvss.n1362 36.1417
R17335 dvss.n1398 dvss.n896 36.1417
R17336 dvss.n5726 dvss.n896 36.1417
R17337 dvss.n5726 dvss.n5725 36.1417
R17338 dvss.n5725 dvss.n898 36.1417
R17339 dvss.n5721 dvss.n898 36.1417
R17340 dvss.n5720 dvss.n903 36.1417
R17341 dvss.n910 dvss.n903 36.1417
R17342 dvss.n5713 dvss.n910 36.1417
R17343 dvss.n5713 dvss.n5712 36.1417
R17344 dvss.n5712 dvss.n913 36.1417
R17345 dvss.n921 dvss.n913 36.1417
R17346 dvss.n5704 dvss.n921 36.1417
R17347 dvss.n5704 dvss.n5703 36.1417
R17348 dvss.n5703 dvss.n924 36.1417
R17349 dvss.n930 dvss.n924 36.1417
R17350 dvss.n5693 dvss.n930 36.1417
R17351 dvss.n5693 dvss.n5692 36.1417
R17352 dvss.n5692 dvss.n933 36.1417
R17353 dvss.n1042 dvss.n933 36.1417
R17354 dvss.n1043 dvss.n1042 36.1417
R17355 dvss.n1043 dvss.n977 36.1417
R17356 dvss.n977 dvss.n945 36.1417
R17357 dvss.n5677 dvss.n945 36.1417
R17358 dvss.n5677 dvss.n5676 36.1417
R17359 dvss.n5676 dvss.n948 36.1417
R17360 dvss.n5672 dvss.n948 36.1417
R17361 dvss.n5665 dvss.n955 36.1417
R17362 dvss.n5665 dvss.n5664 36.1417
R17363 dvss.n5664 dvss.n5663 36.1417
R17364 dvss.n5663 dvss.n964 36.1417
R17365 dvss.n1088 dvss.n964 36.1417
R17366 dvss.n1090 dvss.n1088 36.1417
R17367 dvss.n1090 dvss.n1089 36.1417
R17368 dvss.n1089 dvss.n1077 36.1417
R17369 dvss.n5647 dvss.n1077 36.1417
R17370 dvss.n5647 dvss.n5646 36.1417
R17371 dvss.n5646 dvss.n1080 36.1417
R17372 dvss.n5639 dvss.n1080 36.1417
R17373 dvss.n5639 dvss.n5638 36.1417
R17374 dvss.n5638 dvss.n1104 36.1417
R17375 dvss.n5626 dvss.n1104 36.1417
R17376 dvss.n5626 dvss.n5625 36.1417
R17377 dvss.n5625 dvss.n796 36.1417
R17378 dvss.n6129 dvss.n796 36.1417
R17379 dvss.n6154 dvss.n6129 36.1417
R17380 dvss.n6154 dvss.n6153 36.1417
R17381 dvss.n6153 dvss.n6131 36.1417
R17382 dvss.n6149 dvss.n786 36.1417
R17383 dvss.n6163 dvss.n786 36.1417
R17384 dvss.n6163 dvss.n782 36.1417
R17385 dvss.n6170 dvss.n782 36.1417
R17386 dvss.n6170 dvss.n774 36.1417
R17387 dvss.n6183 dvss.n774 36.1417
R17388 dvss.n6183 dvss.n764 36.1417
R17389 dvss.n6191 dvss.n764 36.1417
R17390 dvss.n6191 dvss.n533 36.1417
R17391 dvss.n6203 dvss.n533 36.1417
R17392 dvss.n6203 dvss.n6202 36.1417
R17393 dvss.n6202 dvss.n535 36.1417
R17394 dvss.n619 dvss.n535 36.1417
R17395 dvss.n642 dvss.n619 36.1417
R17396 dvss.n643 dvss.n642 36.1417
R17397 dvss.n643 dvss.n613 36.1417
R17398 dvss.n613 dvss.n540 36.1417
R17399 dvss.n754 dvss.n540 36.1417
R17400 dvss.n754 dvss.n753 36.1417
R17401 dvss.n753 dvss.n543 36.1417
R17402 dvss.n749 dvss.n543 36.1417
R17403 dvss.n748 dvss.n549 36.1417
R17404 dvss.n556 dvss.n549 36.1417
R17405 dvss.n741 dvss.n556 36.1417
R17406 dvss.n741 dvss.n740 36.1417
R17407 dvss.n740 dvss.n559 36.1417
R17408 dvss.n567 dvss.n559 36.1417
R17409 dvss.n732 dvss.n567 36.1417
R17410 dvss.n732 dvss.n731 36.1417
R17411 dvss.n731 dvss.n570 36.1417
R17412 dvss.n576 dvss.n570 36.1417
R17413 dvss.n721 dvss.n576 36.1417
R17414 dvss.n721 dvss.n720 36.1417
R17415 dvss.n720 dvss.n579 36.1417
R17416 dvss.n696 dvss.n579 36.1417
R17417 dvss.n696 dvss.n590 36.1417
R17418 dvss.n704 dvss.n590 36.1417
R17419 dvss.n704 dvss.n130 36.1417
R17420 dvss.n6710 dvss.n130 36.1417
R17421 dvss.n6710 dvss.n6709 36.1417
R17422 dvss.n6709 dvss.n132 36.1417
R17423 dvss.n6705 dvss.n132 36.1417
R17424 dvss.n6704 dvss.n137 36.1417
R17425 dvss.n144 dvss.n137 36.1417
R17426 dvss.n6697 dvss.n144 36.1417
R17427 dvss.n6697 dvss.n6696 36.1417
R17428 dvss.n6696 dvss.n147 36.1417
R17429 dvss.n155 dvss.n147 36.1417
R17430 dvss.n6688 dvss.n155 36.1417
R17431 dvss.n6688 dvss.n6687 36.1417
R17432 dvss.n6687 dvss.n158 36.1417
R17433 dvss.n164 dvss.n158 36.1417
R17434 dvss.n6677 dvss.n164 36.1417
R17435 dvss.n6677 dvss.n6676 36.1417
R17436 dvss.n6676 dvss.n167 36.1417
R17437 dvss.n177 dvss.n167 36.1417
R17438 dvss.n6663 dvss.n177 36.1417
R17439 dvss.n6663 dvss.n6662 36.1417
R17440 dvss.n6662 dvss.n72 36.1417
R17441 dvss.n6870 dvss.n72 36.1417
R17442 dvss.n6895 dvss.n6870 36.1417
R17443 dvss.n6895 dvss.n6894 36.1417
R17444 dvss.n6894 dvss.n6872 36.1417
R17445 dvss.n6890 dvss.n62 36.1417
R17446 dvss.n6904 dvss.n62 36.1417
R17447 dvss.n6904 dvss.n58 36.1417
R17448 dvss.n6911 dvss.n58 36.1417
R17449 dvss.n6911 dvss.n50 36.1417
R17450 dvss.n6924 dvss.n50 36.1417
R17451 dvss.n6924 dvss.n40 36.1417
R17452 dvss.n6932 dvss.n40 36.1417
R17453 dvss.n6932 dvss.n31 36.1417
R17454 dvss.n6944 dvss.n31 36.1417
R17455 dvss.n6944 dvss.n6943 36.1417
R17456 dvss.n6943 dvss.n33 36.1417
R17457 dvss.n6462 dvss.n33 36.1417
R17458 dvss.n6462 dvss.n6444 36.1417
R17459 dvss.n6474 dvss.n6444 36.1417
R17460 dvss.n6474 dvss.n6440 36.1417
R17461 dvss.n6482 dvss.n6440 36.1417
R17462 dvss.n6482 dvss.n6435 36.1417
R17463 dvss.n6493 dvss.n6435 36.1417
R17464 dvss.n6493 dvss.n6432 36.1417
R17465 dvss.n6499 dvss.n6432 36.1417
R17466 dvss.n7055 dvss.n0 36.1417
R17467 dvss.n7055 dvss.n7054 36.1417
R17468 dvss.n7054 dvss.n3 36.1417
R17469 dvss.n2287 dvss.n3 36.1417
R17470 dvss.n2287 dvss.n1242 36.1417
R17471 dvss.n2283 dvss.n1242 36.1417
R17472 dvss.n2283 dvss.n2282 36.1417
R17473 dvss.n2282 dvss.n1245 36.1417
R17474 dvss.n2276 dvss.n1245 36.1417
R17475 dvss.n2276 dvss.n2275 36.1417
R17476 dvss.n2275 dvss.n1249 36.1417
R17477 dvss.n2268 dvss.n1249 36.1417
R17478 dvss.n2268 dvss.n2267 36.1417
R17479 dvss.n2267 dvss.n1254 36.1417
R17480 dvss.n2261 dvss.n1254 36.1417
R17481 dvss.n2261 dvss.n2260 36.1417
R17482 dvss.n2256 dvss.n1259 36.1417
R17483 dvss.n2256 dvss.n2255 36.1417
R17484 dvss.n2255 dvss.n1262 36.1417
R17485 dvss.n1265 dvss.n1262 36.1417
R17486 dvss.n2247 dvss.n1265 36.1417
R17487 dvss.n2247 dvss.n2246 36.1417
R17488 dvss.n2246 dvss.n1268 36.1417
R17489 dvss.n2238 dvss.n1268 36.1417
R17490 dvss.n2238 dvss.n2237 36.1417
R17491 dvss.n2237 dvss.n1274 36.1417
R17492 dvss.n2230 dvss.n1274 36.1417
R17493 dvss.n2230 dvss.n2229 36.1417
R17494 dvss.n2229 dvss.n1278 36.1417
R17495 dvss.n1282 dvss.n1278 36.1417
R17496 dvss.n2220 dvss.n1282 36.1417
R17497 dvss.n2220 dvss.n2219 36.1417
R17498 dvss.n2219 dvss.n1285 36.1417
R17499 dvss.n2215 dvss.n1285 36.1417
R17500 dvss.n2215 dvss.n2214 36.1417
R17501 dvss.n2214 dvss.n1288 36.1417
R17502 dvss.n2210 dvss.n1288 36.1417
R17503 dvss.n2210 dvss.n2209 36.1417
R17504 dvss.n2209 dvss.n1291 36.1417
R17505 dvss.n2205 dvss.n1291 36.1417
R17506 dvss.n2205 dvss.n2204 36.1417
R17507 dvss.n2204 dvss.n1294 36.1417
R17508 dvss.n2197 dvss.n1294 36.1417
R17509 dvss.n2197 dvss.n2196 36.1417
R17510 dvss.n2196 dvss.n1299 36.1417
R17511 dvss.n2188 dvss.n1299 36.1417
R17512 dvss.n2188 dvss.n2187 36.1417
R17513 dvss.n2187 dvss.n1305 36.1417
R17514 dvss.n2180 dvss.n1305 36.1417
R17515 dvss.n2180 dvss.n2179 36.1417
R17516 dvss.n2179 dvss.n1309 36.1417
R17517 dvss.n1313 dvss.n1309 36.1417
R17518 dvss.n2170 dvss.n1313 36.1417
R17519 dvss.n2170 dvss.n2169 36.1417
R17520 dvss.n2169 dvss.n1316 36.1417
R17521 dvss.n2160 dvss.n1316 36.1417
R17522 dvss.n2160 dvss.n2159 36.1417
R17523 dvss.n2159 dvss.n1319 36.1417
R17524 dvss.n2155 dvss.n1319 36.1417
R17525 dvss.n2155 dvss.n2154 36.1417
R17526 dvss.n2154 dvss.n1322 36.1417
R17527 dvss.n2150 dvss.n1322 36.1417
R17528 dvss.n2150 dvss.n2149 36.1417
R17529 dvss.n2149 dvss.n1325 36.1417
R17530 dvss.n2142 dvss.n1325 36.1417
R17531 dvss.n2142 dvss.n2141 36.1417
R17532 dvss.n2141 dvss.n1330 36.1417
R17533 dvss.n2133 dvss.n1330 36.1417
R17534 dvss.n2133 dvss.n2132 36.1417
R17535 dvss.n2132 dvss.n1336 36.1417
R17536 dvss.n2125 dvss.n1336 36.1417
R17537 dvss.n2125 dvss.n2124 36.1417
R17538 dvss.n2124 dvss.n1340 36.1417
R17539 dvss.n1345 dvss.n1340 36.1417
R17540 dvss.n2115 dvss.n1345 36.1417
R17541 dvss.n2115 dvss.n885 36.1417
R17542 dvss.n5735 dvss.n885 36.1417
R17543 dvss.n5735 dvss.n878 36.1417
R17544 dvss.n5749 dvss.n878 36.1417
R17545 dvss.n5749 dvss.n879 36.1417
R17546 dvss.n5745 dvss.n879 36.1417
R17547 dvss.n5745 dvss.n5744 36.1417
R17548 dvss.n5744 dvss.n872 36.1417
R17549 dvss.n5756 dvss.n872 36.1417
R17550 dvss.n5756 dvss.n870 36.1417
R17551 dvss.n5765 dvss.n870 36.1417
R17552 dvss.n5765 dvss.n866 36.1417
R17553 dvss.n5771 dvss.n866 36.1417
R17554 dvss.n5771 dvss.n864 36.1417
R17555 dvss.n5783 dvss.n864 36.1417
R17556 dvss.n5783 dvss.n860 36.1417
R17557 dvss.n5789 dvss.n860 36.1417
R17558 dvss.n5789 dvss.n859 36.1417
R17559 dvss.n5797 dvss.n859 36.1417
R17560 dvss.n5797 dvss.n855 36.1417
R17561 dvss.n5803 dvss.n855 36.1417
R17562 dvss.n5803 dvss.n852 36.1417
R17563 dvss.n5818 dvss.n852 36.1417
R17564 dvss.n5818 dvss.n847 36.1417
R17565 dvss.n5826 dvss.n847 36.1417
R17566 dvss.n5826 dvss.n846 36.1417
R17567 dvss.n5831 dvss.n846 36.1417
R17568 dvss.n5831 dvss.n843 36.1417
R17569 dvss.n5837 dvss.n843 36.1417
R17570 dvss.n5837 dvss.n842 36.1417
R17571 dvss.n5843 dvss.n842 36.1417
R17572 dvss.n5843 dvss.n838 36.1417
R17573 dvss.n5849 dvss.n838 36.1417
R17574 dvss.n5849 dvss.n834 36.1417
R17575 dvss.n5858 dvss.n834 36.1417
R17576 dvss.n5858 dvss.n830 36.1417
R17577 dvss.n5865 dvss.n830 36.1417
R17578 dvss.n5865 dvss.n824 36.1417
R17579 dvss.n5873 dvss.n824 36.1417
R17580 dvss.n5873 dvss.n821 36.1417
R17581 dvss.n5880 dvss.n821 36.1417
R17582 dvss.n5880 dvss.n816 36.1417
R17583 dvss.n5888 dvss.n816 36.1417
R17584 dvss.n5888 dvss.n813 36.1417
R17585 dvss.n5894 dvss.n813 36.1417
R17586 dvss.n5894 dvss.n811 36.1417
R17587 dvss.n6116 dvss.n811 36.1417
R17588 dvss.n6116 dvss.n812 36.1417
R17589 dvss.n6112 dvss.n812 36.1417
R17590 dvss.n6112 dvss.n6111 36.1417
R17591 dvss.n6111 dvss.n5904 36.1417
R17592 dvss.n6107 dvss.n5904 36.1417
R17593 dvss.n6107 dvss.n6106 36.1417
R17594 dvss.n6106 dvss.n5907 36.1417
R17595 dvss.n5910 dvss.n5907 36.1417
R17596 dvss.n6098 dvss.n5910 36.1417
R17597 dvss.n6098 dvss.n6097 36.1417
R17598 dvss.n6097 dvss.n5913 36.1417
R17599 dvss.n6089 dvss.n5913 36.1417
R17600 dvss.n6089 dvss.n6088 36.1417
R17601 dvss.n6088 dvss.n5935 36.1417
R17602 dvss.n6081 dvss.n5935 36.1417
R17603 dvss.n6081 dvss.n6080 36.1417
R17604 dvss.n6080 dvss.n5939 36.1417
R17605 dvss.n5943 dvss.n5939 36.1417
R17606 dvss.n6071 dvss.n5943 36.1417
R17607 dvss.n6071 dvss.n6070 36.1417
R17608 dvss.n6070 dvss.n5946 36.1417
R17609 dvss.n6066 dvss.n5946 36.1417
R17610 dvss.n6066 dvss.n6065 36.1417
R17611 dvss.n6065 dvss.n5949 36.1417
R17612 dvss.n6061 dvss.n5949 36.1417
R17613 dvss.n6061 dvss.n6060 36.1417
R17614 dvss.n6060 dvss.n5952 36.1417
R17615 dvss.n6056 dvss.n5952 36.1417
R17616 dvss.n6056 dvss.n6055 36.1417
R17617 dvss.n6055 dvss.n5955 36.1417
R17618 dvss.n6048 dvss.n5955 36.1417
R17619 dvss.n6048 dvss.n6047 36.1417
R17620 dvss.n6047 dvss.n5960 36.1417
R17621 dvss.n6039 dvss.n5960 36.1417
R17622 dvss.n6039 dvss.n6038 36.1417
R17623 dvss.n6038 dvss.n5966 36.1417
R17624 dvss.n6031 dvss.n5966 36.1417
R17625 dvss.n6031 dvss.n6030 36.1417
R17626 dvss.n6030 dvss.n5970 36.1417
R17627 dvss.n5974 dvss.n5970 36.1417
R17628 dvss.n6021 dvss.n5974 36.1417
R17629 dvss.n6021 dvss.n6020 36.1417
R17630 dvss.n6020 dvss.n118 36.1417
R17631 dvss.n6720 dvss.n118 36.1417
R17632 dvss.n6720 dvss.n117 36.1417
R17633 dvss.n6725 dvss.n117 36.1417
R17634 dvss.n6725 dvss.n114 36.1417
R17635 dvss.n6731 dvss.n114 36.1417
R17636 dvss.n6731 dvss.n113 36.1417
R17637 dvss.n6737 dvss.n113 36.1417
R17638 dvss.n6737 dvss.n109 36.1417
R17639 dvss.n6743 dvss.n109 36.1417
R17640 dvss.n6743 dvss.n105 36.1417
R17641 dvss.n6752 dvss.n105 36.1417
R17642 dvss.n6752 dvss.n101 36.1417
R17643 dvss.n6759 dvss.n101 36.1417
R17644 dvss.n6759 dvss.n95 36.1417
R17645 dvss.n6767 dvss.n95 36.1417
R17646 dvss.n6767 dvss.n92 36.1417
R17647 dvss.n6774 dvss.n92 36.1417
R17648 dvss.n6774 dvss.n87 36.1417
R17649 dvss.n6782 dvss.n87 36.1417
R17650 dvss.n6782 dvss.n84 36.1417
R17651 dvss.n6788 dvss.n84 36.1417
R17652 dvss.n6788 dvss.n82 36.1417
R17653 dvss.n6857 dvss.n82 36.1417
R17654 dvss.n6857 dvss.n83 36.1417
R17655 dvss.n6853 dvss.n83 36.1417
R17656 dvss.n6853 dvss.n6852 36.1417
R17657 dvss.n6852 dvss.n6793 36.1417
R17658 dvss.n6848 dvss.n6793 36.1417
R17659 dvss.n6848 dvss.n6847 36.1417
R17660 dvss.n6847 dvss.n6796 36.1417
R17661 dvss.n6799 dvss.n6796 36.1417
R17662 dvss.n6839 dvss.n6799 36.1417
R17663 dvss.n6839 dvss.n6838 36.1417
R17664 dvss.n6838 dvss.n6802 36.1417
R17665 dvss.n6830 dvss.n6802 36.1417
R17666 dvss.n6830 dvss.n6829 36.1417
R17667 dvss.n6829 dvss.n21 36.1417
R17668 dvss.n6953 dvss.n21 36.1417
R17669 dvss.n6953 dvss.n20 36.1417
R17670 dvss.n6965 dvss.n20 36.1417
R17671 dvss.n6965 dvss.n16 36.1417
R17672 dvss.n6971 dvss.n16 36.1417
R17673 dvss.n6971 dvss.n14 36.1417
R17674 dvss.n6978 dvss.n14 36.1417
R17675 dvss.n6978 dvss.n15 36.1417
R17676 dvss.n15 dvss.n10 36.1417
R17677 dvss.n10 dvss.n7 36.1417
R17678 dvss.n6987 dvss.n7 36.1417
R17679 dvss.n5585 dvss.t764 36.0406
R17680 dvss.n2431 dvss.t1204 36.0005
R17681 dvss.n2818 dvss.t376 36.0005
R17682 dvss.n2812 dvss.t769 36.0005
R17683 dvss.n3663 dvss.t2190 36.0005
R17684 dvss.n4198 dvss.t99 36.0005
R17685 dvss.n2260 dvss.n1259 35.7652
R17686 dvss.n6292 dvss.t1477 35.6569
R17687 dvss.n6220 dvss.t1378 35.6569
R17688 dvss.t677 dvss 35.4902
R17689 dvss.t2207 dvss.n7040 35.4058
R17690 dvss.n7040 dvss.t2062 35.4058
R17691 dvss.n4351 dvss.n4331 34.6358
R17692 dvss.n2641 dvss.n2423 34.6358
R17693 dvss.n2939 dvss.n2933 34.6358
R17694 dvss.n2945 dvss.n2944 34.6358
R17695 dvss.n2950 dvss.n2949 34.6358
R17696 dvss.n2949 dvss.n2929 34.6358
R17697 dvss.n2958 dvss.n2957 34.6358
R17698 dvss.n2997 dvss.n2996 34.6358
R17699 dvss.n3005 dvss.n2865 34.6358
R17700 dvss.n3009 dvss.n2865 34.6358
R17701 dvss.n3010 dvss.n3009 34.6358
R17702 dvss.n3012 dvss.n2858 34.6358
R17703 dvss.n3029 dvss.n2858 34.6358
R17704 dvss.n3030 dvss.n3029 34.6358
R17705 dvss.n3031 dvss.n3030 34.6358
R17706 dvss.n3040 dvss.n3039 34.6358
R17707 dvss.n3041 dvss.n3040 34.6358
R17708 dvss.n3047 dvss.n2847 34.6358
R17709 dvss.n3123 dvss.n2847 34.6358
R17710 dvss.n3118 dvss.n3117 34.6358
R17711 dvss.n3425 dvss.n3424 34.6358
R17712 dvss.n2822 dvss.n2821 34.6358
R17713 dvss.n2829 dvss.n2815 34.6358
R17714 dvss.n2825 dvss.n2815 34.6358
R17715 dvss.n2843 dvss.n2806 34.6358
R17716 dvss.n2730 dvss.n2711 34.6358
R17717 dvss.n2736 dvss.n2709 34.6358
R17718 dvss.n2845 dvss.n2686 34.6358
R17719 dvss.n3717 dvss.n3705 34.6358
R17720 dvss.n3734 dvss.n3701 34.6358
R17721 dvss.n3730 dvss.n3701 34.6358
R17722 dvss.n3730 dvss.n3729 34.6358
R17723 dvss.n3729 dvss.n3728 34.6358
R17724 dvss.n3728 dvss.n3703 34.6358
R17725 dvss.n3744 dvss.n3743 34.6358
R17726 dvss.n3743 dvss.n3699 34.6358
R17727 dvss.n3739 dvss.n3699 34.6358
R17728 dvss.n3739 dvss.n3738 34.6358
R17729 dvss.n3752 dvss.n3697 34.6358
R17730 dvss.n3748 dvss.n3697 34.6358
R17731 dvss.n3754 dvss.n3653 34.6358
R17732 dvss.n3687 dvss.n3658 34.6358
R17733 dvss.n3681 dvss.n3662 34.6358
R17734 dvss.n3675 dvss.n3665 34.6358
R17735 dvss.n3786 dvss.n3785 34.6358
R17736 dvss.n3803 dvss.n3802 34.6358
R17737 dvss.n3904 dvss.n3839 34.6358
R17738 dvss.n3900 dvss.n3839 34.6358
R17739 dvss.n3892 dvss.n3891 34.6358
R17740 dvss.n3888 dvss.n3846 34.6358
R17741 dvss.n3883 dvss.n3882 34.6358
R17742 dvss.n3882 dvss.n3849 34.6358
R17743 dvss.n3876 dvss.n3854 34.6358
R17744 dvss.n3872 dvss.n3854 34.6358
R17745 dvss.n3943 dvss.n3917 34.6358
R17746 dvss.n3951 dvss.n3915 34.6358
R17747 dvss.n3947 dvss.n3915 34.6358
R17748 dvss.n3947 dvss.n3946 34.6358
R17749 dvss.n3962 dvss.n3961 34.6358
R17750 dvss.n3961 dvss.n3913 34.6358
R17751 dvss.n3957 dvss.n3913 34.6358
R17752 dvss.n3969 dvss.n3910 34.6358
R17753 dvss.n3965 dvss.n3910 34.6358
R17754 dvss.n3973 dvss.n3464 34.6358
R17755 dvss.n3987 dvss.n3986 34.6358
R17756 dvss.n3986 dvss.n3985 34.6358
R17757 dvss.n3985 dvss.n3462 34.6358
R17758 dvss.n3991 dvss.n3457 34.6358
R17759 dvss.n3483 dvss.n3453 34.6358
R17760 dvss.n3999 dvss.n3453 34.6358
R17761 dvss.n3997 dvss.n3455 34.6358
R17762 dvss.n3549 dvss.n3548 34.6358
R17763 dvss.n3559 dvss.n3558 34.6358
R17764 dvss.n4347 dvss.n4346 34.6358
R17765 dvss.n4426 dvss.n4425 34.6358
R17766 dvss.n4425 dvss.n2397 34.6358
R17767 dvss.n4418 dvss.n2401 34.6358
R17768 dvss.n4299 dvss.n2401 34.6358
R17769 dvss.n4406 dvss.n4299 34.6358
R17770 dvss.n4398 dvss.n4306 34.6358
R17771 dvss.n4732 dvss.n4731 34.6358
R17772 dvss.n4731 dvss.n4730 34.6358
R17773 dvss.n4715 dvss.n4558 34.6358
R17774 dvss.n4574 dvss.n4568 34.6358
R17775 dvss.n4703 dvss.n4577 34.6358
R17776 dvss.n4957 dvss.n4956 34.6358
R17777 dvss.n4956 dvss.n4912 34.6358
R17778 dvss.n4949 dvss.n4915 34.6358
R17779 dvss.n4945 dvss.n4915 34.6358
R17780 dvss.n4933 dvss.n4932 34.6358
R17781 dvss.n5092 dvss.n1218 34.6358
R17782 dvss.n5092 dvss.n5091 34.6358
R17783 dvss.n5088 dvss.n5087 34.6358
R17784 dvss.n5087 dvss.n5086 34.6358
R17785 dvss.n5070 dvss.n5069 34.6358
R17786 dvss.n5067 dvss.n5007 34.6358
R17787 dvss.n5063 dvss.n5062 34.6358
R17788 dvss.n5062 dvss.n5061 34.6358
R17789 dvss.n5061 dvss.n5011 34.6358
R17790 dvss.n5057 dvss.n5011 34.6358
R17791 dvss.n5053 dvss.n5013 34.6358
R17792 dvss.n5046 dvss.n5045 34.6358
R17793 dvss.n5045 dvss.n5015 34.6358
R17794 dvss.n5041 dvss.n5040 34.6358
R17795 dvss.n5040 dvss.n5039 34.6358
R17796 dvss.n4108 dvss.n4107 34.6358
R17797 dvss.n4105 dvss.n4041 34.6358
R17798 dvss.n4077 dvss.n4076 34.6358
R17799 dvss.n4069 dvss.n4058 34.6358
R17800 dvss.n4173 dvss.n4151 34.6358
R17801 dvss.n4287 dvss.n4013 34.6358
R17802 dvss.n4272 dvss.n4271 34.6358
R17803 dvss.n4260 dvss.n4259 34.6358
R17804 dvss.n4259 dvss.n4199 34.6358
R17805 dvss.n4255 dvss.n4199 34.6358
R17806 dvss.n4252 dvss.n4202 34.6358
R17807 dvss.n4247 dvss.n4246 34.6358
R17808 dvss.n4246 dvss.n4204 34.6358
R17809 dvss.n4241 dvss.n4240 34.6358
R17810 dvss.n4235 dvss.n4211 34.6358
R17811 dvss.n4231 dvss.n4211 34.6358
R17812 dvss.n6459 dvss.t1066 34.5917
R17813 dvss.n6651 dvss.t909 34.5917
R17814 dvss.t1559 dvss.n597 34.5917
R17815 dvss.n629 dvss.t1368 34.5917
R17816 dvss.n5615 dvss.t484 34.5917
R17817 dvss.t2159 dvss.n989 34.5917
R17818 dvss.n1380 dvss.t607 34.5917
R17819 dvss.n1954 dvss.t277 34.5917
R17820 dvss.t109 dvss.n1524 34.5917
R17821 dvss.n2707 dvss.t969 34.506
R17822 dvss.n3661 dvss.t167 34.506
R17823 dvss.n3853 dvss.t1434 34.506
R17824 dvss.n3459 dvss.t775 34.506
R17825 dvss.n2388 dvss.t81 34.506
R17826 dvss.n2399 dvss.t83 34.506
R17827 dvss.n4587 dvss.t1387 34.506
R17828 dvss.n4578 dvss.t747 34.506
R17829 dvss.n4585 dvss.t972 34.506
R17830 dvss.n5017 dvss.t1212 34.506
R17831 dvss.n5047 dvss.t2212 34.506
R17832 dvss.n5054 dvss.t943 34.506
R17833 dvss.n1219 dvss.t1109 34.506
R17834 dvss.n4922 dvss.t1032 34.506
R17835 dvss.n4920 dvss.t524 34.506
R17836 dvss.n4043 dvss.t987 34.506
R17837 dvss.n4158 dvss.t2071 34.506
R17838 dvss.n2895 dvss.t2252 34.2973
R17839 dvss.n3355 dvss.t2283 34.2973
R17840 dvss.n3579 dvss.t2241 34.2973
R17841 dvss.n4609 dvss.t2306 34.2973
R17842 dvss.n4684 dvss.t2299 34.2973
R17843 dvss.n2801 dvss.n2797 34.2593
R17844 dvss.n3246 dvss 33.9483
R17845 dvss.n6465 dvss 33.9483
R17846 dvss.n6672 dvss 33.9483
R17847 dvss.n716 dvss 33.9483
R17848 dvss.n638 dvss 33.9483
R17849 dvss.n5635 dvss 33.9483
R17850 dvss.n5688 dvss 33.9483
R17851 dvss.n1386 dvss 33.9483
R17852 dvss.n1975 dvss 33.9483
R17853 dvss.n1843 dvss 33.9483
R17854 dvss.n6962 dvss 33.9483
R17855 dvss.n6778 dvss 33.9483
R17856 dvss.n6026 dvss 33.9483
R17857 dvss.n6076 dvss 33.9483
R17858 dvss.n5884 dvss 33.9483
R17859 dvss.n5807 dvss 33.9483
R17860 dvss.n2120 dvss 33.9483
R17861 dvss.n2175 dvss 33.9483
R17862 dvss.n2225 dvss 33.9483
R17863 dvss.n3034 dvss.n2856 33.8829
R17864 dvss.n2839 dvss.n2838 33.8829
R17865 dvss.n3999 dvss.n3998 33.8829
R17866 dvss.t2152 dvss.t673 33.717
R17867 dvss.t1221 dvss.t1990 33.717
R17868 dvss.t571 dvss.t1931 33.717
R17869 dvss.t626 dvss.t459 33.717
R17870 dvss.t2067 dvss.t1527 33.717
R17871 dvss.t2063 dvss.t1547 33.717
R17872 dvss.t1511 dvss.t1235 33.717
R17873 dvss.t1249 dvss.t1275 33.717
R17874 dvss dvss.t207 33.717
R17875 dvss.t935 dvss.t717 33.717
R17876 dvss.t1197 dvss.t2002 33.717
R17877 dvss.n3970 dvss.n3969 33.5064
R17878 dvss.n3548 dvss.n3534 33.5064
R17879 dvss.n3360 dvss.t2154 33.462
R17880 dvss.n3360 dvss.t1324 33.462
R17881 dvss.n4330 dvss.t2012 33.462
R17882 dvss.n4330 dvss.t1216 33.462
R17883 dvss.n4327 dvss.t1417 33.462
R17884 dvss.n4327 dvss.t635 33.462
R17885 dvss.n4630 dvss.t697 33.462
R17886 dvss.n4630 dvss.t1322 33.462
R17887 dvss.n3119 dvss.n3118 33.1299
R17888 dvss.n3107 dvss.n3057 33.1299
R17889 dvss.n3973 dvss.n3972 33.1299
R17890 dvss.n3796 dvss.n3642 32.7534
R17891 dvss.t1515 dvss.n6357 32.1345
R17892 dvss.n6517 dvss.t1074 32.1345
R17893 dvss.n3869 dvss.n3868 32.0005
R17894 dvss.n3544 dvss.n3543 32.0005
R17895 dvss.n3554 dvss.n3553 32.0005
R17896 dvss.n4432 dvss.n2394 32.0005
R17897 dvss.n4735 dvss.n4547 32.0005
R17898 dvss.n4091 dvss.n4090 32.0005
R17899 dvss.n3815 dvss.n3636 31.624
R17900 dvss.n4107 dvss.n4106 31.624
R17901 dvss.t1305 dvss.n6543 31.6138
R17902 dvss.n3549 dvss.n3533 31.2476
R17903 dvss.t1064 dvss.t1080 31.1326
R17904 dvss.t907 dvss.t1523 31.1326
R17905 dvss.t1563 dvss.t1483 31.1326
R17906 dvss.t1364 dvss.t1384 31.1326
R17907 dvss.t1541 dvss.t486 31.1326
R17908 dvss.t2053 dvss.t2163 31.1326
R17909 dvss.t613 dvss.t514 31.1326
R17910 dvss.t281 dvss.t682 31.1326
R17911 dvss.t44 dvss.t113 31.1326
R17912 dvss.n1123 dvss.t1539 31.0696
R17913 dvss.n2741 dvss.n2708 30.8711
R17914 dvss.n3682 dvss.n3681 30.8711
R17915 dvss.n3878 dvss.n3877 30.8711
R17916 dvss.n4421 dvss.n4420 30.8711
R17917 dvss.n4101 dvss.n4098 30.8711
R17918 dvss.n4261 dvss.n4260 30.8711
R17919 dvss.n3113 dvss.n3112 30.7665
R17920 dvss.n1615 dvss.n1614 30.6481
R17921 dvss.n1251 dvss.n1250 30.6481
R17922 dvss.n2825 dvss.n2824 30.4946
R17923 dvss.n3765 dvss.n3651 30.4946
R17924 dvss.n3769 dvss.n3648 30.4946
R17925 dvss.n3485 dvss.n3484 30.4946
R17926 dvss.n4347 dvss.n4333 30.4946
R17927 dvss.n4023 dvss.t88 30.462
R17928 dvss.n3693 dvss.n3654 30.2506
R17929 dvss.n3777 dvss.n3776 30.1181
R17930 dvss.n4281 dvss.n4017 30.1181
R17931 dvss.n1570 dvss.t40 30.054
R17932 dvss.n2943 dvss.n2933 29.7417
R17933 dvss.n3001 dvss.n2867 29.7417
R17934 dvss.n3724 dvss.n3723 29.7417
R17935 dvss.n3939 dvss.n3938 29.7417
R17936 dvss.n4248 dvss.n4202 29.7417
R17937 dvss.n4242 dvss.n4241 29.7417
R17938 dvss.n4023 dvss.t2016 29.539
R17939 dvss.n2325 dvss.n2306 29.2505
R17940 dvss.n4798 dvss.n2306 29.2505
R17941 dvss.n4802 dvss.n2307 29.2505
R17942 dvss.n4798 dvss.n2307 29.2505
R17943 dvss.n3497 dvss.n3496 28.9887
R17944 dvss.n4950 dvss.n4949 28.9887
R17945 dvss.n4275 dvss.n4021 28.9887
R17946 dvss.n4117 dvss.n4116 28.9609
R17947 dvss.n2432 dvss.t2150 28.7917
R17948 dvss.n3923 dvss.t837 28.7917
R17949 dvss.n3535 dvss.t1190 28.7917
R17950 dvss.n3532 dvss.t548 28.7917
R17951 dvss.n4334 dvss.t2079 28.7917
R17952 dvss.n4610 dvss.t5 28.7917
R17953 dvss.n4546 dvss.t1501 28.7917
R17954 dvss.n4622 dvss.t2231 28.7917
R17955 dvss.n4895 dvss.t1975 28.7917
R17956 dvss.n4900 dvss.t1487 28.7917
R17957 dvss.n4905 dvss.t752 28.7917
R17958 dvss.n4910 dvss.t2087 28.7917
R17959 dvss.n1222 dvss.t1361 28.7917
R17960 dvss.n1227 dvss.t966 28.7917
R17961 dvss.t1519 dvss.n6646 28.7399
R17962 dvss.n6520 dvss.t1078 28.7399
R17963 dvss.n3660 dvss.t94 28.6159
R17964 dvss.n3660 dvss.t2049 28.6159
R17965 dvss.n4216 dvss.t920 28.3801
R17966 dvss.n1230 dvss.t1620 28.3205
R17967 dvss.n1230 dvss.t1641 28.3205
R17968 dvss.n4117 dvss.n4034 28.2358
R17969 dvss.n3129 dvss.t2225 28.1205
R17970 dvss.n6880 dvss.t1430 28.1205
R17971 dvss.n140 dvss.t2059 28.1205
R17972 dvss.n552 dvss.t1974 28.1205
R17973 dvss.n6139 dvss.t1987 28.1205
R17974 dvss.n959 dvss.t479 28.1205
R17975 dvss.n906 dvss.t312 28.1205
R17976 dvss.n2036 dvss.t358 28.1205
R17977 dvss.n1894 dvss.t133 28.1205
R17978 dvss.n1779 dvss.t298 28.1205
R17979 dvss.n6375 dvss.t661 28.1205
R17980 dvss.n6324 dvss.t1447 28.1205
R17981 dvss.n6258 dvss.t676 28.1205
R17982 dvss.n5555 dvss.t765 28.1205
R17983 dvss.n5501 dvss.t894 28.1205
R17984 dvss.n5251 dvss.t2057 28.1205
R17985 dvss.n5212 dvss.t518 28.1205
R17986 dvss.n5173 dvss.t686 28.1205
R17987 dvss.n5134 dvss.t1011 28.1205
R17988 dvss.n2951 dvss.n2950 27.8593
R17989 dvss.n2836 dvss.n2835 27.8593
R17990 dvss.n4726 dvss.n4725 27.8593
R17991 dvss.n3117 dvss.n3051 27.6711
R17992 dvss.n3828 dvss.n3827 27.6711
R17993 dvss.n3013 dvss.n3010 27.4829
R17994 dvss.n3047 dvss.n3046 27.4829
R17995 dvss.n3981 dvss.n3978 27.4829
R17996 dvss.n3566 dvss.n3529 27.4829
R17997 dvss.n4275 dvss.n4274 27.4829
R17998 dvss.n2539 dvss.n2538 27.366
R17999 dvss.n44 dvss.n43 27.2737
R18000 dvss.n222 dvss.n183 27.2737
R18001 dvss.n685 dvss.n684 27.2737
R18002 dvss.n768 dvss.n767 27.2737
R18003 dvss.n1120 dvss.n1119 27.2737
R18004 dvss.n1030 dvss.n1029 27.2737
R18005 dvss.n1418 dvss.n1417 27.2737
R18006 dvss.n1934 dvss.n1471 27.2737
R18007 dvss.n1820 dvss.n1819 27.2737
R18008 dvss.n4932 dvss.n4931 27.2385
R18009 dvss.n5049 dvss.n5013 27.2385
R18010 dvss.n5603 dvss.t1539 27.1069
R18011 dvss.n3112 dvss.n3111 27.1064
R18012 dvss.n3818 dvss.n3816 27.1064
R18013 dvss.n4444 dvss.n2384 27.1064
R18014 dvss.n4404 dvss.n4301 27.1064
R18015 dvss.n4286 dvss.n4285 27.1064
R18016 dvss.n3664 dvss.t1339 26.8576
R18017 dvss.n4057 dvss.t1967 26.8576
R18018 dvss.n4817 dvss.n2304 26.7719
R18019 dvss.n4313 dvss.n4312 26.7039
R18020 dvss.n2627 dvss.n2626 26.6009
R18021 dvss.n3411 dvss.n3340 26.6009
R18022 dvss.n4873 dvss.n4872 26.6009
R18023 dvss.n3224 dvss.t539 26.5065
R18024 dvss.n4448 dvss.n4447 26.314
R18025 dvss.n2962 dvss.n2961 26.314
R18026 dvss.n4352 dvss.n4351 26.314
R18027 dvss.n4636 dvss.n4635 26.314
R18028 dvss.n2835 dvss.n2813 25.977
R18029 dvss.n3612 dvss.n3511 25.977
R18030 dvss.n4236 dvss.n4235 25.977
R18031 dvss.n2535 dvss.t1008 25.9346
R18032 dvss.n2674 dvss.t1218 25.9346
R18033 dvss.n3471 dvss.t1566 25.9346
R18034 dvss.n3465 dvss.t2145 25.9346
R18035 dvss.n3525 dvss.t731 25.9346
R18036 dvss.n4914 dvss.t1485 25.9346
R18037 dvss.n4716 dvss.n4715 25.7355
R18038 dvss.n4872 dvss.n4864 25.7355
R18039 dvss.n4996 dvss.n4995 25.7355
R18040 dvss.n4983 dvss.n4982 25.7355
R18041 dvss.n4970 dvss.n4969 25.7355
R18042 dvss.n4945 dvss.n4944 25.7355
R18043 dvss.n4938 dvss.n4937 25.7355
R18044 dvss.n2631 dvss.n2630 25.6926
R18045 dvss.n3419 dvss.n2680 25.6926
R18046 dvss.n2821 dvss.n2820 25.6926
R18047 dvss.n2794 dvss.n2690 25.6926
R18048 dvss.n3567 dvss.n3566 25.6926
R18049 dvss.n4433 dvss.n4432 25.6926
R18050 dvss.n4676 dvss.n4600 25.6926
R18051 dvss.n5039 dvss.n5019 25.6926
R18052 dvss.n4129 dvss.n4029 25.6926
R18053 dvss.n2563 dvss.n2533 25.6005
R18054 dvss.n2795 dvss.n2794 25.6005
R18055 dvss.n3487 dvss.n3485 25.6005
R18056 dvss.n3492 dvss.n3470 25.6005
R18057 dvss.n3543 dvss.n3536 25.6005
R18058 dvss.n3554 dvss.n3531 25.6005
R18059 dvss.n4342 dvss.n4341 25.6005
R18060 dvss.n5001 dvss.n5000 25.6005
R18061 dvss.n4988 dvss.n4987 25.6005
R18062 dvss.n4975 dvss.n4974 25.6005
R18063 dvss.n4962 dvss.n4961 25.6005
R18064 dvss.n5082 dvss.n5081 25.6005
R18065 dvss.n5076 dvss.n1225 25.6005
R18066 dvss.n4077 dvss.n4053 25.5564
R18067 dvss.n2461 dvss.n2460 25.5168
R18068 dvss.n2341 dvss.n2340 25.5168
R18069 dvss.n5510 dvss.n1145 25.4771
R18070 dvss.n2994 dvss.t1445 25.4291
R18071 dvss.n4937 dvss.n4918 25.3891
R18072 dvss.n5057 dvss.n5056 25.3891
R18073 dvss.t549 dvss.t2128 25.2879
R18074 dvss.t442 dvss.t134 25.2879
R18075 dvss.t152 dvss.t1393 25.2879
R18076 dvss.t742 dvss.t733 25.2879
R18077 dvss.t696 dvss.t2230 25.2879
R18078 dvss.n3775 dvss.n3648 25.224
R18079 dvss.n3776 dvss.n3775 25.224
R18080 dvss.n3615 dvss.n3511 25.224
R18081 dvss.n4121 dvss.n4034 25.224
R18082 dvss.n4122 dvss.n4121 25.224
R18083 dvss.n4065 dvss.n4064 25.224
R18084 dvss.n4281 dvss.n4280 25.224
R18085 dvss.n4280 dvss.n4279 25.224
R18086 dvss.n2527 dvss.n2433 25.1912
R18087 dvss.n2431 dvss.t1010 24.9236
R18088 dvss.n2418 dvss.t882 24.9236
R18089 dvss.n2925 dvss.t564 24.9236
R18090 dvss.n2925 dvss.t562 24.9236
R18091 dvss.n2855 dvss.t1578 24.9236
R18092 dvss.n2855 dvss.t1580 24.9236
R18093 dvss.n2818 dvss.t928 24.9236
R18094 dvss.n2812 dvss.t550 24.9236
R18095 dvss.n3663 dvss.t1045 24.9236
R18096 dvss.n3633 dvss.t1175 24.9236
R18097 dvss.n3979 dvss.t2178 24.9236
R18098 dvss.n3454 dvss.t387 24.9236
R18099 dvss.n3454 dvss.t385 24.9236
R18100 dvss.n3469 dvss.t92 24.9236
R18101 dvss.n3469 dvss.t2018 24.9236
R18102 dvss.n3467 dvss.t2064 24.9236
R18103 dvss.n3467 dvss.t119 24.9236
R18104 dvss.n3517 dvss.t303 24.9236
R18105 dvss.n3517 dvss.t1532 24.9236
R18106 dvss.n4300 dvss.t214 24.9236
R18107 dvss.n4300 dvss.t216 24.9236
R18108 dvss.n4309 dvss.t375 24.9236
R18109 dvss.n4309 dvss.t373 24.9236
R18110 dvss.n4551 dvss.t2124 24.9236
R18111 dvss.n4551 dvss.t797 24.9236
R18112 dvss.n4565 dvss.t2120 24.9236
R18113 dvss.n4565 dvss.t777 24.9236
R18114 dvss.n4602 dvss.t1449 24.9236
R18115 dvss.n4602 dvss.t2116 24.9236
R18116 dvss.n5009 dvss.t788 24.9236
R18117 dvss.n5009 dvss.t1123 24.9236
R18118 dvss.n4048 dvss.t301 24.9236
R18119 dvss.n4048 dvss.t989 24.9236
R18120 dvss.n4198 dvss.t2014 24.9236
R18121 dvss.n378 dvss.t806 24.9236
R18122 dvss.n378 dvss.t808 24.9236
R18123 dvss.n374 dvss.t220 24.9236
R18124 dvss.n374 dvss.t226 24.9236
R18125 dvss.n313 dvss.t1188 24.9236
R18126 dvss.n313 dvss.t1186 24.9236
R18127 dvss.n287 dvss.t69 24.9236
R18128 dvss.n287 dvss.t65 24.9236
R18129 dvss.n286 dvss.t77 24.9236
R18130 dvss.n286 dvss.t71 24.9236
R18131 dvss.n294 dvss.t67 24.9236
R18132 dvss.n294 dvss.t79 24.9236
R18133 dvss.n283 dvss.t73 24.9236
R18134 dvss.n283 dvss.t55 24.9236
R18135 dvss.n303 dvss.t51 24.9236
R18136 dvss.n303 dvss.t57 24.9236
R18137 dvss.n280 dvss.t49 24.9236
R18138 dvss.n280 dvss.t75 24.9236
R18139 dvss.n309 dvss.t59 24.9236
R18140 dvss.n309 dvss.t53 24.9236
R18141 dvss.n382 dvss.t822 24.9236
R18142 dvss.n382 dvss.t824 24.9236
R18143 dvss.n396 dvss.t234 24.9236
R18144 dvss.n396 dvss.t230 24.9236
R18145 dvss.n398 dvss.t242 24.9236
R18146 dvss.n398 dvss.t236 24.9236
R18147 dvss.n393 dvss.t232 24.9236
R18148 dvss.n393 dvss.t244 24.9236
R18149 dvss.n407 dvss.t238 24.9236
R18150 dvss.n407 dvss.t252 24.9236
R18151 dvss.n390 dvss.t248 24.9236
R18152 dvss.n390 dvss.t254 24.9236
R18153 dvss.n387 dvss.t246 24.9236
R18154 dvss.n387 dvss.t240 24.9236
R18155 dvss.n386 dvss.t256 24.9236
R18156 dvss.n386 dvss.t250 24.9236
R18157 dvss.n244 dvss.t802 24.9236
R18158 dvss.n244 dvss.t804 24.9236
R18159 dvss.n258 dvss.t1145 24.9236
R18160 dvss.n258 dvss.t1141 24.9236
R18161 dvss.n260 dvss.t1153 24.9236
R18162 dvss.n260 dvss.t1147 24.9236
R18163 dvss.n255 dvss.t1143 24.9236
R18164 dvss.n255 dvss.t1155 24.9236
R18165 dvss.n269 dvss.t1149 24.9236
R18166 dvss.n269 dvss.t1163 24.9236
R18167 dvss.n252 dvss.t1159 24.9236
R18168 dvss.n252 dvss.t1165 24.9236
R18169 dvss.n249 dvss.t1157 24.9236
R18170 dvss.n249 dvss.t1151 24.9236
R18171 dvss.n248 dvss.t1167 24.9236
R18172 dvss.n248 dvss.t1161 24.9236
R18173 dvss.n346 dvss.t331 24.9236
R18174 dvss.n346 dvss.t325 24.9236
R18175 dvss.n348 dvss.t337 24.9236
R18176 dvss.n348 dvss.t327 24.9236
R18177 dvss.n343 dvss.t339 24.9236
R18178 dvss.n343 dvss.t349 24.9236
R18179 dvss.n357 dvss.t329 24.9236
R18180 dvss.n357 dvss.t341 24.9236
R18181 dvss.n340 dvss.t333 24.9236
R18182 dvss.n340 dvss.t345 24.9236
R18183 dvss.n366 dvss.t355 24.9236
R18184 dvss.n366 dvss.t351 24.9236
R18185 dvss.n337 dvss.t347 24.9236
R18186 dvss.n337 dvss.t343 24.9236
R18187 dvss.n2528 dvss.n2527 24.8476
R18188 dvss.n3039 dvss.n2854 24.8476
R18189 dvss.n3753 dvss.n3752 24.8476
R18190 dvss.n3779 dvss.n3645 24.8476
R18191 dvss.n3827 dvss.n3632 24.8476
R18192 dvss.n3868 dvss.n3859 24.8476
R18193 dvss.n3965 dvss.n3964 24.8476
R18194 dvss.n4346 dvss.n4335 24.8476
R18195 dvss.n4635 dvss.n4623 24.8476
R18196 dvss.n4996 dvss.n4896 24.8476
R18197 dvss.n4983 dvss.n4901 24.8476
R18198 dvss.n4970 dvss.n4906 24.8476
R18199 dvss.n4957 dvss.n4911 24.8476
R18200 dvss.n5086 dvss.n1223 24.8476
R18201 dvss.n5075 dvss.n5074 24.8476
R18202 dvss.n4097 dvss.n4044 24.8476
R18203 dvss.n4267 dvss.n4024 24.8476
R18204 dvss.n4265 dvss.n4196 24.8476
R18205 dvss.n4229 dvss.n4228 24.8476
R18206 dvss.n4226 dvss.n4217 24.8476
R18207 dvss.n4566 dvss.t795 24.6931
R18208 dvss.n4605 dvss.t858 24.6931
R18209 dvss.n5006 dvss.t861 24.6931
R18210 dvss.n4723 dvss.n4722 24.6061
R18211 dvss.n3627 dvss.n3506 24.5331
R18212 dvss.n3423 dvss.n2680 24.4711
R18213 dvss.n3487 dvss.n3472 24.4711
R18214 dvss.n3492 dvss.n3491 24.4711
R18215 dvss.n4443 dvss.n4442 24.4711
R18216 dvss.n4070 dvss.n4069 24.4711
R18217 dvss.n3621 dvss.n3618 24.3205
R18218 dvss.n3688 dvss.n3687 24.3177
R18219 dvss.n3897 dvss.n3896 24.0946
R18220 dvss.n3992 dvss.n3991 24.0946
R18221 dvss.n3491 dvss.n3472 24.0946
R18222 dvss.n3558 dvss.n3531 24.0946
R18223 dvss.n4444 dvss.n4443 24.0946
R18224 dvss.n4506 dvss.n4499 24.0946
R18225 dvss.n5081 dvss.n5080 24.0946
R18226 dvss.n5080 dvss.n1225 24.0946
R18227 dvss.n4227 dvss.n4226 24.0946
R18228 dvss.n2817 dvss.t876 24.0005
R18229 dvss.n4332 dvss.t922 24.0005
R18230 dvss.n2460 dvss.n2457 23.7181
R18231 dvss.n2564 dvss.n2563 23.7181
R18232 dvss.n2990 dvss.n2870 23.7181
R18233 dvss.n2990 dvss.n2869 23.7181
R18234 dvss.n3035 dvss.n3034 23.7181
R18235 dvss.n2830 dvss.n2829 23.7181
R18236 dvss.n2726 dvss.n2711 23.7181
R18237 dvss.n2737 dvss.n2736 23.7181
R18238 dvss.n2743 dvss.n2741 23.7181
R18239 dvss.n3412 dvss.n3411 23.7181
R18240 dvss.n3758 dvss.n3653 23.7181
R18241 dvss.n3758 dvss.n3654 23.7181
R18242 dvss.n3671 dvss.n3669 23.7181
R18243 dvss.n3761 dvss.n3651 23.7181
R18244 dvss.n3905 dvss.n3630 23.7181
R18245 dvss.n3905 dvss.n3904 23.7181
R18246 dvss.n3864 dvss.n3863 23.7181
R18247 dvss.n3977 dvss.n3464 23.7181
R18248 dvss.n3978 dvss.n3977 23.7181
R18249 dvss.n3628 dvss.n3627 23.7181
R18250 dvss.n3616 dvss.n3615 23.7181
R18251 dvss.n3612 dvss.n3611 23.7181
R18252 dvss.n2340 dvss.n2337 23.7181
R18253 dvss.n4442 dvss.n2386 23.7181
R18254 dvss.n4401 dvss.n4400 23.7181
R18255 dvss.n4502 dvss.n4499 23.7181
R18256 dvss.n4736 dvss.n4735 23.7181
R18257 dvss.n4677 dvss.n4676 23.7181
R18258 dvss.n4912 dvss.n1228 23.7181
R18259 dvss.n4951 dvss.n1228 23.7181
R18260 dvss.n5074 dvss.n5004 23.7181
R18261 dvss.n5070 dvss.n5004 23.7181
R18262 dvss.n4093 dvss.n4092 23.7181
R18263 dvss.n4090 dvss.n4051 23.7181
R18264 dvss.n4064 dvss.n4061 23.7181
R18265 dvss.n4267 dvss.n4266 23.7181
R18266 dvss.n4266 dvss.n4265 23.7181
R18267 dvss.n4237 dvss.n4236 23.7181
R18268 dvss.n4222 dvss.n4221 23.7181
R18269 dvss.n4829 dvss.n1233 23.628
R18270 dvss.n5563 dvss.t764 23.613
R18271 dvss.n4811 dvss.t1638 23.5222
R18272 dvss.n1232 dvss.n1229 23.4005
R18273 dvss.n1230 dvss.n1229 23.4005
R18274 dvss.n4853 dvss.n1231 23.4005
R18275 dvss.n1231 dvss.n1230 23.4005
R18276 dvss.n4933 dvss.n4921 23.0907
R18277 dvss.n5055 dvss.n5053 23.0907
R18278 dvss.n2996 dvss.n2995 22.9652
R18279 dvss.n3107 dvss.n3106 22.9652
R18280 dvss.n3723 dvss.n3722 22.9652
R18281 dvss.n3892 dvss.n3844 22.9652
R18282 dvss.n3884 dvss.n3846 22.9652
R18283 dvss.n3938 dvss.n3937 22.9652
R18284 dvss.n3501 dvss.n3468 22.9652
R18285 dvss.n4406 dvss.n4405 22.9652
R18286 dvss.n4308 dvss.n4306 22.9652
R18287 dvss.n4726 dvss.n4552 22.9652
R18288 dvss.n2831 dvss.n2830 22.5887
R18289 dvss.n4179 dvss.n4142 22.5887
R18290 dvss.n4179 dvss.n4178 22.5887
R18291 dvss.n1611 dvss.n1609 22.5639
R18292 dvss.n5115 dvss.n5113 22.5639
R18293 dvss.n3515 dvss.n3514 22.5419
R18294 dvss.n6901 dvss.t1231 22.5415
R18295 dvss.n671 dvss.t365 22.5415
R18296 dvss.n6160 dvss.t778 22.5415
R18297 dvss.n1016 dvss.t14 22.5415
R18298 dvss.n2057 dvss.t1348 22.5415
R18299 dvss.t981 dvss.n1901 22.5415
R18300 dvss.n1792 dvss.t2222 22.5415
R18301 dvss.t1128 dvss.n207 22.5415
R18302 dvss.n5661 dvss.t1295 22.5415
R18303 dvss.n2682 dvss.t450 22.3257
R18304 dvss.n3560 dvss.t2043 22.3257
R18305 dvss.n2642 dvss.n2641 22.2123
R18306 dvss.n3424 dvss.n3423 22.2123
R18307 dvss.n2732 dvss.n2709 22.2123
R18308 dvss.n4065 dvss.n4058 22.2123
R18309 dvss.n2778 dvss.n2777 22.1728
R18310 dvss.n4541 dvss.t2000 22.0959
R18311 dvss.n1565 dvss.t1030 22.0013
R18312 dvss.n1255 dvss.t129 22.0013
R18313 dvss.n2956 dvss.n2955 21.8358
R18314 dvss.n3246 dvss.n3245 21.8222
R18315 dvss.n6465 dvss.n6464 21.8222
R18316 dvss.n6673 dvss.n6672 21.8222
R18317 dvss.n717 dvss.n716 21.8222
R18318 dvss.n638 dvss.n637 21.8222
R18319 dvss.n5636 dvss.n5635 21.8222
R18320 dvss.n5689 dvss.n5688 21.8222
R18321 dvss.n1386 dvss.n1385 21.8222
R18322 dvss.n1976 dvss.n1975 21.8222
R18323 dvss.n1844 dvss.n1843 21.8222
R18324 dvss.n6963 dvss.n6962 21.8222
R18325 dvss.n6778 dvss.n6777 21.8222
R18326 dvss.n6027 dvss.n6026 21.8222
R18327 dvss.n6077 dvss.n6076 21.8222
R18328 dvss.n5884 dvss.n5883 21.8222
R18329 dvss.n5807 dvss.n853 21.8222
R18330 dvss.n2121 dvss.n2120 21.8222
R18331 dvss.n2176 dvss.n2175 21.8222
R18332 dvss.n2226 dvss.n2225 21.8222
R18333 dvss.n4549 dvss.t736 21.795
R18334 dvss.n4556 dvss.t723 21.795
R18335 dvss.n2559 dvss.n2558 21.4593
R18336 dvss.n2995 dvss.n2869 21.4593
R18337 dvss.n3013 dvss.n3012 21.4593
R18338 dvss.n3722 dvss.n3705 21.4593
R18339 dvss.n3717 dvss.n3716 21.4593
R18340 dvss.n3754 dvss.n3753 21.4593
R18341 dvss.n3896 dvss.n3844 21.4593
R18342 dvss.n3884 dvss.n3883 21.4593
R18343 dvss.n3864 dvss.n3859 21.4593
R18344 dvss.n3937 dvss.n3919 21.4593
R18345 dvss.n3993 dvss.n3455 21.4593
R18346 dvss.n3497 dvss.n3468 21.4593
R18347 dvss.n3562 dvss.n3529 21.4593
R18348 dvss.n4405 dvss.n4404 21.4593
R18349 dvss.n4399 dvss.n4398 21.4593
R18350 dvss.n4730 dvss.n4552 21.4593
R18351 dvss.n4703 dvss.n4702 21.4593
R18352 dvss.n4951 dvss.n4950 21.4593
R18353 dvss.n4125 dvss.n4029 21.4593
R18354 dvss.n4093 dvss.n4044 21.4593
R18355 dvss.n4271 dvss.n4024 21.4593
R18356 dvss.n4222 dvss.n4217 21.4593
R18357 dvss.n3585 dvss.n3521 21.3338
R18358 dvss.n3129 dvss.t1038 21.2805
R18359 dvss.n6880 dvss.t740 21.2805
R18360 dvss.n140 dvss.t2196 21.2805
R18361 dvss.n552 dvss.t763 21.2805
R18362 dvss.n6139 dvss.t1989 21.2805
R18363 dvss.n959 dvss.t2194 21.2805
R18364 dvss.n906 dvss.t1254 21.2805
R18365 dvss.n2036 dvss.t2035 21.2805
R18366 dvss.n1894 dvss.t2086 21.2805
R18367 dvss.n1779 dvss.t1041 21.2805
R18368 dvss.n1610 dvss.t399 21.2805
R18369 dvss.n1610 dvss.t398 21.2805
R18370 dvss.n6375 dvss.t1306 21.2805
R18371 dvss.n6324 dvss.t1086 21.2805
R18372 dvss.n6258 dvss.t1320 21.2805
R18373 dvss.n5555 dvss.t767 21.2805
R18374 dvss.n5501 dvss.t1504 21.2805
R18375 dvss.n5251 dvss.t1567 21.2805
R18376 dvss.n5212 dvss.t628 21.2805
R18377 dvss.n5173 dvss.t629 21.2805
R18378 dvss.n5134 dvss.t633 21.2805
R18379 dvss.n5114 dvss.t761 21.2805
R18380 dvss.n5114 dvss.t756 21.2805
R18381 dvss.n3683 dvss.n3658 21.0829
R18382 dvss.n2801 dvss.n2800 21.0829
R18383 dvss.n3787 dvss.n3786 21.0829
R18384 dvss.n3004 dvss.n3001 20.7064
R18385 dvss.n4279 dvss.n4021 20.7064
R18386 dvss.n3302 dvss.t1460 20.507
R18387 dvss.n4923 dvss.n1218 20.4554
R18388 dvss.n5048 dvss.n5046 20.4554
R18389 dvss.n1761 dvss.t552 20.3576
R18390 dvss.n5124 dvss.t1278 20.3576
R18391 dvss.n2627 dvss.n2568 20.3299
R18392 dvss.n2937 dvss.n2870 20.3299
R18393 dvss.n3120 dvss.n2849 20.3299
R18394 dvss.n3767 dvss.n3766 20.3299
R18395 dvss.n4419 dvss.n4418 20.3299
R18396 dvss.n3170 dvss.t1467 20.0005
R18397 dvss.n3170 dvss.t818 20.0005
R18398 dvss.n6449 dvss.t1081 20.0005
R18399 dvss.n6449 dvss.t218 20.0005
R18400 dvss.n174 dvss.t1524 20.0005
R18401 dvss.n174 dvss.t1302 20.0005
R18402 dvss.n583 dvss.t1484 20.0005
R18403 dvss.n583 dvss.t2110 20.0005
R18404 dvss.n622 dvss.t1385 20.0005
R18405 dvss.n622 dvss.t2097 20.0005
R18406 dvss.n1107 dvss.t1542 20.0005
R18407 dvss.n1107 dvss.t1615 20.0005
R18408 dvss.n937 dvss.t2054 20.0005
R18409 dvss.n937 dvss.t1591 20.0005
R18410 dvss.n1371 dvss.t515 20.0005
R18411 dvss.n1371 dvss.t1588 20.0005
R18412 dvss.n1947 dvss.t683 20.0005
R18413 dvss.n1947 dvss.t1603 20.0005
R18414 dvss.n1841 dvss.t45 20.0005
R18415 dvss.n1841 dvss.t2143 20.0005
R18416 dvss.n6957 dvss.t1071 20.0005
R18417 dvss.n6957 dvss.t1327 20.0005
R18418 dvss.n88 dvss.t906 20.0005
R18419 dvss.n88 dvss.t2024 20.0005
R18420 dvss.n5972 dvss.t1558 20.0005
R18421 dvss.n5972 dvss.t1534 20.0005
R18422 dvss.n5941 dvss.t1367 20.0005
R18423 dvss.n5941 dvss.t2108 20.0005
R18424 dvss.n817 dvss.t481 20.0005
R18425 dvss.n817 dvss.t1657 20.0005
R18426 dvss.n854 dvss.t2158 20.0005
R18427 dvss.n854 dvss.t1612 20.0005
R18428 dvss.n1342 dvss.t606 20.0005
R18429 dvss.n1342 dvss.t1609 20.0005
R18430 dvss.n1311 dvss.t272 20.0005
R18431 dvss.n1311 dvss.t1633 20.0005
R18432 dvss.n1280 dvss.t116 20.0005
R18433 dvss.n1280 dvss.t1024 20.0005
R18434 dvss.n3898 dvss.n3897 19.9534
R18435 dvss.n3933 dvss.n3932 19.9534
R18436 dvss.n3618 dvss.n3617 19.9534
R18437 dvss.n4176 dvss.n4175 19.9534
R18438 dvss.n3890 dvss.n3889 19.577
R18439 dvss.n4342 dvss.n4335 19.577
R18440 dvss.n5000 dvss.n4896 19.577
R18441 dvss.n4987 dvss.n4901 19.577
R18442 dvss.n4974 dvss.n4906 19.577
R18443 dvss.n4961 dvss.n4911 19.577
R18444 dvss.n5082 dvss.n1223 19.577
R18445 dvss.n5076 dvss.n5075 19.577
R18446 dvss.n4073 dvss.n4072 19.577
R18447 dvss.n4254 dvss.n4253 19.577
R18448 dvss.n4209 dvss.n4207 19.577
R18449 dvss.n7022 dvss.t1443 19.2955
R18450 dvss.n4106 dvss.n4105 19.2005
R18451 dvss.t535 dvss.n3207 18.9334
R18452 dvss.n972 dvss.n953 18.8324
R18453 dvss.n6900 dvss.n64 18.8324
R18454 dvss.n663 dvss.n662 18.8324
R18455 dvss.n6159 dvss.n788 18.8324
R18456 dvss.n1008 dvss.n1007 18.8324
R18457 dvss.n2056 dvss.n1438 18.8324
R18458 dvss.n1503 dvss.n1491 18.8324
R18459 dvss.n190 dvss.n189 18.8324
R18460 dvss.n2559 dvss.n2533 18.824
R18461 dvss.n2961 dvss.n2923 18.824
R18462 dvss.n3425 dvss.n2678 18.824
R18463 dvss.n2844 dvss.n2843 18.824
R18464 dvss.n3711 dvss.n3652 18.824
R18465 dvss.n4577 dvss.n4576 18.824
R18466 dvss.n1675 dvss.t402 18.6559
R18467 dvss.n1594 dvss.n1557 18.6144
R18468 dvss.n2831 dvss.n2813 18.4476
R18469 dvss.n3677 dvss.n3662 18.4476
R18470 dvss.n6820 dvss.t1101 18.3666
R18471 dvss.n6757 dvss.t1410 18.3666
R18472 dvss.n5932 dvss.t2197 18.3666
R18473 dvss.n6005 dvss.t999 18.3666
R18474 dvss.n5863 dvss.t669 18.3666
R18475 dvss.n5785 dvss.t1115 18.3666
R18476 dvss.t1488 dvss.n1348 18.3666
R18477 dvss.n1986 dvss.t1309 18.3666
R18478 dvss.t261 dvss.n1634 18.3666
R18479 dvss.n4468 dvss.n4467 18.2791
R18480 dvss.n2426 dvss.n2423 18.1815
R18481 dvss.n3816 dvss.n3815 18.0711
R18482 dvss.n3628 dvss.n3466 18.0711
R18483 dvss.n3289 dvss 18.0711
R18484 dvss.n5464 dvss 18.0711
R18485 dvss.n5461 dvss 18.0711
R18486 dvss.n5420 dvss 18.0711
R18487 dvss.n5417 dvss 18.0711
R18488 dvss.n5376 dvss 18.0711
R18489 dvss.n5373 dvss 18.0711
R18490 dvss.n5332 dvss 18.0711
R18491 dvss.n5329 dvss 18.0711
R18492 dvss.n5288 dvss 18.0711
R18493 dvss dvss.n1149 18.0711
R18494 dvss.n5590 dvss 18.0711
R18495 dvss dvss.n5589 18.0711
R18496 dvss.n6248 dvss 18.0711
R18497 dvss dvss.n500 18.0711
R18498 dvss.n6322 dvss 18.0711
R18499 dvss.n6332 dvss 18.0711
R18500 dvss.n6547 dvss 18.0711
R18501 dvss dvss.n6546 18.0711
R18502 dvss.n6505 dvss 18.0711
R18503 dvss.n1586 dvss 18.0711
R18504 dvss.n1495 dvss 18.0711
R18505 dvss dvss.n1489 18.0711
R18506 dvss dvss.n2028 18.0711
R18507 dvss.n2046 dvss 18.0711
R18508 dvss.n5721 dvss 18.0711
R18509 dvss dvss.n5720 18.0711
R18510 dvss.n5672 dvss 18.0711
R18511 dvss.n955 dvss 18.0711
R18512 dvss dvss.n6131 18.0711
R18513 dvss.n6149 dvss 18.0711
R18514 dvss.n749 dvss 18.0711
R18515 dvss dvss.n748 18.0711
R18516 dvss.n6705 dvss 18.0711
R18517 dvss dvss.n6704 18.0711
R18518 dvss dvss.n6872 18.0711
R18519 dvss.n6890 dvss 18.0711
R18520 dvss.n6499 dvss 18.0711
R18521 dvss.n7011 dvss.t1651 18.0005
R18522 dvss.n4823 dvss.t1599 17.7798
R18523 dvss.n2932 dvss.n2929 17.6946
R18524 dvss.n3041 dvss.n2852 17.6946
R18525 dvss.n3748 dvss.n3747 17.6946
R18526 dvss.n3871 dvss.n3870 17.6946
R18527 dvss.n3957 dvss.n3956 17.6946
R18528 dvss.n3461 dvss.n3460 17.6946
R18529 dvss.n4428 dvss.n4427 17.6946
R18530 dvss.n4101 dvss.n4100 17.6946
R18531 dvss dvss.n1555 17.6946
R18532 dvss.n421 dvss.t649 17.4005
R18533 dvss.n421 dvss.t1585 17.4005
R18534 dvss.n423 dvss.t820 17.4005
R18535 dvss.n423 dvss.t653 17.4005
R18536 dvss.n7005 dvss.t2022 17.4005
R18537 dvss.n7005 dvss.t1618 17.4005
R18538 dvss.n7004 dvss.t530 17.4005
R18539 dvss.n7004 dvss.t1678 17.4005
R18540 dvss.n7003 dvss.t2020 17.4005
R18541 dvss.n7003 dvss.t292 17.4005
R18542 dvss.n7011 dvss.t296 17.4005
R18543 dvss.n6998 dvss.t1675 17.4005
R18544 dvss.n6998 dvss.t2100 17.4005
R18545 dvss.n3712 dvss.n3707 17.3181
R18546 dvss.n3617 dvss.n3616 17.3181
R18547 dvss.n4598 dvss.n4597 17.2527
R18548 dvss.n6639 dvss.n236 17.2441
R18549 dvss.n7033 dvss.n7032 17.1002
R18550 dvss.n2551 dvss.n2540 16.9936
R18551 dvss.n4386 dvss.n4314 16.9936
R18552 dvss.n4386 dvss.n4385 16.9936
R18553 dvss.n2529 dvss.n2429 16.9417
R18554 dvss.n3046 dvss.n3044 16.9417
R18555 dvss.n3870 dvss.n3869 16.9417
R18556 dvss.n3981 dvss.n3462 16.9417
R18557 dvss.n4428 dvss.n2394 16.9417
R18558 dvss.n4228 dvss.n4227 16.9417
R18559 dvss.n7034 dvss.n7033 16.9365
R18560 dvss.t1007 dvss.t647 16.8587
R18561 dvss.t2006 dvss.t833 16.8587
R18562 dvss.t1531 dvss.t1694 16.8587
R18563 dvss.t2209 dvss.t1972 16.8587
R18564 dvss.t792 dvss.t1948 16.8587
R18565 dvss.t383 dvss.t2184 16.8587
R18566 dvss.n2724 dvss.n2723 16.8353
R18567 dvss.t1462 dvss.n3309 16.8072
R18568 dvss.n4695 dvss.n4694 16.7924
R18569 dvss.n2167 dvss.n2166 16.666
R18570 dvss.n884 dvss.n883 16.6189
R18571 dvss.n5816 dvss.n5815 16.6189
R18572 dvss.n3097 dvss.n3065 16.6166
R18573 dvss.n1453 dvss.n1452 16.615
R18574 dvss.n986 dvss.n985 16.615
R18575 dvss.n803 dvss.n802 16.611
R18576 dvss.n1404 dvss.n1403 16.6032
R18577 dvss.n5900 dvss.n5899 16.5915
R18578 dvss.n2558 dvss.n2557 16.5652
R18579 dvss.n4124 dvss.n4123 16.5652
R18580 dvss.n2552 dvss.n2551 16.5522
R18581 dvss.n4845 dvss.t1660 16.5305
R18582 dvss.n4845 dvss.t1645 16.5305
R18583 dvss.n4832 dvss.t1648 16.5305
R18584 dvss.n4832 dvss.t1636 16.5305
R18585 dvss.n4836 dvss.t1669 16.5305
R18586 dvss.n4836 dvss.t1621 16.5305
R18587 dvss.n4840 dvss.t1642 16.5305
R18588 dvss.n4840 dvss.t1627 16.5305
R18589 dvss.n2313 dvss.t1624 16.5305
R18590 dvss.n2313 dvss.t1672 16.5305
R18591 dvss.n2314 dvss.t1663 16.5305
R18592 dvss.n2314 dvss.t1594 16.5305
R18593 dvss.n2308 dvss.t1597 16.5305
R18594 dvss.n2308 dvss.t1630 16.5305
R18595 dvss.n7025 dvss.n6996 16.3843
R18596 dvss.n296 dvss.n293 16.3561
R18597 dvss.n300 dvss.n284 16.3561
R18598 dvss.n305 dvss.n302 16.3561
R18599 dvss.n327 dvss.n326 16.3561
R18600 dvss.n323 dvss.n322 16.3561
R18601 dvss.n319 dvss.n318 16.3561
R18602 dvss.n318 dvss.n317 16.3561
R18603 dvss.n266 dvss.n256 16.3561
R18604 dvss.n271 dvss.n268 16.3561
R18605 dvss.n275 dvss.n253 16.3561
R18606 dvss.n6619 dvss.n6618 16.3561
R18607 dvss.n6624 dvss.n6622 16.3561
R18608 dvss.n6628 dvss.n245 16.3561
R18609 dvss.n6629 dvss.n6628 16.3561
R18610 dvss.n219 dvss.n218 16.2674
R18611 dvss.n1118 dvss.n1117 16.2674
R18612 dvss.n6930 dvss.n45 16.2668
R18613 dvss.n683 dvss.n600 16.2668
R18614 dvss.n6189 dvss.n769 16.2668
R18615 dvss.n1028 dvss.n992 16.2668
R18616 dvss.n2086 dvss.n1419 16.2668
R18617 dvss.n1931 dvss.n1930 16.2668
R18618 dvss.n1818 dvss.n1817 16.2668
R18619 dvss.n2732 dvss.n2731 16.1887
R18620 dvss.n3766 dvss.n3765 16.1887
R18621 dvss.n3785 dvss.n3645 16.1887
R18622 dvss.n4287 dvss.n4286 16.1887
R18623 dvss.n291 dvss.n288 16.1783
R18624 dvss.n262 dvss.n259 16.1783
R18625 dvss.n4490 dvss.n4489 16.1689
R18626 dvss.n5523 dvss.t1543 16.1564
R18627 dvss.n404 dvss.n394 16.132
R18628 dvss.n409 dvss.n406 16.132
R18629 dvss.n413 dvss.n391 16.132
R18630 dvss.n444 dvss.n443 16.132
R18631 dvss.n449 dvss.n447 16.132
R18632 dvss.n453 dvss.n383 16.132
R18633 dvss.n454 dvss.n453 16.132
R18634 dvss.t759 dvss.n1570 16.1286
R18635 dvss.n1685 dvss.t1035 15.9908
R18636 dvss.n400 dvss.n397 15.9567
R18637 dvss.n2506 dvss.n2505 15.849
R18638 dvss.n329 dvss.n328 15.8227
R18639 dvss.n6617 dvss.n6616 15.8227
R18640 dvss.n2958 dvss.n2923 15.8123
R18641 dvss.n2780 dvss.n2694 15.8123
R18642 dvss.n2845 dvss.n2844 15.8123
R18643 dvss.n3502 dvss.n3466 15.8123
R18644 dvss.n333 dvss.n332 15.6449
R18645 dvss.n6613 dvss.n6612 15.6449
R18646 dvss.n442 dvss.n441 15.606
R18647 dvss.n2557 dvss.n2556 15.5708
R18648 dvss.n3822 dvss.n3634 15.4358
R18649 dvss.n3502 dvss.n3501 15.4358
R18650 dvss.n2643 dvss.n2642 15.3963
R18651 dvss.n3365 dvss.n3364 15.3963
R18652 dvss.n4737 dvss.n4736 15.3963
R18653 dvss.n5002 dvss.n4857 15.3963
R18654 dvss.n317 dvss.n314 15.2894
R18655 dvss.n6630 dvss.n6629 15.2894
R18656 dvss.n4989 dvss.n4988 15.1944
R18657 dvss.n4976 dvss.n4975 15.1944
R18658 dvss.n4963 dvss.n4962 15.1944
R18659 dvss.n3430 dvss.n3429 15.1514
R18660 dvss.n2723 dvss.n2712 15.1259
R18661 dvss.n455 dvss.n454 15.08
R18662 dvss.n3670 dvss.n3665 15.0593
R18663 dvss.n3801 dvss.n3800 15.0593
R18664 dvss.n4073 dvss.n4054 15.0593
R18665 dvss.n4072 dvss.n4071 15.0593
R18666 dvss.n2553 dvss.n2538 15.0266
R18667 dvss.n319 dvss.n311 14.9338
R18668 dvss.n6623 dvss.n245 14.9338
R18669 dvss.n5032 dvss.n5031 14.8179
R18670 dvss.n3413 dvss.n3412 14.775
R18671 dvss.n4191 dvss.n4025 14.775
R18672 dvss.n4191 dvss.n4026 14.775
R18673 dvss.n4183 dvss.n4142 14.775
R18674 dvss.n448 dvss.n383 14.7293
R18675 dvss.n354 dvss.n344 14.7205
R18676 dvss.n359 dvss.n356 14.7205
R18677 dvss.n363 dvss.n341 14.7205
R18678 dvss.n368 dvss.n365 14.7205
R18679 dvss.n6602 dvss.n338 14.7205
R18680 dvss.n6598 dvss.n6597 14.7205
R18681 dvss.n6594 dvss.n6593 14.7205
R18682 dvss.n6593 dvss.n6592 14.7205
R18683 dvss.n6589 dvss.n6588 14.7205
R18684 dvss.n6585 dvss.n6584 14.7205
R18685 dvss.n6584 dvss.n6583 14.7205
R18686 dvss.n2944 dvss.n2943 14.6829
R18687 dvss.n2997 dvss.n2867 14.6829
R18688 dvss.n3761 dvss.n3652 14.6829
R18689 dvss.n3712 dvss.n3711 14.6829
R18690 dvss.n3724 dvss.n3703 14.6829
R18691 dvss.n3933 dvss.n3919 14.6829
R18692 dvss.n3939 dvss.n3917 14.6829
R18693 dvss.n4576 dvss.n4575 14.6829
R18694 dvss.n4248 dvss.n4247 14.6829
R18695 dvss.n4242 dvss.n4204 14.6829
R18696 dvss.n2610 dvss.n2609 14.5992
R18697 dvss.n350 dvss.n347 14.5605
R18698 dvss.n438 dvss.n437 14.5539
R18699 dvss.n3106 dvss.n3105 14.4946
R18700 dvss.n2630 dvss.n2568 14.3064
R18701 dvss.n3123 dvss.n2849 14.3064
R18702 dvss.n3770 dvss.n3767 14.3064
R18703 dvss.n3823 dvss.n3822 14.3064
R18704 dvss.n4420 dvss.n4419 14.3064
R18705 dvss.n4255 dvss.n4254 14.3064
R18706 dvss.n4237 dvss.n4209 14.3064
R18707 dvss.n2482 dvss.n2447 14.2735
R18708 dvss.n2590 dvss.n2589 14.2735
R18709 dvss.n3077 dvss.n3076 14.2735
R18710 dvss.n2360 dvss.n2326 14.2735
R18711 dvss.n329 dvss.n281 14.0449
R18712 dvss.n326 dvss.n310 14.0449
R18713 dvss.n6616 dvss.n250 14.0449
R18714 dvss.n6619 dvss.n246 14.0449
R18715 dvss.n3877 dvss.n3876 13.9299
R18716 dvss.n4421 dvss.n2397 13.9299
R18717 dvss.n4098 dvss.n4097 13.9299
R18718 dvss.n4162 dvss.n4159 13.9299
R18719 dvss.n441 dvss.n388 13.8526
R18720 dvss.n444 dvss.n384 13.8526
R18721 dvss.n3622 dvss.n3621 13.8383
R18722 dvss.n3835 dvss.n3834 13.8253
R18723 dvss.n6592 dvss.n375 13.7605
R18724 dvss.n7049 dvss.n6995 13.7086
R18725 dvss.n292 dvss.n291 13.6894
R18726 dvss.n262 dvss.n261 13.6894
R18727 dvss.n5542 dvss.t1545 13.6709
R18728 dvss.n2938 dvss.n2937 13.5534
R18729 dvss.n2839 dvss.n2809 13.5534
R18730 dvss.n3788 dvss.n3787 13.5534
R18731 dvss.n400 dvss.n399 13.5019
R18732 dvss.n6594 dvss.n372 13.4405
R18733 dvss.n6585 dvss.n376 13.4405
R18734 dvss.n7031 dvss.n7025 13.3982
R18735 dvss.n6583 dvss.n379 13.2077
R18736 dvss.n2564 dvss.n2429 13.177
R18737 dvss.n3928 dvss.n3927 13.177
R18738 dvss.n3539 dvss.n3536 13.177
R18739 dvss.n4341 dvss.n4340 13.177
R18740 dvss.n4629 dvss.n4628 13.177
R18741 dvss.n4631 dvss.n4629 13.177
R18742 dvss.n5002 dvss.n5001 13.177
R18743 dvss.n4125 dvss.n4124 13.177
R18744 dvss.n4177 dvss.n4176 13.177
R18745 dvss.n6813 dvss.t1097 13.1192
R18746 dvss.t1406 dvss.n6740 13.1192
R18747 dvss.n5925 dvss.t2199 13.1192
R18748 dvss.t997 dvss.n5999 13.1192
R18749 dvss.t667 dvss.n5846 13.1192
R18750 dvss.n5753 dvss.t1119 13.1192
R18751 dvss.n2011 dvss.t1494 13.1192
R18752 dvss.n1642 dvss.t1315 13.1192
R18753 dvss.n1669 dvss.t267 13.1192
R18754 dvss.n7031 dvss.n7030 13.0828
R18755 dvss.n2884 dvss.n2881 12.8005
R18756 dvss.n2957 dvss.n2956 12.8005
R18757 dvss.n2719 dvss.n2718 12.8005
R18758 dvss.n3716 dvss.n3707 12.8005
R18759 dvss.n4677 dvss.n4599 12.8005
R18760 dvss.n367 dvss.n336 12.6405
R18761 dvss.n371 dvss.n338 12.6405
R18762 dvss.n4657 dvss.n4611 12.5658
R18763 dvss.n3246 dvss.n3173 12.5222
R18764 dvss.n6465 dvss.n6454 12.5222
R18765 dvss.n6672 dvss.n173 12.5222
R18766 dvss.n716 dvss.n582 12.5222
R18767 dvss.n638 dvss.n625 12.5222
R18768 dvss.n5635 dvss.n1106 12.5222
R18769 dvss.n5688 dvss.n936 12.5222
R18770 dvss.n1386 dvss.n1375 12.5222
R18771 dvss.n1975 dvss.n1946 12.5222
R18772 dvss.n1843 dvss.n1840 12.5222
R18773 dvss.n6962 dvss.n6956 12.5222
R18774 dvss.n6778 dvss.n91 12.5222
R18775 dvss.n6026 dvss.n5971 12.5222
R18776 dvss.n6076 dvss.n5940 12.5222
R18777 dvss.n5884 dvss.n820 12.5222
R18778 dvss.n5808 dvss.n5807 12.5222
R18779 dvss.n2120 dvss.n1341 12.5222
R18780 dvss.n2175 dvss.n1310 12.5222
R18781 dvss.n2225 dvss.n1279 12.5222
R18782 dvss.n3928 dvss.n3922 12.424
R18783 dvss.n350 dvss.n349 12.3205
R18784 dvss.n2743 dvss.n2706 12.285
R18785 dvss.n1612 dvss.n1611 12.2361
R18786 dvss.n5116 dvss.n5115 12.2361
R18787 dvss.t517 dvss.t754 12.1889
R18788 dvss.n1616 dvss.n1615 12.1422
R18789 dvss.n2272 dvss.n1251 12.1422
R18790 dvss.n3586 dvss.n3585 12.1268
R18791 dvss.n4400 dvss.n4399 12.0476
R18792 dvss.t754 dvss.t1277 11.8304
R18793 dvss.n2784 dvss.n2694 11.7632
R18794 dvss.n2800 dvss.n2799 11.6711
R18795 dvss.n4161 dvss.n4013 11.6711
R18796 dvss.n218 dvss.t1132 11.3667
R18797 dvss.n1118 dvss.t1297 11.3667
R18798 dvss.t1225 dvss.n45 11.3663
R18799 dvss.n683 dvss.t367 11.3663
R18800 dvss.t786 dvss.n769 11.3663
R18801 dvss.n1028 dvss.t10 11.3663
R18802 dvss.t1342 dvss.n1419 11.3663
R18803 dvss.n1930 dvss.t975 11.3663
R18804 dvss.n1818 dvss.t2216 11.3663
R18805 dvss.n3802 dvss.n3801 11.2946
R18806 dvss.n304 dvss.n279 11.2005
R18807 dvss.n277 dvss.n276 11.2005
R18808 dvss.n4817 dvss.n4816 11.1237
R18809 dvss.n415 dvss.n414 11.0471
R18810 dvss.n3429 dvss.n2678 10.9181
R18811 dvss.n3388 dvss.n3387 10.9091
R18812 dvss.n296 dvss.n295 10.8449
R18813 dvss.n267 dvss.n266 10.8449
R18814 dvss.n6581 dvss.n379 10.7826
R18815 dvss.n2719 dvss.n2714 10.7135
R18816 dvss.n2726 dvss.n2725 10.7135
R18817 dvss.n3611 dvss.n3512 10.7135
R18818 dvss.n405 dvss.n404 10.6964
R18819 dvss.n3272 dvss.t1459 10.6405
R18820 dvss.n3272 dvss.t1463 10.6405
R18821 dvss.n3276 dvss.t1465 10.6405
R18822 dvss.n3276 dvss.t1461 10.6405
R18823 dvss.n3180 dvss.t532 10.6405
R18824 dvss.n3180 dvss.t540 10.6405
R18825 dvss.n3189 dvss.t536 10.6405
R18826 dvss.n3189 dvss.t534 10.6405
R18827 dvss.n36 dvss.t1228 10.6405
R18828 dvss.n36 dvss.t1226 10.6405
R18829 dvss.n53 dvss.t1232 10.6405
R18830 dvss.n53 dvss.t1230 10.6405
R18831 dvss.n152 dvss.t1127 10.6405
R18832 dvss.n152 dvss.t1133 10.6405
R18833 dvss.n150 dvss.t1129 10.6405
R18834 dvss.n150 dvss.t1125 10.6405
R18835 dvss.n564 dvss.t364 10.6405
R18836 dvss.n564 dvss.t368 10.6405
R18837 dvss.n562 dvss.t366 10.6405
R18838 dvss.n562 dvss.t360 10.6405
R18839 dvss.n760 dvss.t783 10.6405
R18840 dvss.n760 dvss.t787 10.6405
R18841 dvss.n777 dvss.t779 10.6405
R18842 dvss.n777 dvss.t785 10.6405
R18843 dvss.n1094 dvss.t1292 10.6405
R18844 dvss.n1094 dvss.t1298 10.6405
R18845 dvss.n1083 dvss.t1296 10.6405
R18846 dvss.n1083 dvss.t1300 10.6405
R18847 dvss.n918 dvss.t9 10.6405
R18848 dvss.n918 dvss.t11 10.6405
R18849 dvss.n916 dvss.t15 10.6405
R18850 dvss.n916 dvss.t13 10.6405
R18851 dvss.n1410 dvss.t1345 10.6405
R18852 dvss.n1410 dvss.t1343 10.6405
R18853 dvss.n1427 dvss.t1349 10.6405
R18854 dvss.n1427 dvss.t1347 10.6405
R18855 dvss.n1921 dvss.t978 10.6405
R18856 dvss.n1921 dvss.t976 10.6405
R18857 dvss.n1907 dvss.t982 10.6405
R18858 dvss.n1907 dvss.t980 10.6405
R18859 dvss.n1806 dvss.t2219 10.6405
R18860 dvss.n1806 dvss.t2217 10.6405
R18861 dvss.n1783 dvss.t2223 10.6405
R18862 dvss.n1783 dvss.t2221 10.6405
R18863 dvss.n35 dvss.t1069 10.6405
R18864 dvss.n35 dvss.t1067 10.6405
R18865 dvss.n6450 dvss.t1065 10.6405
R18866 dvss.n6450 dvss.t1063 10.6405
R18867 dvss.n168 dvss.t912 10.6405
R18868 dvss.n168 dvss.t910 10.6405
R18869 dvss.n6666 dvss.t908 10.6405
R18870 dvss.n6666 dvss.t904 10.6405
R18871 dvss.n587 dvss.t1562 10.6405
R18872 dvss.n587 dvss.t1560 10.6405
R18873 dvss.n710 dvss.t1564 10.6405
R18874 dvss.n710 dvss.t1556 10.6405
R18875 dvss.n759 dvss.t1373 10.6405
R18876 dvss.n759 dvss.t1369 10.6405
R18877 dvss.n536 dvss.t1365 10.6405
R18878 dvss.n536 dvss.t1363 10.6405
R18879 dvss.n5642 dvss.t489 10.6405
R18880 dvss.n5642 dvss.t485 10.6405
R18881 dvss.n5629 dvss.t487 10.6405
R18882 dvss.n5629 dvss.t483 10.6405
R18883 dvss.n941 dvss.t2166 10.6405
R18884 dvss.n941 dvss.t2160 10.6405
R18885 dvss.n5682 dvss.t2164 10.6405
R18886 dvss.n5682 dvss.t2168 10.6405
R18887 dvss.n1409 dvss.t610 10.6405
R18888 dvss.n1409 dvss.t608 10.6405
R18889 dvss.n1359 dvss.t614 10.6405
R18890 dvss.n1359 dvss.t616 10.6405
R18891 dvss.n1465 dvss.t274 10.6405
R18892 dvss.n1465 dvss.t278 10.6405
R18893 dvss.n1969 dvss.t282 10.6405
R18894 dvss.n1969 dvss.t280 10.6405
R18895 dvss.n1512 dvss.t106 10.6405
R18896 dvss.n1512 dvss.t110 10.6405
R18897 dvss.n1515 dvss.t114 10.6405
R18898 dvss.n1515 dvss.t108 10.6405
R18899 dvss.n6412 dvss.t1083 10.6405
R18900 dvss.n6412 dvss.t1079 10.6405
R18901 dvss.n6416 dvss.t1077 10.6405
R18902 dvss.n6416 dvss.t1075 10.6405
R18903 dvss.n6561 dvss.t1522 10.6405
R18904 dvss.n6561 dvss.t1520 10.6405
R18905 dvss.n6346 dvss.t1518 10.6405
R18906 dvss.n6346 dvss.t1516 10.6405
R18907 dvss.n481 dvss.t1480 10.6405
R18908 dvss.n481 dvss.t1478 10.6405
R18909 dvss.n484 dvss.t1482 10.6405
R18910 dvss.n484 dvss.t1476 10.6405
R18911 dvss.n510 dvss.t1383 10.6405
R18912 dvss.n510 dvss.t1379 10.6405
R18913 dvss.n513 dvss.t1377 10.6405
R18914 dvss.n513 dvss.t1375 10.6405
R18915 dvss.n1137 dvss.t1544 10.6405
R18916 dvss.n1137 dvss.t1538 10.6405
R18917 dvss.n5532 dvss.t1540 10.6405
R18918 dvss.n5532 dvss.t1536 10.6405
R18919 dvss.n5271 dvss.t2055 10.6405
R18920 dvss.n5271 dvss.t2050 10.6405
R18921 dvss.n5275 dvss.t2052 10.6405
R18922 dvss.n5275 dvss.t2056 10.6405
R18923 dvss.n5232 dvss.t511 10.6405
R18924 dvss.n5232 dvss.t510 10.6405
R18925 dvss.n5236 dvss.t513 10.6405
R18926 dvss.n5236 dvss.t516 10.6405
R18927 dvss.n5193 dvss.t679 10.6405
R18928 dvss.n5193 dvss.t681 10.6405
R18929 dvss.n5197 dvss.t685 10.6405
R18930 dvss.n5197 dvss.t684 10.6405
R18931 dvss.n5154 dvss.t41 10.6405
R18932 dvss.n5154 dvss.t43 10.6405
R18933 dvss.n5158 dvss.t47 10.6405
R18934 dvss.n5158 dvss.t42 10.6405
R18935 dvss.n6804 dvss.t1104 10.6405
R18936 dvss.n6804 dvss.t1102 10.6405
R18937 dvss.n6797 dvss.t1098 10.6405
R18938 dvss.n6797 dvss.t1106 10.6405
R18939 dvss.n98 dvss.t1415 10.6405
R18940 dvss.n98 dvss.t1411 10.6405
R18941 dvss.n107 dvss.t1407 10.6405
R18942 dvss.n107 dvss.t1413 10.6405
R18943 dvss.n5962 dvss.t1006 10.6405
R18944 dvss.n5962 dvss.t1000 10.6405
R18945 dvss.n5956 dvss.t998 10.6405
R18946 dvss.n5956 dvss.t1002 10.6405
R18947 dvss.n5915 dvss.t2204 10.6405
R18948 dvss.n5915 dvss.t2198 10.6405
R18949 dvss.n5908 dvss.t2200 10.6405
R18950 dvss.n5908 dvss.t2206 10.6405
R18951 dvss.n827 dvss.t664 10.6405
R18952 dvss.n827 dvss.t670 10.6405
R18953 dvss.n836 dvss.t668 10.6405
R18954 dvss.n836 dvss.t672 10.6405
R18955 dvss.n5776 dvss.t1114 10.6405
R18956 dvss.n5776 dvss.t1116 10.6405
R18957 dvss.n5760 dvss.t1120 10.6405
R18958 dvss.n5760 dvss.t1118 10.6405
R18959 dvss.n1332 dvss.t1491 10.6405
R18960 dvss.n1332 dvss.t1489 10.6405
R18961 dvss.n1326 dvss.t1495 10.6405
R18962 dvss.n1326 dvss.t1493 10.6405
R18963 dvss.n1301 dvss.t1312 10.6405
R18964 dvss.n1301 dvss.t1310 10.6405
R18965 dvss.n1295 dvss.t1316 10.6405
R18966 dvss.n1295 dvss.t1314 10.6405
R18967 dvss.n1270 dvss.t264 10.6405
R18968 dvss.n1270 dvss.t262 10.6405
R18969 dvss.n1263 dvss.t268 10.6405
R18970 dvss.n1263 dvss.t266 10.6405
R18971 dvss.n3201 dvss.n3190 10.64
R18972 dvss.n6909 dvss.n54 10.64
R18973 dvss.n151 dvss.n149 10.64
R18974 dvss.n563 dvss.n561 10.64
R18975 dvss.n6168 dvss.n778 10.64
R18976 dvss.n1084 dvss.n1082 10.64
R18977 dvss.n917 dvss.n915 10.64
R18978 dvss.n2065 dvss.n1428 10.64
R18979 dvss.n1908 dvss.n1906 10.64
R18980 dvss.n1788 dvss.n1787 10.64
R18981 dvss.n6844 dvss.n6843 10.64
R18982 dvss.n6734 dvss.n108 10.64
R18983 dvss.n6053 dvss.n6052 10.64
R18984 dvss.n6103 dvss.n6102 10.64
R18985 dvss.n5840 dvss.n837 10.64
R18986 dvss.n5761 dvss.n5759 10.64
R18987 dvss.n2147 dvss.n2146 10.64
R18988 dvss.n2202 dvss.n2201 10.64
R18989 dvss.n2252 dvss.n2251 10.64
R18990 dvss.n7036 dvss.n7018 10.6369
R18991 dvss.n7040 dvss.n7018 10.6369
R18992 dvss.n7039 dvss.n7038 10.6369
R18993 dvss.n7040 dvss.n7039 10.6369
R18994 dvss.n7016 dvss.n7015 10.6369
R18995 dvss.n7019 dvss.n7016 10.6369
R18996 dvss.n7045 dvss.n7002 10.6369
R18997 dvss.n7019 dvss.n7002 10.6369
R18998 dvss.n2885 dvss.n2884 10.5983
R18999 dvss.n315 dvss.n314 10.3672
R19000 dvss.n6631 dvss.n6630 10.3672
R19001 dvss.n456 dvss.n455 10.3526
R19002 dvss.n3005 dvss.n3004 10.1652
R19003 dvss.n4071 dvss.n4070 10.1652
R19004 dvss.n365 dvss.n364 10.0805
R19005 dvss.n6605 dvss.t346 10.0615
R19006 dvss.n5091 dvss.n1220 10.0265
R19007 dvss.n5018 dvss.n5015 10.0265
R19008 dvss.n3780 dvss.n3779 9.78874
R19009 dvss.n4262 dvss.n4196 9.78874
R19010 dvss.n1209 dvss.n241 9.76206
R19011 dvss.n355 dvss.n354 9.7605
R19012 dvss.n4865 dvss 9.74003
R19013 dvss.n5026 dvss.n5025 9.71789
R19014 dvss.n3561 dvss.n3559 9.41227
R19015 dvss.n4567 dvss.n4558 9.41227
R19016 dvss.n5069 dvss.n5068 9.41227
R19017 dvss.n2755 dvss.n2753 9.36527
R19018 dvss.t1659 dvss.n1145 9.32101
R19019 dvss.n3334 dvss 9.31486
R19020 dvss dvss.n3199 9.31486
R19021 dvss.n5493 dvss 9.31486
R19022 dvss dvss.n0 9.30735
R19023 dvss.n3581 dvss.n3521 9.30134
R19024 dvss.n1699 dvss.n1698 9.30085
R19025 dvss.n2591 dvss.n2590 9.3005
R19026 dvss.n2593 dvss.n2592 9.3005
R19027 dvss.n2594 dvss.n2584 9.3005
R19028 dvss.n2596 dvss.n2595 9.3005
R19029 dvss.n2598 dvss.n2597 9.3005
R19030 dvss.n2599 dvss.n2582 9.3005
R19031 dvss.n2601 dvss.n2600 9.3005
R19032 dvss.n2602 dvss.n2581 9.3005
R19033 dvss.n2604 dvss.n2603 9.3005
R19034 dvss.n2605 dvss.n2580 9.3005
R19035 dvss.n2607 dvss.n2606 9.3005
R19036 dvss.n2609 dvss.n2608 9.3005
R19037 dvss.n2460 dvss.n2459 9.3005
R19038 dvss.n2462 dvss.n2461 9.3005
R19039 dvss.n2464 dvss.n2463 9.3005
R19040 dvss.n2465 dvss.n2453 9.3005
R19041 dvss.n2467 dvss.n2466 9.3005
R19042 dvss.n2468 dvss.n2452 9.3005
R19043 dvss.n2470 dvss.n2469 9.3005
R19044 dvss.n2471 dvss.n2451 9.3005
R19045 dvss.n2473 dvss.n2472 9.3005
R19046 dvss.n2475 dvss.n2474 9.3005
R19047 dvss.n2476 dvss.n2449 9.3005
R19048 dvss.n2479 dvss.n2478 9.3005
R19049 dvss.n2480 dvss.n2447 9.3005
R19050 dvss.n2482 dvss.n2481 9.3005
R19051 dvss.n2484 dvss.n2446 9.3005
R19052 dvss.n2488 dvss.n2487 9.3005
R19053 dvss.n2490 dvss.n2489 9.3005
R19054 dvss.n2492 dvss.n2491 9.3005
R19055 dvss.n2494 dvss.n2493 9.3005
R19056 dvss.n2495 dvss.n2443 9.3005
R19057 dvss.n2497 dvss.n2496 9.3005
R19058 dvss.n2499 dvss.n2498 9.3005
R19059 dvss.n2500 dvss.n2441 9.3005
R19060 dvss.n2503 dvss.n2502 9.3005
R19061 dvss.n2505 dvss.n2504 9.3005
R19062 dvss.n2507 dvss.n2506 9.3005
R19063 dvss.n2509 dvss.n2508 9.3005
R19064 dvss.n2510 dvss.n2438 9.3005
R19065 dvss.n2512 dvss.n2511 9.3005
R19066 dvss.n2513 dvss.n2437 9.3005
R19067 dvss.n2515 dvss.n2514 9.3005
R19068 dvss.n2516 dvss.n2436 9.3005
R19069 dvss.n2518 dvss.n2517 9.3005
R19070 dvss.n2520 dvss.n2519 9.3005
R19071 dvss.n2521 dvss.n2434 9.3005
R19072 dvss.n2524 dvss.n2523 9.3005
R19073 dvss.n2525 dvss.n2433 9.3005
R19074 dvss.n2527 dvss.n2526 9.3005
R19075 dvss.n2528 dvss.n2430 9.3005
R19076 dvss.n2530 dvss.n2529 9.3005
R19077 dvss.n2531 dvss.n2429 9.3005
R19078 dvss.n2564 dvss.n2532 9.3005
R19079 dvss.n2563 dvss.n2562 9.3005
R19080 dvss.n2561 dvss.n2533 9.3005
R19081 dvss.n2560 dvss.n2559 9.3005
R19082 dvss.n2558 dvss.n2534 9.3005
R19083 dvss.n2557 dvss.n2536 9.3005
R19084 dvss.n2556 dvss 9.3005
R19085 dvss.n2555 dvss.n2554 9.3005
R19086 dvss.n2551 dvss.n2550 9.3005
R19087 dvss.n2548 dvss.n2547 9.3005
R19088 dvss.n2545 dvss.n2411 9.3005
R19089 dvss.n2415 dvss.n2412 9.3005
R19090 dvss.n2653 dvss.n2652 9.3005
R19091 dvss.n2651 dvss.n2650 9.3005
R19092 dvss.n2649 dvss.n2648 9.3005
R19093 dvss.n2647 dvss.n2417 9.3005
R19094 dvss.n2646 dvss.n2645 9.3005
R19095 dvss.n2644 dvss.n2643 9.3005
R19096 dvss.n2642 dvss.n2422 9.3005
R19097 dvss.n2641 dvss.n2640 9.3005
R19098 dvss.n2639 dvss.n2423 9.3005
R19099 dvss.n2638 dvss.n2637 9.3005
R19100 dvss.n2635 dvss.n2424 9.3005
R19101 dvss.n2634 dvss.n2633 9.3005
R19102 dvss.n2632 dvss.n2631 9.3005
R19103 dvss.n2630 dvss.n2629 9.3005
R19104 dvss.n2628 dvss.n2627 9.3005
R19105 dvss.n2626 dvss.n2625 9.3005
R19106 dvss.n2624 dvss.n2623 9.3005
R19107 dvss.n2622 dvss.n2570 9.3005
R19108 dvss.n2621 dvss.n2620 9.3005
R19109 dvss.n2619 dvss.n2571 9.3005
R19110 dvss.n2618 dvss.n2617 9.3005
R19111 dvss.n2616 dvss.n2572 9.3005
R19112 dvss.n2615 dvss.n2614 9.3005
R19113 dvss.n2613 dvss.n2612 9.3005
R19114 dvss.n3078 dvss.n3077 9.3005
R19115 dvss.n3080 dvss.n3079 9.3005
R19116 dvss.n3081 dvss.n3071 9.3005
R19117 dvss.n3083 dvss.n3082 9.3005
R19118 dvss.n3085 dvss.n3084 9.3005
R19119 dvss.n3086 dvss.n3069 9.3005
R19120 dvss.n3088 dvss.n3087 9.3005
R19121 dvss.n3089 dvss.n3068 9.3005
R19122 dvss.n3091 dvss.n3090 9.3005
R19123 dvss.n3092 dvss.n3066 9.3005
R19124 dvss.n3094 dvss.n3093 9.3005
R19125 dvss.n3095 dvss.n3065 9.3005
R19126 dvss.n2884 dvss.n2883 9.3005
R19127 dvss.n2886 dvss.n2878 9.3005
R19128 dvss.n2889 dvss.n2888 9.3005
R19129 dvss.n2890 dvss.n2877 9.3005
R19130 dvss.n2892 dvss.n2891 9.3005
R19131 dvss.n2893 dvss.n2875 9.3005
R19132 dvss.n2899 dvss.n2898 9.3005
R19133 dvss.n2901 dvss.n2900 9.3005
R19134 dvss.n2904 dvss.n2903 9.3005
R19135 dvss.n2906 dvss.n2905 9.3005
R19136 dvss.n2907 dvss.n2872 9.3005
R19137 dvss.n2910 dvss.n2909 9.3005
R19138 dvss.n2911 dvss.n2871 9.3005
R19139 dvss.n2987 dvss.n2912 9.3005
R19140 dvss.n2986 dvss.n2985 9.3005
R19141 dvss.n2984 dvss.n2913 9.3005
R19142 dvss.n2983 dvss.n2982 9.3005
R19143 dvss.n2981 dvss.n2914 9.3005
R19144 dvss.n2980 dvss.n2979 9.3005
R19145 dvss.n2978 dvss.n2977 9.3005
R19146 dvss.n2976 dvss.n2975 9.3005
R19147 dvss.n2974 dvss.n2973 9.3005
R19148 dvss.n2971 dvss.n2919 9.3005
R19149 dvss.n2969 dvss.n2968 9.3005
R19150 dvss.n2967 dvss.n2920 9.3005
R19151 dvss.n2966 dvss.n2965 9.3005
R19152 dvss.n2962 dvss.n2921 9.3005
R19153 dvss.n2961 dvss.n2960 9.3005
R19154 dvss.n2959 dvss.n2958 9.3005
R19155 dvss.n2957 dvss.n2924 9.3005
R19156 dvss.n2955 dvss.n2954 9.3005
R19157 dvss.n2953 dvss.n2952 9.3005
R19158 dvss.n2950 dvss.n2928 9.3005
R19159 dvss.n2949 dvss.n2948 9.3005
R19160 dvss.n2947 dvss.n2929 9.3005
R19161 dvss.n2946 dvss.n2945 9.3005
R19162 dvss.n2944 dvss.n2930 9.3005
R19163 dvss.n2943 dvss.n2942 9.3005
R19164 dvss.n2941 dvss.n2933 9.3005
R19165 dvss.n2940 dvss.n2939 9.3005
R19166 dvss.n2934 dvss.n2870 9.3005
R19167 dvss.n2991 dvss.n2990 9.3005
R19168 dvss.n2992 dvss.n2869 9.3005
R19169 dvss.n2995 dvss.n2993 9.3005
R19170 dvss.n2996 dvss.n2868 9.3005
R19171 dvss.n2998 dvss.n2997 9.3005
R19172 dvss.n2999 dvss.n2867 9.3005
R19173 dvss.n3001 dvss.n3000 9.3005
R19174 dvss.n3004 dvss.n2866 9.3005
R19175 dvss.n3006 dvss.n3005 9.3005
R19176 dvss.n3007 dvss.n2865 9.3005
R19177 dvss.n3009 dvss.n3008 9.3005
R19178 dvss.n3010 dvss.n2864 9.3005
R19179 dvss.n3014 dvss.n3013 9.3005
R19180 dvss.n3012 dvss.n2863 9.3005
R19181 dvss.n3020 dvss.n2858 9.3005
R19182 dvss.n3029 dvss.n3028 9.3005
R19183 dvss.n3030 dvss.n2857 9.3005
R19184 dvss.n3032 dvss.n3031 9.3005
R19185 dvss.n3034 dvss.n3033 9.3005
R19186 dvss.n3036 dvss.n3035 9.3005
R19187 dvss.n3037 dvss.n2854 9.3005
R19188 dvss.n3039 dvss.n3038 9.3005
R19189 dvss.n3040 dvss.n2853 9.3005
R19190 dvss.n3042 dvss.n3041 9.3005
R19191 dvss.n3044 dvss.n3043 9.3005
R19192 dvss.n3046 dvss.n2850 9.3005
R19193 dvss.n3048 dvss.n3047 9.3005
R19194 dvss.n3049 dvss.n2847 9.3005
R19195 dvss.n3123 dvss.n3122 9.3005
R19196 dvss.n3121 dvss.n3120 9.3005
R19197 dvss.n3118 dvss.n3050 9.3005
R19198 dvss.n3117 dvss.n3116 9.3005
R19199 dvss.n3115 dvss.n3051 9.3005
R19200 dvss.n3114 dvss.n3113 9.3005
R19201 dvss.n3112 dvss.n3052 9.3005
R19202 dvss.n3110 dvss.n3109 9.3005
R19203 dvss.n3108 dvss.n3107 9.3005
R19204 dvss.n3106 dvss.n3058 9.3005
R19205 dvss.n3105 dvss.n3104 9.3005
R19206 dvss.n3103 dvss.n3102 9.3005
R19207 dvss.n3100 dvss.n3061 9.3005
R19208 dvss.n3097 dvss.n3096 9.3005
R19209 dvss.n3365 dvss.n3359 9.3005
R19210 dvss.n3368 dvss.n3367 9.3005
R19211 dvss.n3369 dvss.n3358 9.3005
R19212 dvss.n3371 dvss.n3370 9.3005
R19213 dvss.n3373 dvss.n3357 9.3005
R19214 dvss.n3375 dvss.n3374 9.3005
R19215 dvss.n3376 dvss.n3356 9.3005
R19216 dvss.n3378 dvss.n3377 9.3005
R19217 dvss.n3354 dvss.n3353 9.3005
R19218 dvss.n3384 dvss.n3383 9.3005
R19219 dvss.n3386 dvss.n3385 9.3005
R19220 dvss.n3352 dvss.n3350 9.3005
R19221 dvss.n2720 dvss.n2719 9.3005
R19222 dvss.n2727 dvss.n2726 9.3005
R19223 dvss.n2728 dvss.n2711 9.3005
R19224 dvss.n2730 dvss.n2729 9.3005
R19225 dvss.n2733 dvss.n2732 9.3005
R19226 dvss.n2734 dvss.n2709 9.3005
R19227 dvss.n2736 dvss.n2735 9.3005
R19228 dvss.n2738 dvss.n2737 9.3005
R19229 dvss.n2739 dvss.n2708 9.3005
R19230 dvss.n2741 dvss.n2740 9.3005
R19231 dvss.n2744 dvss.n2743 9.3005
R19232 dvss.n2746 dvss.n2745 9.3005
R19233 dvss.n2748 dvss.n2705 9.3005
R19234 dvss.n2751 dvss.n2750 9.3005
R19235 dvss.n2753 dvss.n2752 9.3005
R19236 dvss.n2758 dvss.n2757 9.3005
R19237 dvss.n2759 dvss.n2703 9.3005
R19238 dvss.n2761 dvss.n2760 9.3005
R19239 dvss.n2762 dvss.n2702 9.3005
R19240 dvss.n2764 dvss.n2763 9.3005
R19241 dvss.n2766 dvss.n2765 9.3005
R19242 dvss.n2767 dvss.n2699 9.3005
R19243 dvss.n2769 dvss.n2768 9.3005
R19244 dvss.n2771 dvss.n2770 9.3005
R19245 dvss.n2772 dvss.n2697 9.3005
R19246 dvss.n2775 dvss.n2774 9.3005
R19247 dvss.n2777 dvss.n2776 9.3005
R19248 dvss.n2778 dvss.n2695 9.3005
R19249 dvss.n2781 dvss.n2780 9.3005
R19250 dvss.n2782 dvss.n2694 9.3005
R19251 dvss.n2784 dvss.n2783 9.3005
R19252 dvss.n2786 dvss.n2691 9.3005
R19253 dvss.n2792 dvss.n2791 9.3005
R19254 dvss.n2793 dvss.n2690 9.3005
R19255 dvss.n2794 dvss 9.3005
R19256 dvss.n2796 dvss.n2687 9.3005
R19257 dvss.n2802 dvss.n2801 9.3005
R19258 dvss.n2803 dvss.n2686 9.3005
R19259 dvss.n2845 dvss.n2804 9.3005
R19260 dvss.n2843 dvss.n2842 9.3005
R19261 dvss.n2841 dvss.n2806 9.3005
R19262 dvss.n2840 dvss.n2839 9.3005
R19263 dvss.n2837 dvss.n2807 9.3005
R19264 dvss.n2835 dvss.n2834 9.3005
R19265 dvss.n2833 dvss.n2813 9.3005
R19266 dvss.n2832 dvss.n2831 9.3005
R19267 dvss.n2830 dvss.n2814 9.3005
R19268 dvss.n2829 dvss.n2828 9.3005
R19269 dvss.n2827 dvss.n2815 9.3005
R19270 dvss.n2826 dvss.n2825 9.3005
R19271 dvss.n2822 dvss.n2816 9.3005
R19272 dvss.n2821 dvss.n2670 9.3005
R19273 dvss.n2820 dvss.n2671 9.3005
R19274 dvss.n3435 dvss.n3434 9.3005
R19275 dvss.n3433 dvss.n3432 9.3005
R19276 dvss.n3431 dvss.n3430 9.3005
R19277 dvss.n3429 dvss.n3428 9.3005
R19278 dvss.n3427 dvss.n2678 9.3005
R19279 dvss.n3426 dvss.n3425 9.3005
R19280 dvss.n3424 dvss.n2679 9.3005
R19281 dvss.n3423 dvss.n3422 9.3005
R19282 dvss.n3421 dvss.n2680 9.3005
R19283 dvss.n3420 dvss.n3419 9.3005
R19284 dvss.n3417 dvss.n3416 9.3005
R19285 dvss.n3415 dvss.n2681 9.3005
R19286 dvss.n3414 dvss.n3413 9.3005
R19287 dvss.n3412 dvss.n3339 9.3005
R19288 dvss.n3411 dvss.n3410 9.3005
R19289 dvss.n3409 dvss.n3340 9.3005
R19290 dvss.n3408 dvss.n3407 9.3005
R19291 dvss.n3405 dvss.n3341 9.3005
R19292 dvss.n3404 dvss.n3403 9.3005
R19293 dvss.n3402 dvss.n3401 9.3005
R19294 dvss.n3400 dvss.n3344 9.3005
R19295 dvss.n3399 dvss.n3398 9.3005
R19296 dvss.n3397 dvss.n3396 9.3005
R19297 dvss.n3394 dvss.n3347 9.3005
R19298 dvss.n3393 dvss.n3392 9.3005
R19299 dvss.n3391 dvss.n3390 9.3005
R19300 dvss.n3388 dvss.n3349 9.3005
R19301 dvss.n3672 dvss.n3671 9.3005
R19302 dvss.n3673 dvss.n3665 9.3005
R19303 dvss.n3675 dvss.n3674 9.3005
R19304 dvss.n3678 dvss.n3677 9.3005
R19305 dvss.n3679 dvss.n3662 9.3005
R19306 dvss.n3681 dvss.n3680 9.3005
R19307 dvss.n3682 dvss.n3659 9.3005
R19308 dvss.n3684 dvss.n3683 9.3005
R19309 dvss.n3685 dvss.n3658 9.3005
R19310 dvss.n3687 dvss.n3686 9.3005
R19311 dvss.n3688 dvss.n3655 9.3005
R19312 dvss.n3694 dvss.n3693 9.3005
R19313 dvss.n3695 dvss.n3654 9.3005
R19314 dvss.n3758 dvss.n3757 9.3005
R19315 dvss.n3756 dvss.n3653 9.3005
R19316 dvss.n3755 dvss.n3754 9.3005
R19317 dvss.n3753 dvss.n3696 9.3005
R19318 dvss.n3752 dvss.n3751 9.3005
R19319 dvss.n3750 dvss.n3697 9.3005
R19320 dvss.n3749 dvss.n3748 9.3005
R19321 dvss.n3744 dvss.n3698 9.3005
R19322 dvss.n3743 dvss.n3742 9.3005
R19323 dvss.n3741 dvss.n3699 9.3005
R19324 dvss.n3740 dvss.n3739 9.3005
R19325 dvss.n3738 dvss.n3700 9.3005
R19326 dvss.n3734 dvss.n3733 9.3005
R19327 dvss.n3732 dvss.n3701 9.3005
R19328 dvss.n3731 dvss.n3730 9.3005
R19329 dvss.n3729 dvss.n3702 9.3005
R19330 dvss.n3728 dvss.n3727 9.3005
R19331 dvss.n3726 dvss.n3703 9.3005
R19332 dvss.n3725 dvss.n3724 9.3005
R19333 dvss.n3723 dvss.n3704 9.3005
R19334 dvss.n3722 dvss.n3720 9.3005
R19335 dvss.n3719 dvss.n3705 9.3005
R19336 dvss.n3718 dvss.n3717 9.3005
R19337 dvss.n3716 dvss.n3715 9.3005
R19338 dvss.n3714 dvss.n3707 9.3005
R19339 dvss.n3713 dvss.n3712 9.3005
R19340 dvss.n3711 dvss.n3710 9.3005
R19341 dvss.n3709 dvss.n3652 9.3005
R19342 dvss.n3762 dvss.n3761 9.3005
R19343 dvss.n3763 dvss.n3651 9.3005
R19344 dvss.n3765 dvss.n3764 9.3005
R19345 dvss.n3766 dvss.n3649 9.3005
R19346 dvss.n3771 dvss.n3770 9.3005
R19347 dvss.n3772 dvss.n3648 9.3005
R19348 dvss.n3775 dvss.n3773 9.3005
R19349 dvss.n3776 dvss.n3646 9.3005
R19350 dvss.n3781 dvss.n3780 9.3005
R19351 dvss.n3782 dvss.n3645 9.3005
R19352 dvss.n3785 dvss.n3783 9.3005
R19353 dvss.n3786 dvss.n3643 9.3005
R19354 dvss.n3789 dvss.n3788 9.3005
R19355 dvss.n3796 dvss.n3795 9.3005
R19356 dvss.n3804 dvss.n3803 9.3005
R19357 dvss.n3802 dvss.n3637 9.3005
R19358 dvss.n3812 dvss.n3636 9.3005
R19359 dvss.n3815 dvss.n3813 9.3005
R19360 dvss.n3816 dvss.n3635 9.3005
R19361 dvss.n3819 dvss.n3818 9.3005
R19362 dvss.n3820 dvss.n3634 9.3005
R19363 dvss.n3822 dvss.n3821 9.3005
R19364 dvss.n3824 dvss.n3823 9.3005
R19365 dvss.n3825 dvss.n3632 9.3005
R19366 dvss.n3827 dvss.n3826 9.3005
R19367 dvss.n3828 dvss.n3631 9.3005
R19368 dvss.n3836 dvss.n3835 9.3005
R19369 dvss.n3837 dvss.n3630 9.3005
R19370 dvss.n3905 dvss.n3838 9.3005
R19371 dvss.n3904 dvss.n3903 9.3005
R19372 dvss.n3902 dvss.n3839 9.3005
R19373 dvss.n3901 dvss.n3900 9.3005
R19374 dvss.n3898 dvss.n3840 9.3005
R19375 dvss.n3897 dvss.n3842 9.3005
R19376 dvss.n3896 dvss.n3895 9.3005
R19377 dvss.n3894 dvss.n3844 9.3005
R19378 dvss.n3893 dvss.n3892 9.3005
R19379 dvss.n3891 dvss.n3845 9.3005
R19380 dvss.n3888 dvss.n3887 9.3005
R19381 dvss.n3886 dvss.n3846 9.3005
R19382 dvss.n3885 dvss.n3884 9.3005
R19383 dvss.n3883 dvss.n3847 9.3005
R19384 dvss.n3882 dvss.n3881 9.3005
R19385 dvss.n3880 dvss.n3849 9.3005
R19386 dvss.n3879 dvss.n3878 9.3005
R19387 dvss.n3877 dvss.n3850 9.3005
R19388 dvss.n3876 dvss.n3875 9.3005
R19389 dvss.n3874 dvss.n3854 9.3005
R19390 dvss.n3873 dvss.n3872 9.3005
R19391 dvss.n3870 dvss.n3855 9.3005
R19392 dvss.n3869 dvss.n3857 9.3005
R19393 dvss.n3868 dvss.n3867 9.3005
R19394 dvss.n3866 dvss.n3859 9.3005
R19395 dvss.n3865 dvss.n3864 9.3005
R19396 dvss.n3609 dvss.n3608 9.3005
R19397 dvss.n3605 dvss.n3513 9.3005
R19398 dvss.n3604 dvss.n3603 9.3005
R19399 dvss.n3602 dvss.n3516 9.3005
R19400 dvss.n3601 dvss.n3600 9.3005
R19401 dvss.n3611 dvss.n3610 9.3005
R19402 dvss.n3616 dvss.n3509 9.3005
R19403 dvss.n3625 dvss.n3506 9.3005
R19404 dvss.n3628 dvss.n3505 9.3005
R19405 dvss.n3499 dvss.n3468 9.3005
R19406 dvss.n3494 dvss.n3470 9.3005
R19407 dvss.n3483 dvss.n3482 9.3005
R19408 dvss.n3992 dvss.n3456 9.3005
R19409 dvss.n3971 dvss.n3909 9.3005
R19410 dvss.n3962 dvss.n3911 9.3005
R19411 dvss.n3930 dvss.n3922 9.3005
R19412 dvss.n3929 dvss.n3928 9.3005
R19413 dvss.n3932 dvss.n3931 9.3005
R19414 dvss.n3934 dvss.n3933 9.3005
R19415 dvss.n3935 dvss.n3919 9.3005
R19416 dvss.n3937 dvss.n3936 9.3005
R19417 dvss.n3938 dvss.n3918 9.3005
R19418 dvss.n3940 dvss.n3939 9.3005
R19419 dvss.n3941 dvss.n3917 9.3005
R19420 dvss.n3943 dvss.n3942 9.3005
R19421 dvss.n3946 dvss.n3916 9.3005
R19422 dvss.n3948 dvss.n3947 9.3005
R19423 dvss.n3949 dvss.n3915 9.3005
R19424 dvss.n3951 dvss.n3950 9.3005
R19425 dvss.n3954 dvss.n3914 9.3005
R19426 dvss.n3958 dvss.n3957 9.3005
R19427 dvss.n3959 dvss.n3913 9.3005
R19428 dvss.n3961 dvss.n3960 9.3005
R19429 dvss.n3966 dvss.n3965 9.3005
R19430 dvss.n3967 dvss.n3910 9.3005
R19431 dvss.n3969 dvss.n3968 9.3005
R19432 dvss.n3974 dvss.n3973 9.3005
R19433 dvss.n3975 dvss.n3464 9.3005
R19434 dvss.n3977 dvss.n3976 9.3005
R19435 dvss.n3978 dvss.n3463 9.3005
R19436 dvss.n3982 dvss.n3981 9.3005
R19437 dvss.n3983 dvss.n3462 9.3005
R19438 dvss.n3985 dvss.n3984 9.3005
R19439 dvss.n3986 dvss.n3458 9.3005
R19440 dvss.n3988 dvss.n3987 9.3005
R19441 dvss.n3989 dvss.n3457 9.3005
R19442 dvss.n3991 dvss.n3990 9.3005
R19443 dvss.n3994 dvss.n3993 9.3005
R19444 dvss.n3995 dvss.n3455 9.3005
R19445 dvss.n3997 dvss.n3996 9.3005
R19446 dvss.n4000 dvss.n3999 9.3005
R19447 dvss.n3476 dvss.n3453 9.3005
R19448 dvss.n3485 dvss.n3474 9.3005
R19449 dvss.n3488 dvss.n3487 9.3005
R19450 dvss.n3489 dvss.n3472 9.3005
R19451 dvss.n3491 dvss.n3490 9.3005
R19452 dvss.n3493 dvss.n3492 9.3005
R19453 dvss.n3496 dvss.n3495 9.3005
R19454 dvss.n3498 dvss.n3497 9.3005
R19455 dvss.n3501 dvss.n3500 9.3005
R19456 dvss.n3503 dvss.n3502 9.3005
R19457 dvss.n3504 dvss.n3466 9.3005
R19458 dvss.n3627 dvss.n3626 9.3005
R19459 dvss.n3624 dvss.n3623 9.3005
R19460 dvss.n3617 dvss.n3507 9.3005
R19461 dvss.n3615 dvss 9.3005
R19462 dvss.n3614 dvss.n3511 9.3005
R19463 dvss.n3613 dvss.n3612 9.3005
R19464 dvss.n3597 dvss.n3596 9.3005
R19465 dvss.n3595 dvss.n3594 9.3005
R19466 dvss.n3593 dvss.n3519 9.3005
R19467 dvss.n3592 dvss.n3591 9.3005
R19468 dvss.n3590 dvss.n3520 9.3005
R19469 dvss.n3589 dvss.n3588 9.3005
R19470 dvss.n3585 dvss.n3584 9.3005
R19471 dvss.n3541 dvss.n3536 9.3005
R19472 dvss.n3543 dvss.n3542 9.3005
R19473 dvss.n3546 dvss.n3545 9.3005
R19474 dvss.n3548 dvss.n3547 9.3005
R19475 dvss.n3550 dvss.n3549 9.3005
R19476 dvss.n3552 dvss.n3551 9.3005
R19477 dvss.n3555 dvss.n3554 9.3005
R19478 dvss.n3556 dvss.n3531 9.3005
R19479 dvss.n3558 dvss.n3557 9.3005
R19480 dvss.n3559 dvss.n3530 9.3005
R19481 dvss.n3563 dvss.n3562 9.3005
R19482 dvss.n3564 dvss.n3529 9.3005
R19483 dvss.n3566 dvss.n3565 9.3005
R19484 dvss.n3568 dvss.n3567 9.3005
R19485 dvss.n3570 dvss.n3569 9.3005
R19486 dvss.n3572 dvss.n3524 9.3005
R19487 dvss.n3574 dvss.n3573 9.3005
R19488 dvss.n3575 dvss.n3523 9.3005
R19489 dvss.n3577 dvss.n3576 9.3005
R19490 dvss.n3583 dvss.n3582 9.3005
R19491 dvss.n4358 dvss.n4357 9.3005
R19492 dvss.n4359 dvss.n4324 9.3005
R19493 dvss.n4361 dvss.n4360 9.3005
R19494 dvss.n4362 dvss.n4323 9.3005
R19495 dvss.n4365 dvss.n4364 9.3005
R19496 dvss.n4366 dvss.n4322 9.3005
R19497 dvss.n4368 dvss.n4367 9.3005
R19498 dvss.n4369 dvss.n4321 9.3005
R19499 dvss.n4372 dvss.n4371 9.3005
R19500 dvss.n4356 dvss.n4355 9.3005
R19501 dvss.n4354 dvss.n4328 9.3005
R19502 dvss.n4353 dvss.n4352 9.3005
R19503 dvss.n4349 dvss.n4331 9.3005
R19504 dvss.n4344 dvss.n4335 9.3005
R19505 dvss.n4341 dvss.n4336 9.3005
R19506 dvss.n4343 dvss.n4342 9.3005
R19507 dvss.n4346 dvss.n4345 9.3005
R19508 dvss.n4348 dvss.n4347 9.3005
R19509 dvss.n4351 dvss.n4350 9.3005
R19510 dvss.n2340 dvss.n2339 9.3005
R19511 dvss.n2342 dvss.n2341 9.3005
R19512 dvss.n2344 dvss.n2343 9.3005
R19513 dvss.n2345 dvss.n2333 9.3005
R19514 dvss.n2347 dvss.n2346 9.3005
R19515 dvss.n2348 dvss.n2332 9.3005
R19516 dvss.n2350 dvss.n2349 9.3005
R19517 dvss.n2351 dvss.n2331 9.3005
R19518 dvss.n2354 dvss.n2353 9.3005
R19519 dvss.n2355 dvss.n2330 9.3005
R19520 dvss.n2357 dvss.n2356 9.3005
R19521 dvss.n2358 dvss.n2329 9.3005
R19522 dvss.n2361 dvss.n2360 9.3005
R19523 dvss.n2362 dvss.n2327 9.3005
R19524 dvss.n4487 dvss.n4486 9.3005
R19525 dvss.n4485 dvss.n4484 9.3005
R19526 dvss.n4483 dvss.n2363 9.3005
R19527 dvss.n4482 dvss.n4481 9.3005
R19528 dvss.n4480 dvss.n2364 9.3005
R19529 dvss.n4479 dvss.n4478 9.3005
R19530 dvss.n4477 dvss.n2365 9.3005
R19531 dvss.n4475 dvss.n4474 9.3005
R19532 dvss.n4473 dvss.n2368 9.3005
R19533 dvss.n4472 dvss.n4471 9.3005
R19534 dvss.n4468 dvss.n2369 9.3005
R19535 dvss.n4467 dvss.n4466 9.3005
R19536 dvss.n4465 dvss.n4464 9.3005
R19537 dvss.n4463 dvss.n2372 9.3005
R19538 dvss.n4462 dvss.n4461 9.3005
R19539 dvss.n4460 dvss.n2373 9.3005
R19540 dvss.n4459 dvss.n4458 9.3005
R19541 dvss.n4457 dvss.n2374 9.3005
R19542 dvss.n4456 dvss.n4455 9.3005
R19543 dvss.n4454 dvss.n4453 9.3005
R19544 dvss.n4452 dvss.n4451 9.3005
R19545 dvss.n4450 dvss.n2379 9.3005
R19546 dvss.n4449 dvss.n4448 9.3005
R19547 dvss.n4447 dvss.n4446 9.3005
R19548 dvss.n4445 dvss.n4444 9.3005
R19549 dvss.n4443 dvss.n2382 9.3005
R19550 dvss.n4442 dvss 9.3005
R19551 dvss.n4441 dvss.n2386 9.3005
R19552 dvss.n4440 dvss.n4439 9.3005
R19553 dvss.n4437 dvss.n2387 9.3005
R19554 dvss.n4436 dvss.n4435 9.3005
R19555 dvss.n4434 dvss.n4433 9.3005
R19556 dvss.n4432 dvss.n4431 9.3005
R19557 dvss.n4430 dvss.n2394 9.3005
R19558 dvss.n4429 dvss.n4428 9.3005
R19559 dvss.n4426 dvss.n2395 9.3005
R19560 dvss.n4425 dvss.n4424 9.3005
R19561 dvss.n4423 dvss.n2397 9.3005
R19562 dvss.n4422 dvss.n4421 9.3005
R19563 dvss.n4420 dvss.n2398 9.3005
R19564 dvss.n4418 dvss.n4417 9.3005
R19565 dvss.n4295 dvss.n2401 9.3005
R19566 dvss.n4299 dvss.n4297 9.3005
R19567 dvss.n4407 dvss.n4406 9.3005
R19568 dvss.n4405 dvss.n4298 9.3005
R19569 dvss.n4404 dvss.n4403 9.3005
R19570 dvss.n4402 dvss.n4401 9.3005
R19571 dvss.n4400 dvss.n4303 9.3005
R19572 dvss.n4399 dvss.n4305 9.3005
R19573 dvss.n4398 dvss.n4397 9.3005
R19574 dvss.n4396 dvss.n4306 9.3005
R19575 dvss.n4395 dvss.n4394 9.3005
R19576 dvss.n4391 dvss.n4307 9.3005
R19577 dvss.n4389 dvss.n4388 9.3005
R19578 dvss.n4387 dvss.n4386 9.3005
R19579 dvss.n4384 dvss.n4383 9.3005
R19580 dvss.n4382 dvss.n4317 9.3005
R19581 dvss.n4381 dvss.n4380 9.3005
R19582 dvss.n4379 dvss.n4318 9.3005
R19583 dvss.n4632 dvss.n4631 9.3005
R19584 dvss.n4629 dvss.n4624 9.3005
R19585 dvss.n4633 dvss.n4623 9.3005
R19586 dvss.n4635 dvss.n4634 9.3005
R19587 dvss.n4636 dvss.n4621 9.3005
R19588 dvss.n4640 dvss.n4639 9.3005
R19589 dvss.n4642 dvss.n4641 9.3005
R19590 dvss.n4644 dvss.n4643 9.3005
R19591 dvss.n4645 dvss.n4617 9.3005
R19592 dvss.n4647 dvss.n4646 9.3005
R19593 dvss.n4648 dvss.n4615 9.3005
R19594 dvss.n4650 dvss.n4649 9.3005
R19595 dvss.n4651 dvss.n4614 9.3005
R19596 dvss.n4653 dvss.n4652 9.3005
R19597 dvss.n4655 dvss.n4613 9.3005
R19598 dvss.n4658 dvss.n4657 9.3005
R19599 dvss.n4504 dvss.n4499 9.3005
R19600 dvss.n4506 dvss.n4505 9.3005
R19601 dvss.n4509 dvss.n4508 9.3005
R19602 dvss.n4511 dvss.n4510 9.3005
R19603 dvss.n4512 dvss.n4497 9.3005
R19604 dvss.n4514 dvss.n4513 9.3005
R19605 dvss.n4518 dvss.n4494 9.3005
R19606 dvss.n4522 dvss.n4521 9.3005
R19607 dvss.n4523 dvss.n4492 9.3005
R19608 dvss.n4788 dvss.n4787 9.3005
R19609 dvss.n4786 dvss.n4493 9.3005
R19610 dvss.n4785 dvss.n4784 9.3005
R19611 dvss.n4781 dvss.n4524 9.3005
R19612 dvss.n4780 dvss.n4779 9.3005
R19613 dvss.n4778 dvss.n4777 9.3005
R19614 dvss.n4776 dvss.n4527 9.3005
R19615 dvss.n4775 dvss.n4774 9.3005
R19616 dvss.n4773 dvss.n4772 9.3005
R19617 dvss.n4771 dvss.n4770 9.3005
R19618 dvss.n4769 dvss.n4768 9.3005
R19619 dvss.n4767 dvss.n4531 9.3005
R19620 dvss.n4765 dvss.n4764 9.3005
R19621 dvss.n4763 dvss.n4532 9.3005
R19622 dvss.n4762 dvss.n4761 9.3005
R19623 dvss.n4759 dvss.n4533 9.3005
R19624 dvss.n4758 dvss.n4757 9.3005
R19625 dvss.n4756 dvss.n4755 9.3005
R19626 dvss.n4754 dvss.n4535 9.3005
R19627 dvss.n4753 dvss.n4752 9.3005
R19628 dvss.n4751 dvss.n4750 9.3005
R19629 dvss.n4748 dvss.n4747 9.3005
R19630 dvss.n4746 dvss.n4538 9.3005
R19631 dvss.n4745 dvss.n4744 9.3005
R19632 dvss.n4742 dvss.n4539 9.3005
R19633 dvss.n4741 dvss.n4740 9.3005
R19634 dvss.n4739 dvss.n4540 9.3005
R19635 dvss.n4738 dvss.n4737 9.3005
R19636 dvss.n4736 dvss.n4544 9.3005
R19637 dvss.n4735 dvss.n4734 9.3005
R19638 dvss.n4733 dvss.n4732 9.3005
R19639 dvss.n4731 dvss.n4548 9.3005
R19640 dvss.n4730 dvss.n4729 9.3005
R19641 dvss.n4728 dvss.n4552 9.3005
R19642 dvss.n4727 dvss.n4726 9.3005
R19643 dvss.n4724 dvss.n4553 9.3005
R19644 dvss.n4722 dvss.n4721 9.3005
R19645 dvss.n4720 dvss.n4719 9.3005
R19646 dvss.n4716 dvss.n4555 9.3005
R19647 dvss.n4715 dvss.n4714 9.3005
R19648 dvss.n4713 dvss.n4558 9.3005
R19649 dvss.n4568 dvss.n4559 9.3005
R19650 dvss.n4574 dvss.n4573 9.3005
R19651 dvss.n4577 dvss.n4564 9.3005
R19652 dvss.n4704 dvss.n4703 9.3005
R19653 dvss.n4701 dvss.n4700 9.3005
R19654 dvss.n4699 dvss.n4698 9.3005
R19655 dvss.n4695 dvss.n4581 9.3005
R19656 dvss.n4694 dvss.n4693 9.3005
R19657 dvss.n4692 dvss.n4691 9.3005
R19658 dvss.n4690 dvss.n4584 9.3005
R19659 dvss.n4689 dvss.n4688 9.3005
R19660 dvss.n4687 dvss.n4686 9.3005
R19661 dvss.n4590 dvss.n4589 9.3005
R19662 dvss.n4681 dvss.n4680 9.3005
R19663 dvss.n4679 dvss.n4678 9.3005
R19664 dvss.n4677 dvss.n4594 9.3005
R19665 dvss.n4676 dvss.n4675 9.3005
R19666 dvss.n4674 dvss.n4600 9.3005
R19667 dvss.n4673 dvss.n4672 9.3005
R19668 dvss.n4671 dvss.n4601 9.3005
R19669 dvss.n4669 dvss.n4668 9.3005
R19670 dvss.n4667 dvss.n4606 9.3005
R19671 dvss.n4666 dvss.n4665 9.3005
R19672 dvss.n4612 dvss.n4608 9.3005
R19673 dvss.n4660 dvss.n4659 9.3005
R19674 dvss.n5029 dvss.n5028 9.3005
R19675 dvss.n5031 dvss.n5030 9.3005
R19676 dvss.n5034 dvss.n5020 9.3005
R19677 dvss.n5036 dvss.n5035 9.3005
R19678 dvss.n5037 dvss.n5019 9.3005
R19679 dvss.n5039 dvss.n5038 9.3005
R19680 dvss.n5040 dvss.n5016 9.3005
R19681 dvss.n5042 dvss.n5041 9.3005
R19682 dvss.n5043 dvss.n5015 9.3005
R19683 dvss.n5045 dvss.n5044 9.3005
R19684 dvss.n5046 dvss.n5014 9.3005
R19685 dvss.n5050 dvss.n5049 9.3005
R19686 dvss.n5051 dvss.n5013 9.3005
R19687 dvss.n5053 dvss.n5052 9.3005
R19688 dvss.n5056 dvss.n5012 9.3005
R19689 dvss.n5058 dvss.n5057 9.3005
R19690 dvss.n5059 dvss.n5011 9.3005
R19691 dvss.n5061 dvss.n5060 9.3005
R19692 dvss.n5062 dvss.n5008 9.3005
R19693 dvss.n5064 dvss.n5063 9.3005
R19694 dvss.n5065 dvss.n5007 9.3005
R19695 dvss.n5067 dvss.n5066 9.3005
R19696 dvss.n5069 dvss.n5005 9.3005
R19697 dvss.n5071 dvss.n5070 9.3005
R19698 dvss.n5072 dvss.n5004 9.3005
R19699 dvss.n5074 dvss.n5073 9.3005
R19700 dvss.n5075 dvss.n1226 9.3005
R19701 dvss.n5077 dvss.n5076 9.3005
R19702 dvss.n5078 dvss.n1225 9.3005
R19703 dvss.n5080 dvss.n5079 9.3005
R19704 dvss.n5081 dvss.n1224 9.3005
R19705 dvss.n5083 dvss.n5082 9.3005
R19706 dvss.n5084 dvss.n1223 9.3005
R19707 dvss.n5086 dvss.n5085 9.3005
R19708 dvss.n5087 dvss.n1221 9.3005
R19709 dvss.n5089 dvss.n5088 9.3005
R19710 dvss.n5091 dvss.n5090 9.3005
R19711 dvss.n5093 dvss.n5092 9.3005
R19712 dvss.n1218 dvss.n1216 9.3005
R19713 dvss.n4931 dvss.n4930 9.3005
R19714 dvss.n4932 dvss.n4919 9.3005
R19715 dvss.n4934 dvss.n4933 9.3005
R19716 dvss.n4935 dvss.n4918 9.3005
R19717 dvss.n4937 dvss.n4936 9.3005
R19718 dvss.n4938 dvss.n4917 9.3005
R19719 dvss.n4942 dvss.n4941 9.3005
R19720 dvss.n4944 dvss.n4943 9.3005
R19721 dvss.n4946 dvss.n4945 9.3005
R19722 dvss.n4947 dvss.n4915 9.3005
R19723 dvss.n4949 dvss.n4948 9.3005
R19724 dvss.n4950 dvss.n4913 9.3005
R19725 dvss.n4952 dvss.n4951 9.3005
R19726 dvss.n4953 dvss.n1228 9.3005
R19727 dvss.n4954 dvss.n4912 9.3005
R19728 dvss.n4956 dvss.n4955 9.3005
R19729 dvss.n4958 dvss.n4957 9.3005
R19730 dvss.n4959 dvss.n4911 9.3005
R19731 dvss.n4961 dvss.n4960 9.3005
R19732 dvss.n4962 dvss.n4909 9.3005
R19733 dvss.n4963 dvss.n4908 9.3005
R19734 dvss.n4967 dvss.n4966 9.3005
R19735 dvss.n4969 dvss.n4968 9.3005
R19736 dvss.n4971 dvss.n4970 9.3005
R19737 dvss.n4972 dvss.n4906 9.3005
R19738 dvss.n4974 dvss.n4973 9.3005
R19739 dvss.n4975 dvss.n4904 9.3005
R19740 dvss.n4976 dvss.n4903 9.3005
R19741 dvss.n4980 dvss.n4979 9.3005
R19742 dvss.n4982 dvss.n4981 9.3005
R19743 dvss.n4984 dvss.n4983 9.3005
R19744 dvss.n4985 dvss.n4901 9.3005
R19745 dvss.n4987 dvss.n4986 9.3005
R19746 dvss.n4988 dvss.n4899 9.3005
R19747 dvss.n4989 dvss.n4898 9.3005
R19748 dvss.n4993 dvss.n4992 9.3005
R19749 dvss.n4995 dvss.n4994 9.3005
R19750 dvss.n4997 dvss.n4996 9.3005
R19751 dvss.n4998 dvss.n4896 9.3005
R19752 dvss.n5000 dvss.n4999 9.3005
R19753 dvss.n5001 dvss.n4894 9.3005
R19754 dvss.n5002 dvss.n4893 9.3005
R19755 dvss.n4892 dvss.n4857 9.3005
R19756 dvss.n4891 dvss.n4890 9.3005
R19757 dvss.n4888 dvss.n4858 9.3005
R19758 dvss.n4887 dvss.n4886 9.3005
R19759 dvss.n4885 dvss.n4884 9.3005
R19760 dvss.n4883 dvss.n4860 9.3005
R19761 dvss.n4882 dvss.n4881 9.3005
R19762 dvss.n4880 dvss.n4861 9.3005
R19763 dvss.n4879 dvss.n4878 9.3005
R19764 dvss.n4877 dvss.n4862 9.3005
R19765 dvss.n4876 dvss.n4875 9.3005
R19766 dvss.n4874 dvss.n4873 9.3005
R19767 dvss.n4869 dvss.n4868 9.3005
R19768 dvss.n4870 dvss.n4864 9.3005
R19769 dvss.n4872 dvss.n4871 9.3005
R19770 dvss.n4064 dvss.n4063 9.3005
R19771 dvss.n4066 dvss.n4065 9.3005
R19772 dvss.n4067 dvss.n4058 9.3005
R19773 dvss.n4069 dvss.n4068 9.3005
R19774 dvss.n4071 dvss.n4055 9.3005
R19775 dvss.n4074 dvss.n4073 9.3005
R19776 dvss.n4076 dvss.n4075 9.3005
R19777 dvss.n4078 dvss.n4077 9.3005
R19778 dvss.n4080 dvss.n4079 9.3005
R19779 dvss.n4082 dvss.n4052 9.3005
R19780 dvss.n4086 dvss.n4085 9.3005
R19781 dvss.n4088 dvss.n4051 9.3005
R19782 dvss.n4090 dvss.n4089 9.3005
R19783 dvss.n4091 dvss.n4047 9.3005
R19784 dvss.n4092 dvss.n4045 9.3005
R19785 dvss.n4094 dvss.n4093 9.3005
R19786 dvss.n4095 dvss.n4044 9.3005
R19787 dvss.n4097 dvss.n4096 9.3005
R19788 dvss.n4098 dvss.n4042 9.3005
R19789 dvss.n4102 dvss.n4101 9.3005
R19790 dvss.n4103 dvss.n4041 9.3005
R19791 dvss.n4105 dvss.n4104 9.3005
R19792 dvss.n4106 dvss.n4040 9.3005
R19793 dvss.n4107 dvss.n4038 9.3005
R19794 dvss.n4109 dvss.n4108 9.3005
R19795 dvss.n4111 dvss.n4110 9.3005
R19796 dvss.n4116 dvss.n4035 9.3005
R19797 dvss.n4118 dvss.n4117 9.3005
R19798 dvss.n4119 dvss.n4034 9.3005
R19799 dvss.n4121 dvss.n4120 9.3005
R19800 dvss.n4122 dvss.n4033 9.3005
R19801 dvss.n4123 dvss.n4032 9.3005
R19802 dvss.n4124 dvss.n4030 9.3005
R19803 dvss.n4126 dvss.n4125 9.3005
R19804 dvss.n4127 dvss.n4029 9.3005
R19805 dvss.n4129 dvss.n4128 9.3005
R19806 dvss.n4132 dvss.n4027 9.3005
R19807 dvss.n4136 dvss.n4135 9.3005
R19808 dvss.n4137 dvss.n4025 9.3005
R19809 dvss.n4189 dvss.n4026 9.3005
R19810 dvss.n4188 dvss.n4187 9.3005
R19811 dvss.n4186 dvss.n4138 9.3005
R19812 dvss.n4183 dvss.n4182 9.3005
R19813 dvss.n4181 dvss.n4142 9.3005
R19814 dvss.n4180 dvss.n4179 9.3005
R19815 dvss.n4178 dvss.n4143 9.3005
R19816 dvss.n4177 dvss.n4145 9.3005
R19817 dvss.n4176 dvss.n4146 9.3005
R19818 dvss.n4175 dvss.n4149 9.3005
R19819 dvss.n4173 dvss.n4172 9.3005
R19820 dvss.n4171 dvss.n4151 9.3005
R19821 dvss.n4159 dvss.n4152 9.3005
R19822 dvss.n4163 dvss.n4162 9.3005
R19823 dvss.n4013 dvss.n4011 9.3005
R19824 dvss.n4288 dvss.n4287 9.3005
R19825 dvss.n4286 dvss.n4012 9.3005
R19826 dvss.n4284 dvss.n4283 9.3005
R19827 dvss.n4282 dvss.n4281 9.3005
R19828 dvss.n4280 dvss.n4018 9.3005
R19829 dvss.n4279 dvss.n4278 9.3005
R19830 dvss.n4277 dvss.n4021 9.3005
R19831 dvss.n4276 dvss.n4275 9.3005
R19832 dvss.n4272 dvss.n4022 9.3005
R19833 dvss.n4271 dvss.n4270 9.3005
R19834 dvss.n4269 dvss.n4024 9.3005
R19835 dvss.n4268 dvss.n4267 9.3005
R19836 dvss.n4266 dvss.n4194 9.3005
R19837 dvss.n4265 dvss.n4264 9.3005
R19838 dvss.n4263 dvss.n4262 9.3005
R19839 dvss.n4260 dvss.n4197 9.3005
R19840 dvss.n4259 dvss.n4258 9.3005
R19841 dvss.n4257 dvss.n4199 9.3005
R19842 dvss.n4256 dvss.n4255 9.3005
R19843 dvss.n4252 dvss.n4251 9.3005
R19844 dvss.n4250 dvss.n4202 9.3005
R19845 dvss.n4249 dvss.n4248 9.3005
R19846 dvss.n4247 dvss.n4203 9.3005
R19847 dvss.n4246 dvss.n4245 9.3005
R19848 dvss.n4244 dvss.n4204 9.3005
R19849 dvss.n4243 dvss.n4242 9.3005
R19850 dvss.n4241 dvss.n4205 9.3005
R19851 dvss.n4240 dvss.n4239 9.3005
R19852 dvss.n4238 dvss.n4237 9.3005
R19853 dvss.n4236 dvss.n4210 9.3005
R19854 dvss.n4235 dvss.n4234 9.3005
R19855 dvss.n4233 dvss.n4211 9.3005
R19856 dvss.n4232 dvss.n4231 9.3005
R19857 dvss.n4228 dvss.n4212 9.3005
R19858 dvss.n4227 dvss.n4215 9.3005
R19859 dvss.n4226 dvss.n4225 9.3005
R19860 dvss.n4224 dvss.n4217 9.3005
R19861 dvss.n4223 dvss.n4222 9.3005
R19862 dvss.n4191 dvss.n4190 9.3005
R19863 dvss.n4819 dvss.n4818 9.3005
R19864 dvss.n4850 dvss.n4849 9.3005
R19865 dvss.n2324 dvss.n2323 9.3005
R19866 dvss.n3331 dvss.n3330 9.3005
R19867 dvss.n3332 dvss.n3331 9.3005
R19868 dvss.n3282 dvss.n3281 9.3005
R19869 dvss.n3281 dvss.n3280 9.3005
R19870 dvss.n3278 dvss.n3275 9.3005
R19871 dvss.n3278 dvss.n3277 9.3005
R19872 dvss.n3274 dvss.n3271 9.3005
R19873 dvss.n3274 dvss.n3273 9.3005
R19874 dvss.n3333 dvss.n3128 9.3005
R19875 dvss.n3132 dvss.n3131 9.3005
R19876 dvss.n3329 dvss.n3328 9.3005
R19877 dvss.n3139 dvss.n3133 9.3005
R19878 dvss.n3322 dvss.n3140 9.3005
R19879 dvss.n3321 dvss.n3141 9.3005
R19880 dvss.n3320 dvss.n3142 9.3005
R19881 dvss.n3147 dvss.n3143 9.3005
R19882 dvss.n3314 dvss.n3148 9.3005
R19883 dvss.n3313 dvss.n3149 9.3005
R19884 dvss.n3312 dvss.n3150 9.3005
R19885 dvss.n3270 dvss.n3151 9.3005
R19886 dvss.n3306 dvss.n3155 9.3005
R19887 dvss.n3305 dvss.n3156 9.3005
R19888 dvss.n3304 dvss.n3157 9.3005
R19889 dvss.n3268 dvss.n3158 9.3005
R19890 dvss.n3297 dvss.n3269 9.3005
R19891 dvss.n3296 dvss.n3283 9.3005
R19892 dvss.n3295 dvss.n3284 9.3005
R19893 dvss.n3287 dvss.n3285 9.3005
R19894 dvss.n3289 dvss.n3288 9.3005
R19895 dvss.n3248 dvss.n3247 9.3005
R19896 dvss.n3173 dvss.n3172 9.3005
R19897 dvss.n3231 dvss.n3178 9.3005
R19898 dvss.n3214 dvss.n3213 9.3005
R19899 dvss.n3217 dvss.n3216 9.3005
R19900 dvss.n3229 dvss.n3228 9.3005
R19901 dvss.n3232 dvss.n3231 9.3005
R19902 dvss.n324 dvss.n323 9.3005
R19903 dvss.n322 dvss.n321 9.3005
R19904 dvss.n320 dvss.n319 9.3005
R19905 dvss.n318 dvss.n312 9.3005
R19906 dvss.n317 dvss.n316 9.3005
R19907 dvss.n291 dvss.n290 9.3005
R19908 dvss.n293 dvss.n285 9.3005
R19909 dvss.n297 dvss.n296 9.3005
R19910 dvss.n298 dvss.n284 9.3005
R19911 dvss.n300 dvss.n299 9.3005
R19912 dvss.n302 dvss.n282 9.3005
R19913 dvss.n306 dvss.n305 9.3005
R19914 dvss.n307 dvss.n279 9.3005
R19915 dvss.n332 dvss.n331 9.3005
R19916 dvss.n330 dvss.n329 9.3005
R19917 dvss.n327 dvss.n308 9.3005
R19918 dvss.n326 dvss.n325 9.3005
R19919 dvss.n454 dvss.n381 9.3005
R19920 dvss.n453 dvss.n452 9.3005
R19921 dvss.n451 dvss.n383 9.3005
R19922 dvss.n450 dvss.n449 9.3005
R19923 dvss.n447 dvss.n446 9.3005
R19924 dvss.n401 dvss.n400 9.3005
R19925 dvss.n402 dvss.n394 9.3005
R19926 dvss.n404 dvss.n403 9.3005
R19927 dvss.n406 dvss.n392 9.3005
R19928 dvss.n410 dvss.n409 9.3005
R19929 dvss.n411 dvss.n391 9.3005
R19930 dvss.n413 dvss.n412 9.3005
R19931 dvss.n415 dvss.n389 9.3005
R19932 dvss.n439 dvss.n438 9.3005
R19933 dvss.n441 dvss.n440 9.3005
R19934 dvss.n443 dvss.n385 9.3005
R19935 dvss.n445 dvss.n444 9.3005
R19936 dvss.n6622 dvss.n6621 9.3005
R19937 dvss.n6625 dvss.n6624 9.3005
R19938 dvss.n6626 dvss.n245 9.3005
R19939 dvss.n6628 dvss.n6627 9.3005
R19940 dvss.n6629 dvss.n243 9.3005
R19941 dvss.n263 dvss.n262 9.3005
R19942 dvss.n264 dvss.n256 9.3005
R19943 dvss.n266 dvss.n265 9.3005
R19944 dvss.n268 dvss.n254 9.3005
R19945 dvss.n272 dvss.n271 9.3005
R19946 dvss.n273 dvss.n253 9.3005
R19947 dvss.n275 dvss.n274 9.3005
R19948 dvss.n277 dvss.n251 9.3005
R19949 dvss.n6614 dvss.n6613 9.3005
R19950 dvss.n6616 dvss.n6615 9.3005
R19951 dvss.n6618 dvss.n247 9.3005
R19952 dvss.n6620 dvss.n6619 9.3005
R19953 dvss.n6599 dvss.n6598 9.3005
R19954 dvss.n6597 dvss.n6596 9.3005
R19955 dvss.n6595 dvss.n6594 9.3005
R19956 dvss.n6593 dvss.n373 9.3005
R19957 dvss.n6592 dvss.n6591 9.3005
R19958 dvss.n6590 dvss.n6589 9.3005
R19959 dvss.n6588 dvss.n6587 9.3005
R19960 dvss.n6586 dvss.n6585 9.3005
R19961 dvss.n6584 dvss.n377 9.3005
R19962 dvss.n6583 dvss.n6582 9.3005
R19963 dvss.n351 dvss.n350 9.3005
R19964 dvss.n352 dvss.n344 9.3005
R19965 dvss.n354 dvss.n353 9.3005
R19966 dvss.n356 dvss.n342 9.3005
R19967 dvss.n360 dvss.n359 9.3005
R19968 dvss.n361 dvss.n341 9.3005
R19969 dvss.n363 dvss.n362 9.3005
R19970 dvss.n365 dvss.n339 9.3005
R19971 dvss.n369 dvss.n368 9.3005
R19972 dvss.n370 dvss.n336 9.3005
R19973 dvss.n6602 dvss.n6601 9.3005
R19974 dvss.n6600 dvss.n338 9.3005
R19975 dvss.n1735 dvss.n1612 9.3005
R19976 dvss.n1613 dvss.n1612 9.3005
R19977 dvss.n1763 dvss.n1564 9.3005
R19978 dvss.n1764 dvss.n1763 9.3005
R19979 dvss.n1782 dvss.n1781 9.3005
R19980 dvss.n1781 dvss.n1778 9.3005
R19981 dvss.n1864 dvss.n1509 9.3005
R19982 dvss.n1865 dvss.n1864 9.3005
R19983 dvss.n1862 dvss.n1514 9.3005
R19984 dvss.n1862 dvss.n1861 9.3005
R19985 dvss.n1830 dvss.n1513 9.3005
R19986 dvss.n1533 dvss.n1513 9.3005
R19987 dvss.n1897 dvss.n1896 9.3005
R19988 dvss.n1896 dvss.n1893 9.3005
R19989 dvss.n2024 dvss.n2023 9.3005
R19990 dvss.n2023 dvss.n2022 9.3005
R19991 dvss.n1972 dvss.n1971 9.3005
R19992 dvss.n1971 dvss.n1970 9.3005
R19993 dvss.n1944 dvss.n1943 9.3005
R19994 dvss.n1943 dvss.n1942 9.3005
R19995 dvss.n2038 dvss.n1435 9.3005
R19996 dvss.n2039 dvss.n2038 9.3005
R19997 dvss.n1407 dvss.n895 9.3005
R19998 dvss.n1407 dvss.n1406 9.3005
R19999 dvss.n1372 dvss.n1360 9.3005
R20000 dvss.n1369 dvss.n1360 9.3005
R20001 dvss.n2097 dvss.n2096 9.3005
R20002 dvss.n2096 dvss.n2095 9.3005
R20003 dvss.n5716 dvss.n5715 9.3005
R20004 dvss.n5717 dvss.n5716 9.3005
R20005 dvss.n5680 dvss.n5679 9.3005
R20006 dvss.n5680 dvss.n943 9.3005
R20007 dvss.n5685 dvss.n5684 9.3005
R20008 dvss.n5684 dvss.n5683 9.3005
R20009 dvss.n942 dvss.n940 9.3005
R20010 dvss.n942 dvss.n928 9.3005
R20011 dvss.n962 dvss.n961 9.3005
R20012 dvss.n961 dvss.n958 9.3005
R20013 dvss.n6127 dvss.n6126 9.3005
R20014 dvss.n6126 dvss.n6125 9.3005
R20015 dvss.n5632 dvss.n5631 9.3005
R20016 dvss.n5631 dvss.n5630 9.3005
R20017 dvss.n5643 dvss.n5641 9.3005
R20018 dvss.n5644 dvss.n5643 9.3005
R20019 dvss.n6141 dvss.n785 9.3005
R20020 dvss.n6142 dvss.n6141 9.3005
R20021 dvss.n757 dvss.n756 9.3005
R20022 dvss.n757 dvss.n538 9.3005
R20023 dvss.n623 dvss.n537 9.3005
R20024 dvss.n621 dvss.n537 9.3005
R20025 dvss.n6200 dvss.n6199 9.3005
R20026 dvss.n6199 dvss.n6198 9.3005
R20027 dvss.n744 dvss.n743 9.3005
R20028 dvss.n745 dvss.n744 9.3005
R20029 dvss.n708 dvss.n129 9.3005
R20030 dvss.n708 dvss.n707 9.3005
R20031 dvss.n713 dvss.n712 9.3005
R20032 dvss.n712 dvss.n711 9.3005
R20033 dvss.n588 dvss.n586 9.3005
R20034 dvss.n588 dvss.n574 9.3005
R20035 dvss.n6700 dvss.n6699 9.3005
R20036 dvss.n6701 dvss.n6700 9.3005
R20037 dvss.n6868 dvss.n6867 9.3005
R20038 dvss.n6867 dvss.n6866 9.3005
R20039 dvss.n6669 dvss.n6668 9.3005
R20040 dvss.n6668 dvss.n6667 9.3005
R20041 dvss.n170 dvss.n169 9.3005
R20042 dvss.n169 dvss.n162 9.3005
R20043 dvss.n6882 dvss.n61 9.3005
R20044 dvss.n6883 dvss.n6882 9.3005
R20045 dvss.n6486 dvss.n6485 9.3005
R20046 dvss.n6485 dvss.n6484 9.3005
R20047 dvss.n6452 dvss.n6451 9.3005
R20048 dvss.n6451 dvss.n6448 9.3005
R20049 dvss.n6941 dvss.n6940 9.3005
R20050 dvss.n6940 dvss.n6939 9.3005
R20051 dvss.n1711 dvss.n1710 9.3005
R20052 dvss.n1710 dvss.n1709 9.3005
R20053 dvss.n1767 dvss.n1766 9.3005
R20054 dvss.n1766 dvss.n1765 9.3005
R20055 dvss.n1842 dvss.n1517 9.3005
R20056 dvss.n1840 dvss.n1839 9.3005
R20057 dvss.n1828 dvss.n1827 9.3005
R20058 dvss.n1786 dvss.n1785 9.3005
R20059 dvss.n1805 dvss.n1804 9.3005
R20060 dvss.n1810 dvss.n1809 9.3005
R20061 dvss.n1829 dvss.n1828 9.3005
R20062 dvss.n1974 dvss.n1973 9.3005
R20063 dvss.n1968 dvss.n1946 9.3005
R20064 dvss.n1940 dvss.n1939 9.3005
R20065 dvss.n1910 dvss.n1909 9.3005
R20066 dvss.n1920 dvss.n1919 9.3005
R20067 dvss.n1925 dvss.n1924 9.3005
R20068 dvss.n1941 dvss.n1940 9.3005
R20069 dvss.n1388 dvss.n1387 9.3005
R20070 dvss.n1375 dvss.n1374 9.3005
R20071 dvss.n2093 dvss.n1355 9.3005
R20072 dvss.n2075 dvss.n2074 9.3005
R20073 dvss.n2078 dvss.n2077 9.3005
R20074 dvss.n2091 dvss.n2090 9.3005
R20075 dvss.n2094 dvss.n2093 9.3005
R20076 dvss.n5687 dvss.n5686 9.3005
R20077 dvss.n939 dvss.n936 9.3005
R20078 dvss.n5700 dvss.n5699 9.3005
R20079 dvss.n5710 dvss.n5709 9.3005
R20080 dvss.n5707 dvss.n5706 9.3005
R20081 dvss.n5697 dvss.n5696 9.3005
R20082 dvss.n5699 dvss.n5695 9.3005
R20083 dvss.n5634 dvss.n5633 9.3005
R20084 dvss.n5628 dvss.n1106 9.3005
R20085 dvss.n1099 dvss.n1081 9.3005
R20086 dvss.n1086 dvss.n1085 9.3005
R20087 dvss.n1093 dvss.n1092 9.3005
R20088 dvss.n1097 dvss.n1096 9.3005
R20089 dvss.n1100 dvss.n1099 9.3005
R20090 dvss.n640 dvss.n639 9.3005
R20091 dvss.n625 dvss.n624 9.3005
R20092 dvss.n6196 dvss.n532 9.3005
R20093 dvss.n6178 dvss.n6177 9.3005
R20094 dvss.n6181 dvss.n6180 9.3005
R20095 dvss.n6194 dvss.n6193 9.3005
R20096 dvss.n6197 dvss.n6196 9.3005
R20097 dvss.n715 dvss.n714 9.3005
R20098 dvss.n585 dvss.n582 9.3005
R20099 dvss.n728 dvss.n727 9.3005
R20100 dvss.n738 dvss.n737 9.3005
R20101 dvss.n735 dvss.n734 9.3005
R20102 dvss.n725 dvss.n724 9.3005
R20103 dvss.n727 dvss.n723 9.3005
R20104 dvss.n6671 dvss.n6670 9.3005
R20105 dvss.n6665 dvss.n173 9.3005
R20106 dvss.n6684 dvss.n6683 9.3005
R20107 dvss.n6694 dvss.n6693 9.3005
R20108 dvss.n6691 dvss.n6690 9.3005
R20109 dvss.n6681 dvss.n6680 9.3005
R20110 dvss.n6683 dvss.n6679 9.3005
R20111 dvss.n6467 dvss.n6466 9.3005
R20112 dvss.n6454 dvss.n6453 9.3005
R20113 dvss.n6937 dvss.n30 9.3005
R20114 dvss.n6919 dvss.n6918 9.3005
R20115 dvss.n6922 dvss.n6921 9.3005
R20116 dvss.n6935 dvss.n6934 9.3005
R20117 dvss.n6938 dvss.n6937 9.3005
R20118 dvss.n1616 dvss.n1608 9.3005
R20119 dvss.n1617 dvss.n1616 9.3005
R20120 dvss.n5117 dvss.n5116 9.3005
R20121 dvss.n5116 dvss.n5112 9.3005
R20122 dvss.n5127 dvss.n5126 9.3005
R20123 dvss.n5126 dvss.n5122 9.3005
R20124 dvss.n5137 dvss.n5136 9.3005
R20125 dvss.n5136 dvss.n5133 9.3005
R20126 dvss.n5164 dvss.n5163 9.3005
R20127 dvss.n5163 dvss.n5162 9.3005
R20128 dvss.n5160 dvss.n5157 9.3005
R20129 dvss.n5160 dvss.n5159 9.3005
R20130 dvss.n5156 dvss.n5153 9.3005
R20131 dvss.n5156 dvss.n5155 9.3005
R20132 dvss.n5176 dvss.n5175 9.3005
R20133 dvss.n5175 dvss.n5172 9.3005
R20134 dvss.n5203 dvss.n5202 9.3005
R20135 dvss.n5202 dvss.n5201 9.3005
R20136 dvss.n5199 dvss.n5196 9.3005
R20137 dvss.n5199 dvss.n5198 9.3005
R20138 dvss.n5195 dvss.n5192 9.3005
R20139 dvss.n5195 dvss.n5194 9.3005
R20140 dvss.n5215 dvss.n5214 9.3005
R20141 dvss.n5214 dvss.n5211 9.3005
R20142 dvss.n5242 dvss.n5241 9.3005
R20143 dvss.n5241 dvss.n5240 9.3005
R20144 dvss.n5238 dvss.n5235 9.3005
R20145 dvss.n5238 dvss.n5237 9.3005
R20146 dvss.n5234 dvss.n5231 9.3005
R20147 dvss.n5234 dvss.n5233 9.3005
R20148 dvss.n5254 dvss.n5253 9.3005
R20149 dvss.n5253 dvss.n5250 9.3005
R20150 dvss.n5281 dvss.n5280 9.3005
R20151 dvss.n5280 dvss.n5279 9.3005
R20152 dvss.n5277 dvss.n5274 9.3005
R20153 dvss.n5277 dvss.n5276 9.3005
R20154 dvss.n5273 dvss.n5270 9.3005
R20155 dvss.n5273 dvss.n5272 9.3005
R20156 dvss.n5504 dvss.n5503 9.3005
R20157 dvss.n5503 dvss.n5500 9.3005
R20158 dvss.n5538 dvss.n5537 9.3005
R20159 dvss.n5537 dvss.n5536 9.3005
R20160 dvss.n5534 dvss.n5531 9.3005
R20161 dvss.n5534 dvss.n5533 9.3005
R20162 dvss.n5529 dvss.n1136 9.3005
R20163 dvss.n5529 dvss.n5528 9.3005
R20164 dvss.n5558 dvss.n5557 9.3005
R20165 dvss.n5557 dvss.n5554 9.3005
R20166 dvss.n6233 dvss.n6232 9.3005
R20167 dvss.n6234 dvss.n6233 9.3005
R20168 dvss.n6229 dvss.n512 9.3005
R20169 dvss.n6229 dvss.n6228 9.3005
R20170 dvss.n6215 dvss.n511 9.3005
R20171 dvss.n6213 dvss.n511 9.3005
R20172 dvss.n6261 dvss.n6260 9.3005
R20173 dvss.n6260 dvss.n6257 9.3005
R20174 dvss.n6301 dvss.n474 9.3005
R20175 dvss.n6302 dvss.n6301 9.3005
R20176 dvss.n6299 dvss.n483 9.3005
R20177 dvss.n6299 dvss.n6298 9.3005
R20178 dvss.n6287 dvss.n482 9.3005
R20179 dvss.n6285 dvss.n482 9.3005
R20180 dvss.n6328 dvss.n6327 9.3005
R20181 dvss.n6329 dvss.n6328 9.3005
R20182 dvss.n6557 dvss.n6556 9.3005
R20183 dvss.n6557 dvss.n6349 9.3005
R20184 dvss.n6352 dvss.n6348 9.3005
R20185 dvss.n6348 dvss.n6347 9.3005
R20186 dvss.n6562 dvss.n6560 9.3005
R20187 dvss.n6563 dvss.n6562 9.3005
R20188 dvss.n6378 dvss.n6377 9.3005
R20189 dvss.n6377 dvss.n6374 9.3005
R20190 dvss.n6424 dvss.n6423 9.3005
R20191 dvss.n6423 dvss.n6422 9.3005
R20192 dvss.n6420 dvss.n6415 9.3005
R20193 dvss.n6420 dvss.n6419 9.3005
R20194 dvss.n6414 dvss.n6411 9.3005
R20195 dvss.n6414 dvss.n6413 9.3005
R20196 dvss.n5492 dvss.n1208 9.3005
R20197 dvss.n5491 dvss.n5103 9.3005
R20198 dvss.n5490 dvss.n5104 9.3005
R20199 dvss.n5488 dvss.n5105 9.3005
R20200 dvss.n5485 dvss.n5106 9.3005
R20201 dvss.n5484 dvss.n5107 9.3005
R20202 dvss.n5481 dvss.n5108 9.3005
R20203 dvss.n5480 dvss.n5109 9.3005
R20204 dvss.n5477 dvss.n5110 9.3005
R20205 dvss.n5476 dvss.n5111 9.3005
R20206 dvss.n5473 dvss.n5118 9.3005
R20207 dvss.n5472 dvss.n5119 9.3005
R20208 dvss.n5469 dvss.n5120 9.3005
R20209 dvss.n5468 dvss.n5121 9.3005
R20210 dvss.n5465 dvss.n5128 9.3005
R20211 dvss.n5464 dvss.n5129 9.3005
R20212 dvss.n5461 dvss.n5130 9.3005
R20213 dvss.n5460 dvss.n5131 9.3005
R20214 dvss.n5457 dvss.n5132 9.3005
R20215 dvss.n5456 dvss.n5138 9.3005
R20216 dvss.n5453 dvss.n5139 9.3005
R20217 dvss.n5452 dvss.n5140 9.3005
R20218 dvss.n5449 dvss.n5141 9.3005
R20219 dvss.n5448 dvss.n5142 9.3005
R20220 dvss.n5445 dvss.n5143 9.3005
R20221 dvss.n5444 dvss.n5144 9.3005
R20222 dvss.n5441 dvss.n5145 9.3005
R20223 dvss.n5440 dvss.n5146 9.3005
R20224 dvss.n5437 dvss.n5147 9.3005
R20225 dvss.n5436 dvss.n5148 9.3005
R20226 dvss.n5433 dvss.n5149 9.3005
R20227 dvss.n5432 dvss.n5150 9.3005
R20228 dvss.n5429 dvss.n5151 9.3005
R20229 dvss.n5428 dvss.n5152 9.3005
R20230 dvss.n5425 dvss.n5165 9.3005
R20231 dvss.n5424 dvss.n5166 9.3005
R20232 dvss.n5421 dvss.n5167 9.3005
R20233 dvss.n5420 dvss.n5168 9.3005
R20234 dvss.n5417 dvss.n5169 9.3005
R20235 dvss.n5416 dvss.n5170 9.3005
R20236 dvss.n5413 dvss.n5171 9.3005
R20237 dvss.n5412 dvss.n5177 9.3005
R20238 dvss.n5409 dvss.n5178 9.3005
R20239 dvss.n5408 dvss.n5179 9.3005
R20240 dvss.n5405 dvss.n5180 9.3005
R20241 dvss.n5404 dvss.n5181 9.3005
R20242 dvss.n5401 dvss.n5182 9.3005
R20243 dvss.n5400 dvss.n5183 9.3005
R20244 dvss.n5397 dvss.n5184 9.3005
R20245 dvss.n5396 dvss.n5185 9.3005
R20246 dvss.n5393 dvss.n5186 9.3005
R20247 dvss.n5392 dvss.n5187 9.3005
R20248 dvss.n5389 dvss.n5188 9.3005
R20249 dvss.n5388 dvss.n5189 9.3005
R20250 dvss.n5385 dvss.n5190 9.3005
R20251 dvss.n5384 dvss.n5191 9.3005
R20252 dvss.n5381 dvss.n5204 9.3005
R20253 dvss.n5380 dvss.n5205 9.3005
R20254 dvss.n5377 dvss.n5206 9.3005
R20255 dvss.n5376 dvss.n5207 9.3005
R20256 dvss.n5373 dvss.n5208 9.3005
R20257 dvss.n5372 dvss.n5209 9.3005
R20258 dvss.n5369 dvss.n5210 9.3005
R20259 dvss.n5368 dvss.n5216 9.3005
R20260 dvss.n5365 dvss.n5217 9.3005
R20261 dvss.n5364 dvss.n5218 9.3005
R20262 dvss.n5361 dvss.n5219 9.3005
R20263 dvss.n5360 dvss.n5220 9.3005
R20264 dvss.n5357 dvss.n5221 9.3005
R20265 dvss.n5356 dvss.n5222 9.3005
R20266 dvss.n5353 dvss.n5223 9.3005
R20267 dvss.n5352 dvss.n5224 9.3005
R20268 dvss.n5349 dvss.n5225 9.3005
R20269 dvss.n5348 dvss.n5226 9.3005
R20270 dvss.n5345 dvss.n5227 9.3005
R20271 dvss.n5344 dvss.n5228 9.3005
R20272 dvss.n5341 dvss.n5229 9.3005
R20273 dvss.n5340 dvss.n5230 9.3005
R20274 dvss.n5337 dvss.n5243 9.3005
R20275 dvss.n5336 dvss.n5244 9.3005
R20276 dvss.n5333 dvss.n5245 9.3005
R20277 dvss.n5332 dvss.n5246 9.3005
R20278 dvss.n5329 dvss.n5247 9.3005
R20279 dvss.n5328 dvss.n5248 9.3005
R20280 dvss.n5325 dvss.n5249 9.3005
R20281 dvss.n5324 dvss.n5255 9.3005
R20282 dvss.n5321 dvss.n5256 9.3005
R20283 dvss.n5320 dvss.n5257 9.3005
R20284 dvss.n5317 dvss.n5258 9.3005
R20285 dvss.n5316 dvss.n5259 9.3005
R20286 dvss.n5313 dvss.n5260 9.3005
R20287 dvss.n5312 dvss.n5261 9.3005
R20288 dvss.n5309 dvss.n5262 9.3005
R20289 dvss.n5308 dvss.n5263 9.3005
R20290 dvss.n5305 dvss.n5264 9.3005
R20291 dvss.n5304 dvss.n5265 9.3005
R20292 dvss.n5301 dvss.n5266 9.3005
R20293 dvss.n5300 dvss.n5267 9.3005
R20294 dvss.n5297 dvss.n5268 9.3005
R20295 dvss.n5296 dvss.n5269 9.3005
R20296 dvss.n5293 dvss.n5282 9.3005
R20297 dvss.n5292 dvss.n5283 9.3005
R20298 dvss.n5289 dvss.n5284 9.3005
R20299 dvss.n5288 dvss.n5286 9.3005
R20300 dvss.n5285 dvss.n1149 9.3005
R20301 dvss.n5499 dvss.n5498 9.3005
R20302 dvss.n1150 dvss.n1148 9.3005
R20303 dvss.n5505 dvss.n1147 9.3005
R20304 dvss.n5508 dvss.n5507 9.3005
R20305 dvss.n5506 dvss.n1143 9.3005
R20306 dvss.n5515 dvss.n5514 9.3005
R20307 dvss.n5516 dvss.n1142 9.3005
R20308 dvss.n5519 dvss.n5518 9.3005
R20309 dvss.n5517 dvss.n1138 9.3005
R20310 dvss.n5526 dvss.n5525 9.3005
R20311 dvss.n5527 dvss.n1126 9.3005
R20312 dvss.n5607 dvss.n1127 9.3005
R20313 dvss.n5606 dvss.n1128 9.3005
R20314 dvss.n5605 dvss.n1129 9.3005
R20315 dvss.n5530 dvss.n1130 9.3005
R20316 dvss.n5599 dvss.n1134 9.3005
R20317 dvss.n5598 dvss.n1135 9.3005
R20318 dvss.n5597 dvss.n5539 9.3005
R20319 dvss.n5545 dvss.n5540 9.3005
R20320 dvss.n5591 dvss.n5546 9.3005
R20321 dvss.n5590 dvss.n5547 9.3005
R20322 dvss.n5589 dvss.n5548 9.3005
R20323 dvss.n5553 dvss.n5549 9.3005
R20324 dvss.n5583 dvss.n5552 9.3005
R20325 dvss.n5582 dvss.n5559 9.3005
R20326 dvss.n5581 dvss.n5560 9.3005
R20327 dvss.n5566 dvss.n5561 9.3005
R20328 dvss.n5575 dvss.n5567 9.3005
R20329 dvss.n5574 dvss.n5568 9.3005
R20330 dvss.n5573 dvss.n5570 9.3005
R20331 dvss.n5569 dvss.n522 9.3005
R20332 dvss.n6212 dvss.n6211 9.3005
R20333 dvss.n6214 dvss.n521 9.3005
R20334 dvss.n6218 dvss.n6217 9.3005
R20335 dvss.n6216 dvss.n514 9.3005
R20336 dvss.n6227 dvss.n6226 9.3005
R20337 dvss.n517 dvss.n516 9.3005
R20338 dvss.n515 dvss.n509 9.3005
R20339 dvss.n6236 dvss.n6235 9.3005
R20340 dvss.n6231 dvss.n505 9.3005
R20341 dvss.n6244 dvss.n6243 9.3005
R20342 dvss.n6245 dvss.n504 9.3005
R20343 dvss.n6248 dvss.n6247 9.3005
R20344 dvss.n6246 dvss.n500 9.3005
R20345 dvss.n6256 dvss.n6255 9.3005
R20346 dvss.n499 dvss.n498 9.3005
R20347 dvss.n6264 dvss.n6263 9.3005
R20348 dvss.n6262 dvss.n495 9.3005
R20349 dvss.n6271 dvss.n6270 9.3005
R20350 dvss.n6272 dvss.n494 9.3005
R20351 dvss.n6275 dvss.n6274 9.3005
R20352 dvss.n6273 dvss.n490 9.3005
R20353 dvss.n6283 dvss.n6282 9.3005
R20354 dvss.n6284 dvss.n489 9.3005
R20355 dvss.n6289 dvss.n6288 9.3005
R20356 dvss.n6286 dvss.n485 9.3005
R20357 dvss.n6296 dvss.n6295 9.3005
R20358 dvss.n6297 dvss.n479 9.3005
R20359 dvss.n6306 dvss.n6305 9.3005
R20360 dvss.n6304 dvss.n480 9.3005
R20361 dvss.n6303 dvss.n475 9.3005
R20362 dvss.n6318 dvss.n6317 9.3005
R20363 dvss.n6319 dvss.n472 9.3005
R20364 dvss.n6321 dvss.n6320 9.3005
R20365 dvss.n6323 dvss.n6322 9.3005
R20366 dvss.n6332 dvss.n6331 9.3005
R20367 dvss.n6330 dvss.n471 9.3005
R20368 dvss.n6326 dvss.n468 9.3005
R20369 dvss.n459 dvss.n458 9.3005
R20370 dvss.n6578 dvss.n6577 9.3005
R20371 dvss.n6576 dvss.n6575 9.3005
R20372 dvss.n6574 dvss.n462 9.3005
R20373 dvss.n6573 dvss.n6572 9.3005
R20374 dvss.n6571 dvss.n464 9.3005
R20375 dvss.n6345 dvss.n465 9.3005
R20376 dvss.n6565 dvss.n6564 9.3005
R20377 dvss.n6559 dvss.n230 9.3005
R20378 dvss.n6644 dvss.n231 9.3005
R20379 dvss.n6643 dvss.n232 9.3005
R20380 dvss.n6642 dvss.n233 9.3005
R20381 dvss.n6353 dvss.n234 9.3005
R20382 dvss.n6356 dvss.n6355 9.3005
R20383 dvss.n6354 dvss.n6350 9.3005
R20384 dvss.n6555 dvss.n6554 9.3005
R20385 dvss.n6365 dvss.n6351 9.3005
R20386 dvss.n6548 dvss.n6366 9.3005
R20387 dvss.n6547 dvss.n6367 9.3005
R20388 dvss.n6546 dvss.n6368 9.3005
R20389 dvss.n6373 dvss.n6369 9.3005
R20390 dvss.n6540 dvss.n6372 9.3005
R20391 dvss.n6539 dvss.n6379 9.3005
R20392 dvss.n6538 dvss.n6380 9.3005
R20393 dvss.n6386 dvss.n6381 9.3005
R20394 dvss.n6532 dvss.n6387 9.3005
R20395 dvss.n6531 dvss.n6388 9.3005
R20396 dvss.n6530 dvss.n6389 9.3005
R20397 dvss.n6394 dvss.n6390 9.3005
R20398 dvss.n6524 dvss.n6395 9.3005
R20399 dvss.n6523 dvss.n6396 9.3005
R20400 dvss.n6522 dvss.n6397 9.3005
R20401 dvss.n6417 dvss.n6398 9.3005
R20402 dvss.n6418 dvss.n6402 9.3005
R20403 dvss.n6515 dvss.n6403 9.3005
R20404 dvss.n6514 dvss.n6404 9.3005
R20405 dvss.n6513 dvss.n6405 9.3005
R20406 dvss.n6425 dvss.n6406 9.3005
R20407 dvss.n6507 dvss.n6426 9.3005
R20408 dvss.n6506 dvss.n6427 9.3005
R20409 dvss.n6505 dvss.n6428 9.3005
R20410 dvss.n1700 dvss.n1598 9.3005
R20411 dvss.n1752 dvss.n1599 9.3005
R20412 dvss.n1751 dvss.n1600 9.3005
R20413 dvss.n1750 dvss.n1601 9.3005
R20414 dvss.n1749 dvss.n1602 9.3005
R20415 dvss.n1747 dvss.n1603 9.3005
R20416 dvss.n1744 dvss.n1604 9.3005
R20417 dvss.n1743 dvss.n1605 9.3005
R20418 dvss.n1740 dvss.n1606 9.3005
R20419 dvss.n1739 dvss.n1607 9.3005
R20420 dvss.n1736 dvss.n1735 9.3005
R20421 dvss.n1620 dvss.n1566 9.3005
R20422 dvss.n1758 dvss.n1757 9.3005
R20423 dvss.n1567 dvss.n1563 9.3005
R20424 dvss.n1583 dvss.n1582 9.3005
R20425 dvss.n1585 dvss.n1580 9.3005
R20426 dvss.n1589 dvss.n1588 9.3005
R20427 dvss.n1777 dvss.n1554 9.3005
R20428 dvss.n1553 dvss.n1552 9.3005
R20429 dvss.n1790 dvss.n1789 9.3005
R20430 dvss.n1784 dvss.n1547 9.3005
R20431 dvss.n1800 dvss.n1799 9.3005
R20432 dvss.n1803 dvss.n1542 9.3005
R20433 dvss.n1812 dvss.n1811 9.3005
R20434 dvss.n1543 dvss.n1536 9.3005
R20435 dvss.n1823 dvss.n1822 9.3005
R20436 dvss.n1826 dvss.n1532 9.3005
R20437 dvss.n1832 dvss.n1831 9.3005
R20438 dvss.n1838 dvss.n1527 9.3005
R20439 dvss.n1846 dvss.n1845 9.3005
R20440 dvss.n1860 dvss.n1516 9.3005
R20441 dvss.n1857 dvss.n1855 9.3005
R20442 dvss.n1856 dvss.n1510 9.3005
R20443 dvss.n1867 dvss.n1866 9.3005
R20444 dvss.n1870 dvss.n1868 9.3005
R20445 dvss.n1869 dvss.n1505 9.3005
R20446 dvss.n1884 dvss.n1496 9.3005
R20447 dvss.n1883 dvss.n1497 9.3005
R20448 dvss.n1882 dvss.n1881 9.3005
R20449 dvss.n1892 dvss.n1488 9.3005
R20450 dvss.n1500 dvss.n1487 9.3005
R20451 dvss.n1898 dvss.n1483 9.3005
R20452 dvss.n1905 dvss.n1904 9.3005
R20453 dvss.n1911 dvss.n1479 9.3005
R20454 dvss.n1918 dvss.n1917 9.3005
R20455 dvss.n1926 dvss.n1476 9.3005
R20456 dvss.n1477 dvss.n1473 9.3005
R20457 dvss.n1937 dvss.n1466 9.3005
R20458 dvss.n1938 dvss.n1460 9.3005
R20459 dvss.n1982 dvss.n1981 9.3005
R20460 dvss.n1978 dvss.n1461 9.3005
R20461 dvss.n1977 dvss.n1945 9.3005
R20462 dvss.n1953 dvss.n1948 9.3005
R20463 dvss.n1967 dvss.n1949 9.3005
R20464 dvss.n1964 dvss.n1454 9.3005
R20465 dvss.n2021 dvss.n2020 9.3005
R20466 dvss.n2025 dvss.n1444 9.3005
R20467 dvss.n2053 dvss.n2052 9.3005
R20468 dvss.n2049 dvss.n1445 9.3005
R20469 dvss.n2048 dvss.n2029 9.3005
R20470 dvss.n2047 dvss.n2035 9.3005
R20471 dvss.n2040 dvss.n1433 9.3005
R20472 dvss.n2062 dvss.n2061 9.3005
R20473 dvss.n2064 dvss.n2063 9.3005
R20474 dvss.n2066 dvss.n1429 9.3005
R20475 dvss.n2073 dvss.n2072 9.3005
R20476 dvss.n2079 dvss.n1425 9.3005
R20477 dvss.n1426 dvss.n1421 9.3005
R20478 dvss.n2089 dvss.n1412 9.3005
R20479 dvss.n1413 dvss.n1353 9.3005
R20480 dvss.n2102 dvss.n2101 9.3005
R20481 dvss.n2098 dvss.n1354 9.3005
R20482 dvss.n1377 dvss.n1376 9.3005
R20483 dvss.n1384 dvss.n1383 9.3005
R20484 dvss.n1389 dvss.n1370 9.3005
R20485 dvss.n1373 dvss.n1366 9.3005
R20486 dvss.n1399 dvss.n1361 9.3005
R20487 dvss.n1405 dvss.n893 9.3005
R20488 dvss.n5728 dvss.n5727 9.3005
R20489 dvss.n5724 dvss.n894 9.3005
R20490 dvss.n5723 dvss.n899 9.3005
R20491 dvss.n5722 dvss.n900 9.3005
R20492 dvss.n5719 dvss.n904 9.3005
R20493 dvss.n5718 dvss.n905 9.3005
R20494 dvss.n998 dvss.n908 9.3005
R20495 dvss.n5714 dvss.n909 9.3005
R20496 dvss.n5711 dvss.n914 9.3005
R20497 dvss.n995 dvss.n994 9.3005
R20498 dvss.n997 dvss.n996 9.3005
R20499 dvss.n5705 dvss.n920 9.3005
R20500 dvss.n5702 dvss.n925 9.3005
R20501 dvss.n5701 dvss.n926 9.3005
R20502 dvss.n991 dvss.n927 9.3005
R20503 dvss.n5694 dvss.n929 9.3005
R20504 dvss.n5691 dvss.n934 9.3005
R20505 dvss.n5690 dvss.n935 9.3005
R20506 dvss.n979 dvss.n938 9.3005
R20507 dvss.n1045 dvss.n1044 9.3005
R20508 dvss.n987 dvss.n980 9.3005
R20509 dvss.n981 dvss.n975 9.3005
R20510 dvss.n5678 dvss.n944 9.3005
R20511 dvss.n5675 dvss.n949 9.3005
R20512 dvss.n5674 dvss.n950 9.3005
R20513 dvss.n5673 dvss.n951 9.3005
R20514 dvss.n969 dvss.n968 9.3005
R20515 dvss.n1062 dvss.n956 9.3005
R20516 dvss.n1063 dvss.n957 9.3005
R20517 dvss.n5659 dvss.n963 9.3005
R20518 dvss.n5658 dvss.n1064 9.3005
R20519 dvss.n5657 dvss.n1065 9.3005
R20520 dvss.n1091 dvss.n1066 9.3005
R20521 dvss.n5651 dvss.n1073 9.3005
R20522 dvss.n5650 dvss.n1074 9.3005
R20523 dvss.n5649 dvss.n5648 9.3005
R20524 dvss.n5645 dvss.n1076 9.3005
R20525 dvss.n1115 dvss.n1114 9.3005
R20526 dvss.n5640 dvss.n1101 9.3005
R20527 dvss.n5637 dvss.n1105 9.3005
R20528 dvss.n1112 dvss.n1108 9.3005
R20529 dvss.n5627 dvss.n1109 9.3005
R20530 dvss.n5624 dvss.n804 9.3005
R20531 dvss.n6124 dvss.n6123 9.3005
R20532 dvss.n6128 dvss.n794 9.3005
R20533 dvss.n6156 dvss.n6155 9.3005
R20534 dvss.n6152 dvss.n795 9.3005
R20535 dvss.n6151 dvss.n6132 9.3005
R20536 dvss.n6150 dvss.n6138 9.3005
R20537 dvss.n6143 dvss.n783 9.3005
R20538 dvss.n6165 dvss.n6164 9.3005
R20539 dvss.n6167 dvss.n6166 9.3005
R20540 dvss.n6169 dvss.n779 9.3005
R20541 dvss.n6176 dvss.n6175 9.3005
R20542 dvss.n6182 dvss.n775 9.3005
R20543 dvss.n776 dvss.n771 9.3005
R20544 dvss.n6192 dvss.n762 9.3005
R20545 dvss.n763 dvss.n530 9.3005
R20546 dvss.n6205 dvss.n6204 9.3005
R20547 dvss.n6201 dvss.n531 9.3005
R20548 dvss.n627 dvss.n626 9.3005
R20549 dvss.n636 dvss.n635 9.3005
R20550 dvss.n641 dvss.n615 9.3005
R20551 dvss.n645 dvss.n644 9.3005
R20552 dvss.n618 dvss.n616 9.3005
R20553 dvss.n617 dvss.n611 9.3005
R20554 dvss.n755 dvss.n539 9.3005
R20555 dvss.n752 dvss.n544 9.3005
R20556 dvss.n751 dvss.n545 9.3005
R20557 dvss.n750 dvss.n546 9.3005
R20558 dvss.n747 dvss.n550 9.3005
R20559 dvss.n746 dvss.n551 9.3005
R20560 dvss.n606 dvss.n554 9.3005
R20561 dvss.n742 dvss.n555 9.3005
R20562 dvss.n739 dvss.n560 9.3005
R20563 dvss.n603 dvss.n602 9.3005
R20564 dvss.n605 dvss.n604 9.3005
R20565 dvss.n733 dvss.n566 9.3005
R20566 dvss.n730 dvss.n571 9.3005
R20567 dvss.n729 dvss.n572 9.3005
R20568 dvss.n599 dvss.n573 9.3005
R20569 dvss.n722 dvss.n575 9.3005
R20570 dvss.n719 dvss.n580 9.3005
R20571 dvss.n718 dvss.n581 9.3005
R20572 dvss.n594 dvss.n584 9.3005
R20573 dvss.n596 dvss.n595 9.3005
R20574 dvss.n705 dvss.n589 9.3005
R20575 dvss.n706 dvss.n127 9.3005
R20576 dvss.n6712 dvss.n6711 9.3005
R20577 dvss.n6708 dvss.n128 9.3005
R20578 dvss.n6707 dvss.n133 9.3005
R20579 dvss.n6706 dvss.n134 9.3005
R20580 dvss.n6703 dvss.n138 9.3005
R20581 dvss.n6702 dvss.n139 9.3005
R20582 dvss.n204 dvss.n142 9.3005
R20583 dvss.n6698 dvss.n143 9.3005
R20584 dvss.n6695 dvss.n148 9.3005
R20585 dvss.n212 dvss.n211 9.3005
R20586 dvss.n214 dvss.n213 9.3005
R20587 dvss.n6689 dvss.n154 9.3005
R20588 dvss.n6686 dvss.n159 9.3005
R20589 dvss.n6685 dvss.n160 9.3005
R20590 dvss.n181 dvss.n161 9.3005
R20591 dvss.n6678 dvss.n163 9.3005
R20592 dvss.n6675 dvss.n171 9.3005
R20593 dvss.n6674 dvss.n172 9.3005
R20594 dvss.n180 dvss.n175 9.3005
R20595 dvss.n6664 dvss.n176 9.3005
R20596 dvss.n6661 dvss.n75 9.3005
R20597 dvss.n6865 dvss.n6864 9.3005
R20598 dvss.n6869 dvss.n70 9.3005
R20599 dvss.n6897 dvss.n6896 9.3005
R20600 dvss.n6893 dvss.n71 9.3005
R20601 dvss.n6892 dvss.n6873 9.3005
R20602 dvss.n6891 dvss.n6879 9.3005
R20603 dvss.n6884 dvss.n59 9.3005
R20604 dvss.n6906 dvss.n6905 9.3005
R20605 dvss.n6908 dvss.n6907 9.3005
R20606 dvss.n6910 dvss.n55 9.3005
R20607 dvss.n6917 dvss.n6916 9.3005
R20608 dvss.n6923 dvss.n51 9.3005
R20609 dvss.n52 dvss.n47 9.3005
R20610 dvss.n6933 dvss.n38 9.3005
R20611 dvss.n39 dvss.n28 9.3005
R20612 dvss.n6946 dvss.n6945 9.3005
R20613 dvss.n6942 dvss.n29 9.3005
R20614 dvss.n6457 dvss.n6456 9.3005
R20615 dvss.n6463 dvss.n6447 9.3005
R20616 dvss.n6469 dvss.n6468 9.3005
R20617 dvss.n6475 dvss.n6443 9.3005
R20618 dvss.n6477 dvss.n6476 9.3005
R20619 dvss.n6483 dvss.n6439 9.3005
R20620 dvss.n6488 dvss.n6487 9.3005
R20621 dvss.n6494 dvss.n6433 9.3005
R20622 dvss.n6496 dvss.n6495 9.3005
R20623 dvss.n6498 dvss.n6497 9.3005
R20624 dvss.n3200 dvss.n3195 9.3005
R20625 dvss.n3204 dvss.n3203 9.3005
R20626 dvss.n3202 dvss.n3191 9.3005
R20627 dvss.n3211 dvss.n3210 9.3005
R20628 dvss.n3212 dvss.n3187 9.3005
R20629 dvss.n3219 dvss.n3218 9.3005
R20630 dvss.n3188 dvss.n3183 9.3005
R20631 dvss.n3227 dvss.n3226 9.3005
R20632 dvss.n3182 dvss.n3177 9.3005
R20633 dvss.n3234 dvss.n3233 9.3005
R20634 dvss.n3179 dvss.n3174 9.3005
R20635 dvss.n3243 dvss.n3242 9.3005
R20636 dvss.n3244 dvss.n3169 9.3005
R20637 dvss.n3250 dvss.n3249 9.3005
R20638 dvss.n3171 dvss.n3166 9.3005
R20639 dvss.n3257 dvss.n3256 9.3005
R20640 dvss.n3258 dvss.n3164 9.3005
R20641 dvss.n3262 dvss.n3261 9.3005
R20642 dvss.n3260 dvss.n3165 9.3005
R20643 dvss.n3259 dvss.n240 9.3005
R20644 dvss.n6635 dvss.n6634 9.3005
R20645 dvss.n1699 dvss.n1691 9.3005
R20646 dvss.n1703 dvss.n1702 9.3005
R20647 dvss.n1727 dvss.n1704 9.3005
R20648 dvss.n1726 dvss.n1705 9.3005
R20649 dvss.n1725 dvss.n1706 9.3005
R20650 dvss.n1724 dvss.n1707 9.3005
R20651 dvss.n1722 dvss.n1708 9.3005
R20652 dvss.n1719 dvss.n1712 9.3005
R20653 dvss.n1718 dvss.n1713 9.3005
R20654 dvss.n1715 dvss.n1714 9.3005
R20655 dvss.n1619 dvss.n1618 9.3005
R20656 dvss.n1734 dvss.n1733 9.3005
R20657 dvss.n1622 dvss.n1621 9.3005
R20658 dvss.n1759 dvss.n1561 9.3005
R20659 dvss.n1769 dvss.n1768 9.3005
R20660 dvss.n1584 dvss.n1562 9.3005
R20661 dvss.n1587 dvss.n1586 9.3005
R20662 dvss.n1588 dvss.n1555 9.3005
R20663 dvss.n1777 dvss.n1776 9.3005
R20664 dvss.n1775 dvss.n1553 9.3005
R20665 dvss.n1789 dvss.n1550 9.3005
R20666 dvss.n1784 dvss.n1545 9.3005
R20667 dvss.n1801 dvss.n1800 9.3005
R20668 dvss.n1803 dvss.n1802 9.3005
R20669 dvss.n1811 dvss.n1540 9.3005
R20670 dvss.n1543 dvss.n1534 9.3005
R20671 dvss.n1824 dvss.n1823 9.3005
R20672 dvss.n1826 dvss.n1825 9.3005
R20673 dvss.n1831 dvss.n1528 9.3005
R20674 dvss.n1838 dvss.n1837 9.3005
R20675 dvss.n1845 dvss.n1518 9.3005
R20676 dvss.n1860 dvss.n1859 9.3005
R20677 dvss.n1858 dvss.n1857 9.3005
R20678 dvss.n1856 dvss.n1521 9.3005
R20679 dvss.n1866 dvss.n1508 9.3005
R20680 dvss.n1871 dvss.n1870 9.3005
R20681 dvss.n1869 dvss.n1494 9.3005
R20682 dvss.n1885 dvss.n1884 9.3005
R20683 dvss.n1883 dvss.n1495 9.3005
R20684 dvss.n1882 dvss.n1489 9.3005
R20685 dvss.n1892 dvss.n1891 9.3005
R20686 dvss.n1487 dvss.n1486 9.3005
R20687 dvss.n1899 dvss.n1898 9.3005
R20688 dvss.n1905 dvss.n1482 9.3005
R20689 dvss.n1912 dvss.n1911 9.3005
R20690 dvss.n1918 dvss.n1475 9.3005
R20691 dvss.n1927 dvss.n1926 9.3005
R20692 dvss.n1477 dvss.n1467 9.3005
R20693 dvss.n1937 dvss.n1936 9.3005
R20694 dvss.n1938 dvss.n1462 9.3005
R20695 dvss.n1981 dvss.n1980 9.3005
R20696 dvss.n1979 dvss.n1978 9.3005
R20697 dvss.n1977 dvss.n1464 9.3005
R20698 dvss.n1950 dvss.n1948 9.3005
R20699 dvss.n1967 dvss.n1966 9.3005
R20700 dvss.n1965 dvss.n1964 9.3005
R20701 dvss.n2021 dvss.n1446 9.3005
R20702 dvss.n2026 dvss.n2025 9.3005
R20703 dvss.n2052 dvss.n2051 9.3005
R20704 dvss.n2050 dvss.n2049 9.3005
R20705 dvss.n2048 dvss.n2028 9.3005
R20706 dvss.n2047 dvss.n2046 9.3005
R20707 dvss.n2040 dvss.n1436 9.3005
R20708 dvss.n2061 dvss.n2060 9.3005
R20709 dvss.n2064 dvss.n1432 9.3005
R20710 dvss.n2067 dvss.n2066 9.3005
R20711 dvss.n2073 dvss.n1424 9.3005
R20712 dvss.n2080 dvss.n2079 9.3005
R20713 dvss.n1426 dvss.n1414 9.3005
R20714 dvss.n2089 dvss.n2088 9.3005
R20715 dvss.n1413 dvss.n1356 9.3005
R20716 dvss.n2101 dvss.n2100 9.3005
R20717 dvss.n2099 dvss.n2098 9.3005
R20718 dvss.n1376 dvss.n1358 9.3005
R20719 dvss.n1384 dvss.n1368 9.3005
R20720 dvss.n1390 dvss.n1389 9.3005
R20721 dvss.n1373 dvss.n1362 9.3005
R20722 dvss.n1399 dvss.n1398 9.3005
R20723 dvss.n1405 dvss.n896 9.3005
R20724 dvss.n5727 dvss.n5726 9.3005
R20725 dvss.n5725 dvss.n5724 9.3005
R20726 dvss.n5723 dvss.n898 9.3005
R20727 dvss.n5722 dvss.n5721 9.3005
R20728 dvss.n5720 dvss.n5719 9.3005
R20729 dvss.n5718 dvss.n903 9.3005
R20730 dvss.n910 dvss.n908 9.3005
R20731 dvss.n5714 dvss.n5713 9.3005
R20732 dvss.n5712 dvss.n5711 9.3005
R20733 dvss.n995 dvss.n913 9.3005
R20734 dvss.n996 dvss.n921 9.3005
R20735 dvss.n5705 dvss.n5704 9.3005
R20736 dvss.n5703 dvss.n5702 9.3005
R20737 dvss.n5701 dvss.n924 9.3005
R20738 dvss.n930 dvss.n927 9.3005
R20739 dvss.n5694 dvss.n5693 9.3005
R20740 dvss.n5692 dvss.n5691 9.3005
R20741 dvss.n5690 dvss.n933 9.3005
R20742 dvss.n1042 dvss.n938 9.3005
R20743 dvss.n1044 dvss.n1043 9.3005
R20744 dvss.n987 dvss.n977 9.3005
R20745 dvss.n981 dvss.n945 9.3005
R20746 dvss.n5678 dvss.n5677 9.3005
R20747 dvss.n5676 dvss.n5675 9.3005
R20748 dvss.n5674 dvss.n948 9.3005
R20749 dvss.n5673 dvss.n5672 9.3005
R20750 dvss.n968 dvss.n955 9.3005
R20751 dvss.n5665 dvss.n956 9.3005
R20752 dvss.n5664 dvss.n957 9.3005
R20753 dvss.n5663 dvss.n963 9.3005
R20754 dvss.n1064 dvss.n964 9.3005
R20755 dvss.n1088 dvss.n1065 9.3005
R20756 dvss.n1091 dvss.n1090 9.3005
R20757 dvss.n1089 dvss.n1073 9.3005
R20758 dvss.n1077 dvss.n1074 9.3005
R20759 dvss.n5648 dvss.n5647 9.3005
R20760 dvss.n5646 dvss.n5645 9.3005
R20761 dvss.n1114 dvss.n1080 9.3005
R20762 dvss.n5640 dvss.n5639 9.3005
R20763 dvss.n5638 dvss.n5637 9.3005
R20764 dvss.n1108 dvss.n1104 9.3005
R20765 dvss.n5627 dvss.n5626 9.3005
R20766 dvss.n5625 dvss.n5624 9.3005
R20767 dvss.n6124 dvss.n796 9.3005
R20768 dvss.n6129 dvss.n6128 9.3005
R20769 dvss.n6155 dvss.n6154 9.3005
R20770 dvss.n6153 dvss.n6152 9.3005
R20771 dvss.n6151 dvss.n6131 9.3005
R20772 dvss.n6150 dvss.n6149 9.3005
R20773 dvss.n6143 dvss.n786 9.3005
R20774 dvss.n6164 dvss.n6163 9.3005
R20775 dvss.n6167 dvss.n782 9.3005
R20776 dvss.n6170 dvss.n6169 9.3005
R20777 dvss.n6176 dvss.n774 9.3005
R20778 dvss.n6183 dvss.n6182 9.3005
R20779 dvss.n776 dvss.n764 9.3005
R20780 dvss.n6192 dvss.n6191 9.3005
R20781 dvss.n763 dvss.n533 9.3005
R20782 dvss.n6204 dvss.n6203 9.3005
R20783 dvss.n6202 dvss.n6201 9.3005
R20784 dvss.n626 dvss.n535 9.3005
R20785 dvss.n636 dvss.n619 9.3005
R20786 dvss.n642 dvss.n641 9.3005
R20787 dvss.n644 dvss.n643 9.3005
R20788 dvss.n618 dvss.n613 9.3005
R20789 dvss.n617 dvss.n540 9.3005
R20790 dvss.n755 dvss.n754 9.3005
R20791 dvss.n753 dvss.n752 9.3005
R20792 dvss.n751 dvss.n543 9.3005
R20793 dvss.n750 dvss.n749 9.3005
R20794 dvss.n748 dvss.n747 9.3005
R20795 dvss.n746 dvss.n549 9.3005
R20796 dvss.n556 dvss.n554 9.3005
R20797 dvss.n742 dvss.n741 9.3005
R20798 dvss.n740 dvss.n739 9.3005
R20799 dvss.n603 dvss.n559 9.3005
R20800 dvss.n604 dvss.n567 9.3005
R20801 dvss.n733 dvss.n732 9.3005
R20802 dvss.n731 dvss.n730 9.3005
R20803 dvss.n729 dvss.n570 9.3005
R20804 dvss.n576 dvss.n573 9.3005
R20805 dvss.n722 dvss.n721 9.3005
R20806 dvss.n720 dvss.n719 9.3005
R20807 dvss.n718 dvss.n579 9.3005
R20808 dvss.n696 dvss.n584 9.3005
R20809 dvss.n595 dvss.n590 9.3005
R20810 dvss.n705 dvss.n704 9.3005
R20811 dvss.n706 dvss.n130 9.3005
R20812 dvss.n6711 dvss.n6710 9.3005
R20813 dvss.n6709 dvss.n6708 9.3005
R20814 dvss.n6707 dvss.n132 9.3005
R20815 dvss.n6706 dvss.n6705 9.3005
R20816 dvss.n6704 dvss.n6703 9.3005
R20817 dvss.n6702 dvss.n137 9.3005
R20818 dvss.n144 dvss.n142 9.3005
R20819 dvss.n6698 dvss.n6697 9.3005
R20820 dvss.n6696 dvss.n6695 9.3005
R20821 dvss.n212 dvss.n147 9.3005
R20822 dvss.n213 dvss.n155 9.3005
R20823 dvss.n6689 dvss.n6688 9.3005
R20824 dvss.n6687 dvss.n6686 9.3005
R20825 dvss.n6685 dvss.n158 9.3005
R20826 dvss.n164 dvss.n161 9.3005
R20827 dvss.n6678 dvss.n6677 9.3005
R20828 dvss.n6676 dvss.n6675 9.3005
R20829 dvss.n6674 dvss.n167 9.3005
R20830 dvss.n177 dvss.n175 9.3005
R20831 dvss.n6664 dvss.n6663 9.3005
R20832 dvss.n6662 dvss.n6661 9.3005
R20833 dvss.n6865 dvss.n72 9.3005
R20834 dvss.n6870 dvss.n6869 9.3005
R20835 dvss.n6896 dvss.n6895 9.3005
R20836 dvss.n6894 dvss.n6893 9.3005
R20837 dvss.n6892 dvss.n6872 9.3005
R20838 dvss.n6891 dvss.n6890 9.3005
R20839 dvss.n6884 dvss.n62 9.3005
R20840 dvss.n6905 dvss.n6904 9.3005
R20841 dvss.n6908 dvss.n58 9.3005
R20842 dvss.n6911 dvss.n6910 9.3005
R20843 dvss.n6917 dvss.n50 9.3005
R20844 dvss.n6924 dvss.n6923 9.3005
R20845 dvss.n52 dvss.n40 9.3005
R20846 dvss.n6933 dvss.n6932 9.3005
R20847 dvss.n39 dvss.n31 9.3005
R20848 dvss.n6945 dvss.n6944 9.3005
R20849 dvss.n6943 dvss.n6942 9.3005
R20850 dvss.n6456 dvss.n33 9.3005
R20851 dvss.n6463 dvss.n6462 9.3005
R20852 dvss.n6468 dvss.n6444 9.3005
R20853 dvss.n6475 dvss.n6474 9.3005
R20854 dvss.n6476 dvss.n6440 9.3005
R20855 dvss.n6483 dvss.n6482 9.3005
R20856 dvss.n6487 dvss.n6435 9.3005
R20857 dvss.n6494 dvss.n6493 9.3005
R20858 dvss.n6495 dvss.n6432 9.3005
R20859 dvss.n6499 dvss.n6498 9.3005
R20860 dvss.n2280 dvss.n2279 9.3005
R20861 dvss.n2279 dvss.n1246 9.3005
R20862 dvss.n2264 dvss.n2263 9.3005
R20863 dvss.n2265 dvss.n2264 9.3005
R20864 dvss.n2224 dvss.n2223 9.3005
R20865 dvss.n2222 dvss.n1279 9.3005
R20866 dvss.n2235 dvss.n2234 9.3005
R20867 dvss.n2250 dvss.n2249 9.3005
R20868 dvss.n2244 dvss.n2243 9.3005
R20869 dvss.n2241 dvss.n2240 9.3005
R20870 dvss.n2234 dvss.n2232 9.3005
R20871 dvss.n2174 dvss.n2173 9.3005
R20872 dvss.n2172 dvss.n1310 9.3005
R20873 dvss.n2185 dvss.n2184 9.3005
R20874 dvss.n2200 dvss.n2199 9.3005
R20875 dvss.n2194 dvss.n2193 9.3005
R20876 dvss.n2191 dvss.n2190 9.3005
R20877 dvss.n2184 dvss.n2182 9.3005
R20878 dvss.n2119 dvss.n2118 9.3005
R20879 dvss.n2117 dvss.n1341 9.3005
R20880 dvss.n2130 dvss.n2129 9.3005
R20881 dvss.n2145 dvss.n2144 9.3005
R20882 dvss.n2139 dvss.n2138 9.3005
R20883 dvss.n2136 dvss.n2135 9.3005
R20884 dvss.n2129 dvss.n2127 9.3005
R20885 dvss.n5806 dvss.n5805 9.3005
R20886 dvss.n5809 dvss.n5808 9.3005
R20887 dvss.n5792 dvss.n5791 9.3005
R20888 dvss.n5763 dvss.n5762 9.3005
R20889 dvss.n5775 dvss.n5774 9.3005
R20890 dvss.n5780 dvss.n5779 9.3005
R20891 dvss.n5793 dvss.n5792 9.3005
R20892 dvss.n5886 dvss.n5885 9.3005
R20893 dvss.n820 dvss.n819 9.3005
R20894 dvss.n5870 dvss.n825 9.3005
R20895 dvss.n5853 dvss.n5852 9.3005
R20896 dvss.n5856 dvss.n5855 9.3005
R20897 dvss.n5868 dvss.n5867 9.3005
R20898 dvss.n5871 dvss.n5870 9.3005
R20899 dvss.n6075 dvss.n6074 9.3005
R20900 dvss.n6073 dvss.n5940 9.3005
R20901 dvss.n6086 dvss.n6085 9.3005
R20902 dvss.n6101 dvss.n6100 9.3005
R20903 dvss.n6095 dvss.n6094 9.3005
R20904 dvss.n6092 dvss.n6091 9.3005
R20905 dvss.n6085 dvss.n6083 9.3005
R20906 dvss.n6025 dvss.n6024 9.3005
R20907 dvss.n6023 dvss.n5971 9.3005
R20908 dvss.n6036 dvss.n6035 9.3005
R20909 dvss.n6051 dvss.n6050 9.3005
R20910 dvss.n6045 dvss.n6044 9.3005
R20911 dvss.n6042 dvss.n6041 9.3005
R20912 dvss.n6035 dvss.n6033 9.3005
R20913 dvss.n6780 dvss.n6779 9.3005
R20914 dvss.n91 dvss.n90 9.3005
R20915 dvss.n6764 dvss.n96 9.3005
R20916 dvss.n6747 dvss.n6746 9.3005
R20917 dvss.n6750 dvss.n6749 9.3005
R20918 dvss.n6762 dvss.n6761 9.3005
R20919 dvss.n6765 dvss.n6764 9.3005
R20920 dvss.n6961 dvss.n6960 9.3005
R20921 dvss.n6959 dvss.n6956 9.3005
R20922 dvss.n6827 dvss.n6826 9.3005
R20923 dvss.n6842 dvss.n6841 9.3005
R20924 dvss.n6836 dvss.n6835 9.3005
R20925 dvss.n6833 dvss.n6832 9.3005
R20926 dvss.n6826 dvss.n6824 9.3005
R20927 dvss.n2272 dvss.n2271 9.3005
R20928 dvss.n2273 dvss.n2272 9.3005
R20929 dvss.n7056 dvss.n7055 9.3005
R20930 dvss.n7054 dvss.n7053 9.3005
R20931 dvss.n4 dvss.n3 9.3005
R20932 dvss.n2287 dvss.n2286 9.3005
R20933 dvss.n2285 dvss.n1242 9.3005
R20934 dvss.n2284 dvss.n2283 9.3005
R20935 dvss.n2282 dvss.n2281 9.3005
R20936 dvss.n2278 dvss.n1245 9.3005
R20937 dvss.n2277 dvss.n2276 9.3005
R20938 dvss.n2275 dvss.n2274 9.3005
R20939 dvss.n2270 dvss.n1249 9.3005
R20940 dvss.n2269 dvss.n2268 9.3005
R20941 dvss.n2267 dvss.n2266 9.3005
R20942 dvss.n1256 dvss.n1254 9.3005
R20943 dvss.n2262 dvss.n2261 9.3005
R20944 dvss.n2260 dvss.n2259 9.3005
R20945 dvss.n2258 dvss.n1259 9.3005
R20946 dvss.n2257 dvss.n2256 9.3005
R20947 dvss.n2255 dvss.n2254 9.3005
R20948 dvss.n2253 dvss.n1262 9.3005
R20949 dvss.n1265 dvss.n1264 9.3005
R20950 dvss.n2248 dvss.n2247 9.3005
R20951 dvss.n2246 dvss.n2245 9.3005
R20952 dvss.n1271 dvss.n1268 9.3005
R20953 dvss.n2239 dvss.n2238 9.3005
R20954 dvss.n2237 dvss.n2236 9.3005
R20955 dvss.n1275 dvss.n1274 9.3005
R20956 dvss.n2231 dvss.n2230 9.3005
R20957 dvss.n2229 dvss.n2228 9.3005
R20958 dvss.n2227 dvss.n1278 9.3005
R20959 dvss.n1282 dvss.n1281 9.3005
R20960 dvss.n2221 dvss.n2220 9.3005
R20961 dvss.n2219 dvss.n2218 9.3005
R20962 dvss.n2217 dvss.n1285 9.3005
R20963 dvss.n2216 dvss.n2215 9.3005
R20964 dvss.n2214 dvss.n2213 9.3005
R20965 dvss.n2212 dvss.n1288 9.3005
R20966 dvss.n2211 dvss.n2210 9.3005
R20967 dvss.n2209 dvss.n2208 9.3005
R20968 dvss.n2207 dvss.n1291 9.3005
R20969 dvss.n2206 dvss.n2205 9.3005
R20970 dvss.n2204 dvss.n2203 9.3005
R20971 dvss.n1296 dvss.n1294 9.3005
R20972 dvss.n2198 dvss.n2197 9.3005
R20973 dvss.n2196 dvss.n2195 9.3005
R20974 dvss.n1302 dvss.n1299 9.3005
R20975 dvss.n2189 dvss.n2188 9.3005
R20976 dvss.n2187 dvss.n2186 9.3005
R20977 dvss.n1306 dvss.n1305 9.3005
R20978 dvss.n2181 dvss.n2180 9.3005
R20979 dvss.n2179 dvss.n2178 9.3005
R20980 dvss.n2177 dvss.n1309 9.3005
R20981 dvss.n1313 dvss.n1312 9.3005
R20982 dvss.n2171 dvss.n2170 9.3005
R20983 dvss.n2169 dvss.n2168 9.3005
R20984 dvss.n2162 dvss.n1316 9.3005
R20985 dvss.n2161 dvss.n2160 9.3005
R20986 dvss.n2159 dvss.n2158 9.3005
R20987 dvss.n2157 dvss.n1319 9.3005
R20988 dvss.n2156 dvss.n2155 9.3005
R20989 dvss.n2154 dvss.n2153 9.3005
R20990 dvss.n2152 dvss.n1322 9.3005
R20991 dvss.n2151 dvss.n2150 9.3005
R20992 dvss.n2149 dvss.n2148 9.3005
R20993 dvss.n1327 dvss.n1325 9.3005
R20994 dvss.n2143 dvss.n2142 9.3005
R20995 dvss.n2141 dvss.n2140 9.3005
R20996 dvss.n1333 dvss.n1330 9.3005
R20997 dvss.n2134 dvss.n2133 9.3005
R20998 dvss.n2132 dvss.n2131 9.3005
R20999 dvss.n1337 dvss.n1336 9.3005
R21000 dvss.n2126 dvss.n2125 9.3005
R21001 dvss.n2124 dvss.n2123 9.3005
R21002 dvss.n2122 dvss.n1340 9.3005
R21003 dvss.n1345 dvss.n1343 9.3005
R21004 dvss.n2116 dvss.n2115 9.3005
R21005 dvss.n1344 dvss.n885 9.3005
R21006 dvss.n5736 dvss.n5735 9.3005
R21007 dvss.n5737 dvss.n878 9.3005
R21008 dvss.n5749 dvss.n5748 9.3005
R21009 dvss.n5747 dvss.n879 9.3005
R21010 dvss.n5746 dvss.n5745 9.3005
R21011 dvss.n5744 dvss.n5743 9.3005
R21012 dvss.n5742 dvss.n872 9.3005
R21013 dvss.n5757 dvss.n5756 9.3005
R21014 dvss.n5758 dvss.n870 9.3005
R21015 dvss.n5765 dvss.n5764 9.3005
R21016 dvss.n871 dvss.n866 9.3005
R21017 dvss.n5772 dvss.n5771 9.3005
R21018 dvss.n5773 dvss.n864 9.3005
R21019 dvss.n5783 dvss.n5782 9.3005
R21020 dvss.n5781 dvss.n860 9.3005
R21021 dvss.n5790 dvss.n5789 9.3005
R21022 dvss.n5794 dvss.n859 9.3005
R21023 dvss.n5797 dvss.n5796 9.3005
R21024 dvss.n5795 dvss.n855 9.3005
R21025 dvss.n5804 dvss.n5803 9.3005
R21026 dvss.n5810 dvss.n852 9.3005
R21027 dvss.n5818 dvss.n5817 9.3005
R21028 dvss.n5811 dvss.n847 9.3005
R21029 dvss.n5827 dvss.n5826 9.3005
R21030 dvss.n5828 dvss.n846 9.3005
R21031 dvss.n5831 dvss.n5830 9.3005
R21032 dvss.n5829 dvss.n843 9.3005
R21033 dvss.n5838 dvss.n5837 9.3005
R21034 dvss.n5839 dvss.n842 9.3005
R21035 dvss.n5843 dvss.n5842 9.3005
R21036 dvss.n5841 dvss.n838 9.3005
R21037 dvss.n5850 dvss.n5849 9.3005
R21038 dvss.n5851 dvss.n834 9.3005
R21039 dvss.n5858 dvss.n5857 9.3005
R21040 dvss.n835 dvss.n830 9.3005
R21041 dvss.n5866 dvss.n5865 9.3005
R21042 dvss.n829 dvss.n824 9.3005
R21043 dvss.n5873 dvss.n5872 9.3005
R21044 dvss.n826 dvss.n821 9.3005
R21045 dvss.n5881 dvss.n5880 9.3005
R21046 dvss.n5882 dvss.n816 9.3005
R21047 dvss.n5888 dvss.n5887 9.3005
R21048 dvss.n818 dvss.n813 9.3005
R21049 dvss.n5895 dvss.n5894 9.3005
R21050 dvss.n5901 dvss.n811 9.3005
R21051 dvss.n6116 dvss.n6115 9.3005
R21052 dvss.n6114 dvss.n812 9.3005
R21053 dvss.n6113 dvss.n6112 9.3005
R21054 dvss.n6111 dvss.n6110 9.3005
R21055 dvss.n6109 dvss.n5904 9.3005
R21056 dvss.n6108 dvss.n6107 9.3005
R21057 dvss.n6106 dvss.n6105 9.3005
R21058 dvss.n6104 dvss.n5907 9.3005
R21059 dvss.n5910 dvss.n5909 9.3005
R21060 dvss.n6099 dvss.n6098 9.3005
R21061 dvss.n6097 dvss.n6096 9.3005
R21062 dvss.n5916 dvss.n5913 9.3005
R21063 dvss.n6090 dvss.n6089 9.3005
R21064 dvss.n6088 dvss.n6087 9.3005
R21065 dvss.n5936 dvss.n5935 9.3005
R21066 dvss.n6082 dvss.n6081 9.3005
R21067 dvss.n6080 dvss.n6079 9.3005
R21068 dvss.n6078 dvss.n5939 9.3005
R21069 dvss.n5943 dvss.n5942 9.3005
R21070 dvss.n6072 dvss.n6071 9.3005
R21071 dvss.n6070 dvss.n6069 9.3005
R21072 dvss.n6068 dvss.n5946 9.3005
R21073 dvss.n6067 dvss.n6066 9.3005
R21074 dvss.n6065 dvss.n6064 9.3005
R21075 dvss.n6063 dvss.n5949 9.3005
R21076 dvss.n6062 dvss.n6061 9.3005
R21077 dvss.n6060 dvss.n6059 9.3005
R21078 dvss.n6058 dvss.n5952 9.3005
R21079 dvss.n6057 dvss.n6056 9.3005
R21080 dvss.n6055 dvss.n6054 9.3005
R21081 dvss.n5957 dvss.n5955 9.3005
R21082 dvss.n6049 dvss.n6048 9.3005
R21083 dvss.n6047 dvss.n6046 9.3005
R21084 dvss.n5963 dvss.n5960 9.3005
R21085 dvss.n6040 dvss.n6039 9.3005
R21086 dvss.n6038 dvss.n6037 9.3005
R21087 dvss.n5967 dvss.n5966 9.3005
R21088 dvss.n6032 dvss.n6031 9.3005
R21089 dvss.n6030 dvss.n6029 9.3005
R21090 dvss.n6028 dvss.n5970 9.3005
R21091 dvss.n5974 dvss.n5973 9.3005
R21092 dvss.n6022 dvss.n6021 9.3005
R21093 dvss.n6020 dvss.n6019 9.3005
R21094 dvss.n6018 dvss.n118 9.3005
R21095 dvss.n6721 dvss.n6720 9.3005
R21096 dvss.n6722 dvss.n117 9.3005
R21097 dvss.n6725 dvss.n6724 9.3005
R21098 dvss.n6723 dvss.n114 9.3005
R21099 dvss.n6732 dvss.n6731 9.3005
R21100 dvss.n6733 dvss.n113 9.3005
R21101 dvss.n6737 dvss.n6736 9.3005
R21102 dvss.n6735 dvss.n109 9.3005
R21103 dvss.n6744 dvss.n6743 9.3005
R21104 dvss.n6745 dvss.n105 9.3005
R21105 dvss.n6752 dvss.n6751 9.3005
R21106 dvss.n106 dvss.n101 9.3005
R21107 dvss.n6760 dvss.n6759 9.3005
R21108 dvss.n100 dvss.n95 9.3005
R21109 dvss.n6767 dvss.n6766 9.3005
R21110 dvss.n97 dvss.n92 9.3005
R21111 dvss.n6775 dvss.n6774 9.3005
R21112 dvss.n6776 dvss.n87 9.3005
R21113 dvss.n6782 dvss.n6781 9.3005
R21114 dvss.n89 dvss.n84 9.3005
R21115 dvss.n6789 dvss.n6788 9.3005
R21116 dvss.n6790 dvss.n82 9.3005
R21117 dvss.n6857 dvss.n6856 9.3005
R21118 dvss.n6855 dvss.n83 9.3005
R21119 dvss.n6854 dvss.n6853 9.3005
R21120 dvss.n6852 dvss.n6851 9.3005
R21121 dvss.n6850 dvss.n6793 9.3005
R21122 dvss.n6849 dvss.n6848 9.3005
R21123 dvss.n6847 dvss.n6846 9.3005
R21124 dvss.n6845 dvss.n6796 9.3005
R21125 dvss.n6799 dvss.n6798 9.3005
R21126 dvss.n6840 dvss.n6839 9.3005
R21127 dvss.n6838 dvss.n6837 9.3005
R21128 dvss.n6805 dvss.n6802 9.3005
R21129 dvss.n6831 dvss.n6830 9.3005
R21130 dvss.n6829 dvss.n6828 9.3005
R21131 dvss.n6823 dvss.n21 9.3005
R21132 dvss.n6954 dvss.n6953 9.3005
R21133 dvss.n6955 dvss.n20 9.3005
R21134 dvss.n6965 dvss.n6964 9.3005
R21135 dvss.n6958 dvss.n16 9.3005
R21136 dvss.n6972 dvss.n6971 9.3005
R21137 dvss.n6973 dvss.n14 9.3005
R21138 dvss.n6978 dvss.n6977 9.3005
R21139 dvss.n6976 dvss.n15 9.3005
R21140 dvss.n6975 dvss.n10 9.3005
R21141 dvss.n6974 dvss.n7 9.3005
R21142 dvss.n6988 dvss.n6987 9.3005
R21143 dvss.n2796 dvss.n2795 9.03579
R21144 dvss.n3803 dvss.n3798 9.03579
R21145 dvss.n3823 dvss.n3632 9.03579
R21146 dvss.n4157 dvss.n4151 9.03579
R21147 dvss.n4230 dvss.n4229 9.03579
R21148 dvss.t1638 dvss.n4808 8.72452
R21149 dvss.n4808 dvss.t1599 8.72452
R21150 dvss.n3460 dvss.n3457 8.65932
R21151 dvss.n3496 dvss.n3470 8.65932
R21152 dvss.n1762 dvss.n1760 8.56999
R21153 dvss.n5125 dvss.n5123 8.56999
R21154 dvss.n7049 dvss.n7048 8.56458
R21155 dvss.n3331 dvss.n3130 8.54791
R21156 dvss.n6882 dvss.n6881 8.54791
R21157 dvss.n6700 dvss.n141 8.54791
R21158 dvss.n744 dvss.n553 8.54791
R21159 dvss.n6141 dvss.n6140 8.54791
R21160 dvss.n961 dvss.n960 8.54791
R21161 dvss.n5716 dvss.n907 8.54791
R21162 dvss.n2038 dvss.n2037 8.54791
R21163 dvss.n1896 dvss.n1895 8.54791
R21164 dvss.n1781 dvss.n1780 8.54791
R21165 dvss.n6377 dvss.n6376 8.54791
R21166 dvss.n6328 dvss.n6325 8.54791
R21167 dvss.n6260 dvss.n6259 8.54791
R21168 dvss.n5557 dvss.n5556 8.54791
R21169 dvss.n5503 dvss.n5502 8.54791
R21170 dvss.n5253 dvss.n5252 8.54791
R21171 dvss.n5214 dvss.n5213 8.54791
R21172 dvss.n5175 dvss.n5174 8.54791
R21173 dvss.n5136 dvss.n5135 8.54791
R21174 dvss.n1209 dvss 8.53237
R21175 dvss.n1609 dvss 8.48432
R21176 dvss.n5113 dvss 8.48432
R21177 dvss.n3130 dvss 8.43944
R21178 dvss.n6881 dvss 8.43944
R21179 dvss.n141 dvss 8.43944
R21180 dvss.n553 dvss 8.43944
R21181 dvss.n6140 dvss 8.43944
R21182 dvss.n960 dvss 8.43944
R21183 dvss.n907 dvss 8.43944
R21184 dvss.n2037 dvss 8.43944
R21185 dvss.n1895 dvss 8.43944
R21186 dvss.n1780 dvss 8.43944
R21187 dvss.n6376 dvss 8.43944
R21188 dvss.n6325 dvss 8.43944
R21189 dvss.n6259 dvss 8.43944
R21190 dvss.n5556 dvss 8.43944
R21191 dvss.n5502 dvss 8.43944
R21192 dvss.n5252 dvss 8.43944
R21193 dvss.n5213 dvss 8.43944
R21194 dvss.n5174 dvss 8.43944
R21195 dvss.n5135 dvss 8.43944
R21196 dvss.t2147 dvss.t1203 8.42962
R21197 dvss.n2846 dvss.t573 8.42962
R21198 dvss.t1111 dvss.t2134 8.42962
R21199 dvss.t1112 dvss.t985 8.42962
R21200 dvss.t927 dvss.t875 8.42962
R21201 dvss dvss.t715 8.42962
R21202 dvss.t983 dvss.t1093 8.42962
R21203 dvss.t836 dvss.t32 8.42962
R21204 dvss.t834 dvss.t496 8.42962
R21205 dvss.t2228 dvss.t1321 8.42962
R21206 dvss.n302 dvss.n301 8.35606
R21207 dvss.n270 dvss.n253 8.35606
R21208 dvss.n2304 dvss.n1233 8.34157
R21209 dvss.n4115 dvss.n4112 8.2968
R21210 dvss.n3800 dvss.n3636 8.28285
R21211 dvss.n3964 dvss.n3963 8.28285
R21212 dvss.n3987 dvss.n3461 8.28285
R21213 dvss.n5602 dvss.t1535 8.25063
R21214 dvss.n408 dvss.n391 8.2416
R21215 dvss.n2545 dvss.n2415 8.23546
R21216 dvss.n2652 dvss.n2415 8.23546
R21217 dvss.n2652 dvss.n2651 8.23546
R21218 dvss.n2648 dvss.n2647 8.23546
R21219 dvss.n2647 dvss.n2646 8.23546
R21220 dvss.n2623 dvss.n2622 8.23546
R21221 dvss.n2622 dvss.n2621 8.23546
R21222 dvss.n2621 dvss.n2571 8.23546
R21223 dvss.n2617 dvss.n2616 8.23546
R21224 dvss.n2616 dvss.n2615 8.23546
R21225 dvss.n2969 dvss.n2920 8.23546
R21226 dvss.n2965 dvss.n2920 8.23546
R21227 dvss.n2987 dvss.n2986 8.23546
R21228 dvss.n2761 dvss.n2703 8.23546
R21229 dvss.n2762 dvss.n2761 8.23546
R21230 dvss.n2763 dvss.n2762 8.23546
R21231 dvss.n2767 dvss.n2766 8.23546
R21232 dvss.n2768 dvss.n2767 8.23546
R21233 dvss.n2772 dvss.n2771 8.23546
R21234 dvss.n2774 dvss.n2772 8.23546
R21235 dvss.n3405 dvss.n3404 8.23546
R21236 dvss.n3401 dvss.n3400 8.23546
R21237 dvss.n3400 dvss.n3399 8.23546
R21238 dvss.n3374 dvss.n3356 8.23546
R21239 dvss.n3374 dvss.n3373 8.23546
R21240 dvss.n3371 dvss.n3358 8.23546
R21241 dvss.n3367 dvss.n3358 8.23546
R21242 dvss.n3592 dvss.n3520 8.23546
R21243 dvss.n3593 dvss.n3592 8.23546
R21244 dvss.n3594 dvss.n3593 8.23546
R21245 dvss.n4356 dvss.n4328 8.23546
R21246 dvss.n4484 dvss.n4483 8.23546
R21247 dvss.n4483 dvss.n4482 8.23546
R21248 dvss.n4482 dvss.n2364 8.23546
R21249 dvss.n4478 dvss.n4477 8.23546
R21250 dvss.n4475 dvss.n2368 8.23546
R21251 dvss.n4471 dvss.n2368 8.23546
R21252 dvss.n4464 dvss.n4463 8.23546
R21253 dvss.n4463 dvss.n4462 8.23546
R21254 dvss.n4462 dvss.n2373 8.23546
R21255 dvss.n4458 dvss.n4457 8.23546
R21256 dvss.n4457 dvss.n4456 8.23546
R21257 dvss.n4453 dvss.n4452 8.23546
R21258 dvss.n4452 dvss.n2379 8.23546
R21259 dvss.n4748 dvss.n4538 8.23546
R21260 dvss.n4744 dvss.n4538 8.23546
R21261 dvss.n4742 dvss.n4741 8.23546
R21262 dvss.n4741 dvss.n4540 8.23546
R21263 dvss.n4877 dvss.n4876 8.23546
R21264 dvss.n4878 dvss.n4877 8.23546
R21265 dvss.n4878 dvss.n4861 8.23546
R21266 dvss.n4882 dvss.n4861 8.23546
R21267 dvss.n4883 dvss.n4882 8.23546
R21268 dvss.n4884 dvss.n4883 8.23546
R21269 dvss.n4888 dvss.n4887 8.23546
R21270 dvss.n4890 dvss.n4888 8.23546
R21271 dvss.n3056 dvss.n3053 8.05976
R21272 dvss.n3689 dvss.n3657 8.05976
R21273 dvss.n3832 dvss.n3829 8.05976
R21274 dvss.n3407 dvss.n3406 8.05644
R21275 dvss.n3588 dvss.n3587 8.05644
R21276 dvss.n3597 dvss.n3518 8.05644
R21277 dvss.n4654 dvss.n4653 8.05644
R21278 dvss.n301 dvss.n300 8.0005
R21279 dvss.n271 dvss.n270 8.0005
R21280 dvss.t128 dvss.n1678 7.99565
R21281 dvss.n2952 dvss.n2927 7.90638
R21282 dvss.n3737 dvss.n3734 7.90638
R21283 dvss.n3899 dvss.n3898 7.90638
R21284 dvss.n3852 dvss.n3849 7.90638
R21285 dvss.n3932 dvss.n3922 7.90638
R21286 dvss.n3945 dvss.n3943 7.90638
R21287 dvss.n3953 dvss.n3951 7.90638
R21288 dvss.n409 dvss.n408 7.89091
R21289 dvss.n2973 dvss.n2972 7.87742
R21290 dvss.n3401 dvss.n3343 7.87742
R21291 dvss.n4487 dvss.n2328 7.87742
R21292 dvss.n4639 dvss.n4620 7.87742
R21293 dvss.n4393 dvss.n4310 7.8005
R21294 dvss.n2483 dvss.n2482 7.73676
R21295 dvss.n2646 dvss.n2420 7.6984
R21296 dvss.n2623 dvss.n2569 7.6984
R21297 dvss.n2973 dvss.n2918 7.6984
R21298 dvss.n2756 dvss.n2703 7.6984
R21299 dvss.n3407 dvss.n3342 7.6984
R21300 dvss.n3367 dvss.n3366 7.6984
R21301 dvss.n4329 dvss.n4328 7.6984
R21302 dvss.n4488 dvss.n4487 7.6984
R21303 dvss.n4464 dvss.n2371 7.6984
R21304 dvss.n2380 dvss.n2379 7.6984
R21305 dvss.n4656 dvss.n4655 7.6984
R21306 dvss.n4639 dvss.n4638 7.6984
R21307 dvss.n4876 dvss.n4863 7.6984
R21308 dvss.n4890 dvss.n4889 7.6984
R21309 dvss.n4507 dvss.n4506 7.5961
R21310 dvss.n3111 dvss.n3110 7.52991
R21311 dvss.n2731 dvss.n2730 7.52991
R21312 dvss.n3677 dvss.n3676 7.52991
R21313 dvss.n3891 dvss.n3890 7.52991
R21314 dvss.n3889 dvss.n3888 7.52991
R21315 dvss.n4285 dvss.n4284 7.52991
R21316 dvss.n358 dvss.n341 7.5205
R21317 dvss.n4543 dvss.n4542 7.51938
R21318 dvss.n7050 dvss.n7049 7.49264
R21319 dvss.n4378 dvss.n4377 7.47915
R21320 dvss.n1763 dvss.n1762 7.37677
R21321 dvss.n5126 dvss.n5125 7.37677
R21322 dvss.n7046 dvss.n7000 7.3244
R21323 dvss.n6995 dvss.n6994 7.25358
R21324 dvss.n4312 dvss.n4311 7.23528
R21325 dvss.n4582 dvss.n4579 7.21177
R21326 dvss.n359 dvss.n358 7.2005
R21327 dvss.n6604 dvss.n6603 7.2005
R21328 dvss.n4631 dvss.n4623 7.15344
R21329 dvss.n4178 dvss.n4177 7.15344
R21330 dvss.n2986 dvss.n2913 7.15139
R21331 dvss.n2977 dvss.n2976 7.11268
R21332 dvss.n2987 dvss.n2871 7.11268
R21333 dvss.n4357 dvss.n4356 7.11268
R21334 dvss.n4788 dvss.n4492 7.11268
R21335 dvss.n6604 dvss.n336 7.0405
R21336 dvss.n4788 dvss.n4493 6.90655
R21337 dvss.n3394 dvss.n3393 6.88949
R21338 dvss.n3600 dvss.n3597 6.88949
R21339 dvss.n4653 dvss.n4614 6.88949
R21340 dvss.n4643 dvss.n4642 6.88949
R21341 dvss.n4750 dvss.n4749 6.84415
R21342 dvss.t766 dvss.n5586 6.83569
R21343 dvss.n4377 dvss.n4376 6.79884
R21344 dvss.n2952 dvss.n2951 6.77697
R21345 dvss.n3035 dvss.n2854 6.77697
R21346 dvss.n2837 dvss.n2836 6.77697
R21347 dvss.n3993 dvss.n3992 6.77697
R21348 dvss.n4725 dvss.n4724 6.77697
R21349 dvss.n4123 dvss.n4122 6.77697
R21350 dvss.n3064 dvss.n3060 6.75606
R21351 dvss.n3378 dvss.n3356 6.56535
R21352 dvss.n2573 dvss.n2571 6.44526
R21353 dvss.n2774 dvss.n2773 6.44526
R21354 dvss.n2375 dvss.n2373 6.44526
R21355 dvss.n3562 dvss.n3561 6.4005
R21356 dvss.n4599 dvss.n4595 6.4005
R21357 dvss.n5063 dvss.n5010 6.4005
R21358 dvss.n3173 dvss 6.4005
R21359 dvss.n6454 dvss 6.4005
R21360 dvss.n173 dvss 6.4005
R21361 dvss.n582 dvss 6.4005
R21362 dvss.n625 dvss 6.4005
R21363 dvss.n1106 dvss 6.4005
R21364 dvss.n936 dvss 6.4005
R21365 dvss.n1375 dvss 6.4005
R21366 dvss.n1946 dvss 6.4005
R21367 dvss.n1840 dvss 6.4005
R21368 dvss.n6956 dvss 6.4005
R21369 dvss.n91 dvss 6.4005
R21370 dvss.n5971 dvss 6.4005
R21371 dvss.n5940 dvss 6.4005
R21372 dvss.n820 dvss 6.4005
R21373 dvss.n5808 dvss 6.4005
R21374 dvss.n1341 dvss 6.4005
R21375 dvss.n1310 dvss 6.4005
R21376 dvss.n1279 dvss 6.4005
R21377 dvss.n2547 dvss.n2546 6.26623
R21378 dvss.n4384 dvss.n4317 6.26433
R21379 dvss.n2635 dvss.n2634 6.26433
R21380 dvss.n3417 dvss.n2681 6.26433
R21381 dvss.n3434 dvss.n3433 6.26433
R21382 dvss.n2750 dvss.n2748 6.26433
R21383 dvss.n2791 dvss.n2786 6.26433
R21384 dvss.n3573 dvss.n3572 6.26433
R21385 dvss.n4437 dvss.n4436 6.26433
R21386 dvss.n4380 dvss.n4317 6.26433
R21387 dvss.n4380 dvss.n4379 6.26433
R21388 dvss.n4691 dvss.n4690 6.26433
R21389 dvss.n4690 dvss.n4689 6.26433
R21390 dvss.n4672 dvss.n4671 6.26433
R21391 dvss.n5035 dvss.n5034 6.26433
R21392 dvss.n4135 dvss.n4132 6.26433
R21393 dvss.n4085 dvss.n4082 6.26433
R21394 dvss.n4187 dvss.n4186 6.26433
R21395 dvss.t1537 dvss.n5609 6.21431
R21396 dvss.n4772 dvss.n4771 6.02861
R21397 dvss.n4759 dvss.n4758 6.02861
R21398 dvss.n3798 dvss.n3796 6.02403
R21399 dvss.n2554 dvss.n2537 5.98311
R21400 dvss.n3101 dvss.n3100 5.98311
R21401 dvss.n4868 dvss.n4867 5.98311
R21402 dvss.n4992 dvss.n4897 5.98311
R21403 dvss.n4979 dvss.n4902 5.98311
R21404 dvss.n4966 dvss.n4907 5.98311
R21405 dvss.n4941 dvss.n4916 5.98311
R21406 dvss.n5028 dvss.n5024 5.98311
R21407 dvss.n4698 dvss.n4582 5.91354
R21408 dvss.n2965 dvss.n2964 5.90819
R21409 dvss.n2367 dvss.n2364 5.90819
R21410 dvss.n289 dvss.n288 5.90523
R21411 dvss.n259 dvss.n257 5.90523
R21412 dvss.n4829 dvss.n4828 5.88889
R21413 dvss.n4380 dvss.n4319 5.8885
R21414 dvss.n397 dvss.n395 5.87299
R21415 dvss.n2636 dvss.n2635 5.85582
R21416 dvss.n3418 dvss.n3417 5.85582
R21417 dvss.n2748 dvss.n2747 5.85582
R21418 dvss.n2786 dvss.n2785 5.85582
R21419 dvss.n3570 dvss.n3526 5.85582
R21420 dvss.n4438 dvss.n4437 5.85582
R21421 dvss.n4392 dvss.n4391 5.85582
R21422 dvss.n5035 dvss.n5021 5.85582
R21423 dvss.n4082 dvss.n4081 5.85582
R21424 dvss.n4557 dvss.n4554 5.84398
R21425 dvss.n4781 dvss.n4780 5.82248
R21426 dvss.n4823 dvss.n4822 5.7429
R21427 dvss.n5003 dvss.t523 5.7362
R21428 dvss.n3573 dvss.n3523 5.65809
R21429 dvss.n4669 dvss.n4606 5.65809
R21430 dvss.n347 dvss.n345 5.65757
R21431 dvss.n2547 dvss.n2544 5.63966
R21432 dvss.n2612 dvss.n2611 5.63966
R21433 dvss.n3588 dvss.n3586 5.63966
R21434 dvss.n1132 dvss.t1545 5.59293
R21435 dvss.n3571 dvss.n3570 5.58348
R21436 dvss.n2491 dvss.n2490 5.56058
R21437 dvss.n4314 dvss.n4313 5.51774
R21438 dvss.n4691 dvss.n4586 5.51539
R21439 dvss.n295 dvss.n284 5.51161
R21440 dvss.n268 dvss.n267 5.51161
R21441 dvss.n2903 dvss.n2901 5.48128
R21442 dvss.n3246 dvss 5.45235
R21443 dvss.n6465 dvss 5.45235
R21444 dvss.n6672 dvss 5.45235
R21445 dvss.n716 dvss 5.45235
R21446 dvss.n638 dvss 5.45235
R21447 dvss.n5635 dvss 5.45235
R21448 dvss.n5688 dvss 5.45235
R21449 dvss.n1386 dvss 5.45235
R21450 dvss.n1975 dvss 5.45235
R21451 dvss.n1843 dvss 5.45235
R21452 dvss.n6962 dvss 5.45235
R21453 dvss.n6778 dvss 5.45235
R21454 dvss.n6026 dvss 5.45235
R21455 dvss.n6076 dvss 5.45235
R21456 dvss.n5884 dvss 5.45235
R21457 dvss.n5807 dvss 5.45235
R21458 dvss.n2120 dvss 5.45235
R21459 dvss.n2175 dvss 5.45235
R21460 dvss.n2225 dvss 5.45235
R21461 dvss.n406 dvss.n405 5.43612
R21462 dvss.n7051 dvss.n7050 5.4358
R21463 dvss.n4391 dvss.n4390 5.31114
R21464 dvss.n2384 dvss.n2381 5.27109
R21465 dvss.n4401 dvss.n4302 5.27109
R21466 dvss.n2819 dvss.n2675 5.17497
R21467 dvss.n305 dvss.n304 5.15606
R21468 dvss.n276 dvss.n275 5.15606
R21469 dvss.n2457 dvss.n2455 5.13108
R21470 dvss.n2457 dvss.n2456 5.13108
R21471 dvss.n2610 dvss.n2578 5.13108
R21472 dvss.n2589 dvss.n2586 5.13108
R21473 dvss.n2589 dvss.n2587 5.13108
R21474 dvss.n2881 dvss.n2879 5.13108
R21475 dvss.n2881 dvss.n2880 5.13108
R21476 dvss.n3076 dvss.n3073 5.13108
R21477 dvss.n3076 dvss.n3074 5.13108
R21478 dvss.n2718 dvss.n2715 5.13108
R21479 dvss.n2718 dvss.n2717 5.13108
R21480 dvss.n3364 dvss.n3361 5.13108
R21481 dvss.n3364 dvss.n3362 5.13108
R21482 dvss.n3669 dvss.n3666 5.13108
R21483 dvss.n3669 dvss.n3668 5.13108
R21484 dvss.n3863 dvss.n3860 5.13108
R21485 dvss.n3863 dvss.n3861 5.13108
R21486 dvss.n3927 dvss.n3924 5.13108
R21487 dvss.n3927 dvss.n3926 5.13108
R21488 dvss.n3539 dvss.n3537 5.13108
R21489 dvss.n3539 dvss.n3538 5.13108
R21490 dvss.n4340 dvss.n4337 5.13108
R21491 dvss.n4340 dvss.n4339 5.13108
R21492 dvss.n2337 dvss.n2335 5.13108
R21493 dvss.n2337 dvss.n2336 5.13108
R21494 dvss.n4502 dvss.n4500 5.13108
R21495 dvss.n4502 dvss.n4501 5.13108
R21496 dvss.n4628 dvss.n4625 5.13108
R21497 dvss.n4628 dvss.n4627 5.13108
R21498 dvss.n4061 dvss.n4059 5.13108
R21499 dvss.n4061 dvss.n4060 5.13108
R21500 dvss.n4221 dvss.n4218 5.13108
R21501 dvss.n4221 dvss.n4219 5.13108
R21502 dvss.n1696 dvss.n1695 5.11678
R21503 dvss.n1693 dvss.n1692 5.11678
R21504 dvss.n414 dvss.n413 5.08543
R21505 dvss.n2166 dvss.n2165 4.96991
R21506 dvss.n883 dvss.n882 4.96991
R21507 dvss.n5815 dvss.n5814 4.96991
R21508 dvss.n5899 dvss.n5898 4.96991
R21509 dvss.n1403 dvss.n1402 4.96991
R21510 dvss.n1452 dvss.n1451 4.96991
R21511 dvss.n985 dvss.n984 4.96991
R21512 dvss.n802 dvss.n801 4.96991
R21513 dvss.n356 dvss.n355 4.9605
R21514 dvss.n3818 dvss.n3634 4.89462
R21515 dvss dvss.n6580 4.88722
R21516 dvss.n457 dvss 4.88201
R21517 dvss dvss.n242 4.8781
R21518 dvss.n6632 dvss 4.8729
R21519 dvss.n2896 dvss.n2895 4.85762
R21520 dvss.n3381 dvss.n3355 4.85762
R21521 dvss.n3580 dvss.n3579 4.85762
R21522 dvss.n4663 dvss.n4609 4.85762
R21523 dvss.n4684 dvss.n4683 4.85762
R21524 dvss.n2552 dvss.n2539 4.85567
R21525 dvss.n2766 dvss.n2701 4.83407
R21526 dvss.n6995 dvss.n6989 4.80519
R21527 dvss.n3100 dvss.n3099 4.8005
R21528 dvss.n4719 dvss.n4718 4.8005
R21529 dvss.n4698 dvss.n4697 4.8005
R21530 dvss.n4868 dvss.n4866 4.8005
R21531 dvss.n4992 dvss.n4991 4.8005
R21532 dvss.n4979 dvss.n4978 4.8005
R21533 dvss.n4966 dvss.n4965 4.8005
R21534 dvss.n4941 dvss.n4940 4.8005
R21535 dvss.n5028 dvss.n5027 4.8005
R21536 dvss.n2465 dvss.n2464 4.67352
R21537 dvss.n2466 dvss.n2465 4.67352
R21538 dvss.n2466 dvss.n2452 4.67352
R21539 dvss.n2470 dvss.n2452 4.67352
R21540 dvss.n2471 dvss.n2470 4.67352
R21541 dvss.n2472 dvss.n2471 4.67352
R21542 dvss.n2476 dvss.n2475 4.67352
R21543 dvss.n2478 dvss.n2476 4.67352
R21544 dvss.n2510 dvss.n2509 4.67352
R21545 dvss.n2511 dvss.n2510 4.67352
R21546 dvss.n2511 dvss.n2437 4.67352
R21547 dvss.n2515 dvss.n2437 4.67352
R21548 dvss.n2516 dvss.n2515 4.67352
R21549 dvss.n2517 dvss.n2516 4.67352
R21550 dvss.n2521 dvss.n2520 4.67352
R21551 dvss.n2523 dvss.n2521 4.67352
R21552 dvss.n2606 dvss.n2605 4.67352
R21553 dvss.n2605 dvss.n2604 4.67352
R21554 dvss.n2604 dvss.n2581 4.67352
R21555 dvss.n2600 dvss.n2581 4.67352
R21556 dvss.n2600 dvss.n2599 4.67352
R21557 dvss.n2599 dvss.n2598 4.67352
R21558 dvss.n2595 dvss.n2594 4.67352
R21559 dvss.n2594 dvss.n2593 4.67352
R21560 dvss.n2982 dvss.n2981 4.67352
R21561 dvss.n2981 dvss.n2980 4.67352
R21562 dvss.n2907 dvss.n2906 4.67352
R21563 dvss.n2909 dvss.n2907 4.67352
R21564 dvss.n3093 dvss.n3092 4.67352
R21565 dvss.n3092 dvss.n3091 4.67352
R21566 dvss.n3091 dvss.n3068 4.67352
R21567 dvss.n3087 dvss.n3068 4.67352
R21568 dvss.n3087 dvss.n3086 4.67352
R21569 dvss.n3086 dvss.n3085 4.67352
R21570 dvss.n3082 dvss.n3081 4.67352
R21571 dvss.n3081 dvss.n3080 4.67352
R21572 dvss.n2345 dvss.n2344 4.67352
R21573 dvss.n2346 dvss.n2345 4.67352
R21574 dvss.n2346 dvss.n2332 4.67352
R21575 dvss.n2350 dvss.n2332 4.67352
R21576 dvss.n2351 dvss.n2350 4.67352
R21577 dvss.n2353 dvss.n2351 4.67352
R21578 dvss.n2357 dvss.n2330 4.67352
R21579 dvss.n2358 dvss.n2357 4.67352
R21580 dvss.n4369 dvss.n4368 4.67352
R21581 dvss.n4368 dvss.n4322 4.67352
R21582 dvss.n4364 dvss.n4322 4.67352
R21583 dvss.n4362 dvss.n4361 4.67352
R21584 dvss.n4361 dvss.n4324 4.67352
R21585 dvss.n4777 dvss.n4776 4.67352
R21586 dvss.n4776 dvss.n4775 4.67352
R21587 dvss.n4768 dvss.n4767 4.67352
R21588 dvss.n4765 dvss.n4532 4.67352
R21589 dvss.n4761 dvss.n4532 4.67352
R21590 dvss.n4755 dvss.n4754 4.67352
R21591 dvss.n4754 dvss.n4753 4.67352
R21592 dvss.t1682 dvss.t677 4.66076
R21593 dvss.n3396 dvss.n3346 4.65505
R21594 dvss.n364 dvss.n363 4.6405
R21595 dvss.n4087 dvss.n4051 4.62124
R21596 dvss.n4371 dvss.n4320 4.55559
R21597 dvss.n4518 dvss.n4517 4.55559
R21598 dvss.n2780 dvss.n2778 4.51815
R21599 dvss.n3780 dvss.n3777 4.51815
R21600 dvss.n4092 dvss.n4091 4.51815
R21601 dvss.n4162 dvss.n4161 4.51815
R21602 dvss.n4284 dvss.n4017 4.51815
R21603 dvss.n4274 dvss.n4273 4.51815
R21604 dvss.n2662 dvss.n2409 4.51401
R21605 dvss.n2414 dvss.n2413 4.51401
R21606 dvss.n3017 dvss.n3015 4.51401
R21607 dvss.n3027 dvss.n3026 4.51401
R21608 dvss.n3444 dvss.n2668 4.51401
R21609 dvss.n2673 dvss.n2672 4.51401
R21610 dvss.n3792 dvss.n3790 4.51401
R21611 dvss.n3811 dvss.n3810 4.51401
R21612 dvss.n3478 dvss.n3475 4.51401
R21613 dvss.n3452 dvss.n3449 4.51401
R21614 dvss.n2404 dvss.n2403 4.51401
R21615 dvss.n4409 dvss.n4408 4.51401
R21616 dvss.n4712 dvss.n4711 4.51401
R21617 dvss.n4706 dvss.n4705 4.51401
R21618 dvss.n4926 dvss.n4924 4.51401
R21619 dvss.n1217 dvss.n1213 4.51401
R21620 dvss.n4170 dvss.n4169 4.51401
R21621 dvss.n4290 dvss.n4289 4.51401
R21622 dvss.n2661 dvss.n2660 4.5005
R21623 dvss.n2659 dvss.n2658 4.5005
R21624 dvss.n2655 dvss.n2654 4.5005
R21625 dvss.n3019 dvss.n3018 4.5005
R21626 dvss.n3022 dvss.n3021 4.5005
R21627 dvss.n2860 dvss.n2859 4.5005
R21628 dvss.n3443 dvss.n3442 4.5005
R21629 dvss.n3441 dvss.n3440 4.5005
R21630 dvss.n3437 dvss.n3436 4.5005
R21631 dvss.n3794 dvss.n3793 4.5005
R21632 dvss.n3806 dvss.n3805 4.5005
R21633 dvss.n3641 dvss.n3638 4.5005
R21634 dvss.n3481 dvss.n3480 4.5005
R21635 dvss.n3477 dvss.n3451 4.5005
R21636 dvss.n4002 dvss.n4001 4.5005
R21637 dvss.n4416 dvss.n4415 4.5005
R21638 dvss.n2405 dvss.n2402 4.5005
R21639 dvss.n4296 dvss.n4294 4.5005
R21640 dvss.n4569 dvss.n4560 4.5005
R21641 dvss.n4571 dvss.n4570 4.5005
R21642 dvss.n4572 dvss.n4563 4.5005
R21643 dvss.n4929 dvss.n4928 4.5005
R21644 dvss.n4925 dvss.n1215 4.5005
R21645 dvss.n5095 dvss.n5094 4.5005
R21646 dvss.n4168 dvss.n4167 4.5005
R21647 dvss.n4166 dvss.n4165 4.5005
R21648 dvss.n4155 dvss.n4010 4.5005
R21649 dvss.n2464 dvss.n2454 4.36875
R21650 dvss.n2478 dvss.n2477 4.36875
R21651 dvss.n2509 dvss.n2439 4.36875
R21652 dvss.n2523 dvss.n2522 4.36875
R21653 dvss.n2606 dvss.n2579 4.36875
R21654 dvss.n2593 dvss.n2585 4.36875
R21655 dvss.n2980 dvss.n2917 4.36875
R21656 dvss.n2909 dvss.n2908 4.36875
R21657 dvss.n3093 dvss.n3067 4.36875
R21658 dvss.n3080 dvss.n3072 4.36875
R21659 dvss.n2344 dvss.n2334 4.36875
R21660 dvss.n2359 dvss.n2358 4.36875
R21661 dvss.n4370 dvss.n4369 4.36875
R21662 dvss.n4521 dvss.n4519 4.36875
R21663 dvss.n4521 dvss.n4520 4.36875
R21664 dvss.n4775 dvss.n4529 4.36875
R21665 dvss.n4768 dvss.n4530 4.36875
R21666 dvss.n4761 dvss.n4760 4.36875
R21667 dvss.n4753 dvss.n4537 4.36875
R21668 dvss.n7041 dvss.n7017 4.3437
R21669 dvss.n4470 dvss.n4469 4.297
R21670 dvss.n4385 dvss.n4384 4.28986
R21671 dvss.n5034 dvss.n5033 4.28986
R21672 dvss.n4085 dvss.n4084 4.28986
R21673 dvss.n3606 dvss.n3515 4.2869
R21674 dvss.n5088 dvss.n1220 4.26717
R21675 dvss.n5041 dvss.n5018 4.26717
R21676 dvss.n7047 dvss.n7046 4.25273
R21677 dvss.n3770 dvss.n3769 4.14168
R21678 dvss.n3484 dvss.n3483 4.14168
R21679 dvss.n4333 dvss.n4331 4.14168
R21680 dvss.n2651 dvss.n2416 4.11798
R21681 dvss.n2612 dvss.n2576 4.11798
R21682 dvss.n2971 dvss.n2970 4.11798
R21683 dvss.n2970 dvss.n2969 4.11798
R21684 dvss.n2768 dvss.n2698 4.11798
R21685 dvss.n2771 dvss.n2698 4.11798
R21686 dvss.n3396 dvss.n3395 4.11798
R21687 dvss.n3395 dvss.n3394 4.11798
R21688 dvss.n3373 dvss.n3372 4.11798
R21689 dvss.n3372 dvss.n3371 4.11798
R21690 dvss.n4477 dvss.n4476 4.11798
R21691 dvss.n4476 dvss.n4475 4.11798
R21692 dvss.n4453 dvss.n2378 4.11798
R21693 dvss.n4744 dvss.n4743 4.11798
R21694 dvss.n4743 dvss.n4742 4.11798
R21695 dvss.n4884 dvss.n4859 4.11798
R21696 dvss.n4887 dvss.n4859 4.11798
R21697 dvss.n2543 dvss.n2542 4.09013
R21698 dvss.n4375 dvss.n4374 4.09013
R21699 dvss.n4131 dvss.n4130 4.08561
R21700 dvss.n2725 dvss.n2722 4.07323
R21701 dvss.n2722 dvss.n2714 4.07323
R21702 dvss.n5033 dvss.n5032 4.07323
R21703 dvss.n4084 dvss.n4051 4.07323
R21704 dvss.n2495 dvss.n2494 3.96548
R21705 dvss.n2496 dvss.n2495 3.96548
R21706 dvss.n2500 dvss.n2499 3.96548
R21707 dvss.n2888 dvss.n2877 3.96548
R21708 dvss.n3604 dvss.n3516 3.96548
R21709 dvss.n3605 dvss.n3604 3.96548
R21710 dvss.n4512 dvss.n4511 3.96548
R21711 dvss.n4513 dvss.n4512 3.96548
R21712 dvss.n4649 dvss.n4648 3.96548
R21713 dvss.n4648 dvss.n4647 3.96548
R21714 dvss.n4647 dvss.n4617 3.96548
R21715 dvss.n4670 dvss.n4669 3.94944
R21716 dvss.n2576 dvss.n2575 3.93896
R21717 dvss.n2378 dvss.n2377 3.93896
R21718 dvss.n2389 dvss.n2386 3.90237
R21719 dvss.n2823 dvss.n2822 3.76521
R21720 dvss.n4262 dvss.n4261 3.76521
R21721 dvss.n2487 dvss.n2485 3.7575
R21722 dvss.n4784 dvss.n4525 3.7575
R21723 dvss.n7032 dvss.n7031 3.72777
R21724 dvss.n2494 dvss.n2444 3.7069
R21725 dvss.n2502 dvss.n2440 3.7069
R21726 dvss.n2888 dvss.n2887 3.7069
R21727 dvss.n3390 dvss.n3348 3.7069
R21728 dvss.n3390 dvss.n3389 3.7069
R21729 dvss.n4511 dvss.n4498 3.7069
R21730 dvss.n4649 dvss.n4616 3.7069
R21731 dvss.n3279 dvss.n3278 3.68864
R21732 dvss.n6451 dvss.n34 3.68864
R21733 dvss.n6668 dvss.n74 3.68864
R21734 dvss.n712 dvss.n709 3.68864
R21735 dvss.n758 dvss.n537 3.68864
R21736 dvss.n5631 dvss.n798 3.68864
R21737 dvss.n5684 dvss.n5681 3.68864
R21738 dvss.n1408 dvss.n1360 3.68864
R21739 dvss.n1971 dvss.n1448 3.68864
R21740 dvss.n1863 dvss.n1862 3.68864
R21741 dvss.n6421 dvss.n6420 3.68864
R21742 dvss.n6558 dvss.n6348 3.68864
R21743 dvss.n6300 dvss.n6299 3.68864
R21744 dvss.n6230 dvss.n6229 3.68864
R21745 dvss.n5535 dvss.n5534 3.68864
R21746 dvss.n5278 dvss.n5277 3.68864
R21747 dvss.n5239 dvss.n5238 3.68864
R21748 dvss.n5200 dvss.n5199 3.68864
R21749 dvss.n5161 dvss.n5160 3.68864
R21750 dvss.n2892 dvss.n2877 3.68605
R21751 dvss.n4187 dvss.n4141 3.6771
R21752 dvss.n4111 dvss.n4037 3.63493
R21753 dvss.t523 dvss.t1682 3.58531
R21754 dvss.n3399 dvss.n3346 3.58092
R21755 dvss.n3578 dvss.n3577 3.50735
R21756 dvss.n4685 dvss.n4590 3.50735
R21757 dvss.n4665 dvss.n4607 3.50735
R21758 dvss.n4689 dvss.n4588 3.49783
R21759 dvss.n2725 dvss.n2724 3.47876
R21760 dvss.n2165 dvss 3.46403
R21761 dvss.n882 dvss 3.46403
R21762 dvss.n5814 dvss 3.46403
R21763 dvss.n5898 dvss 3.46403
R21764 dvss.n1402 dvss 3.46403
R21765 dvss.n1451 dvss 3.46403
R21766 dvss.n984 dvss 3.46403
R21767 dvss.n801 dvss 3.46403
R21768 dvss.n2413 dvss.n2407 3.43925
R21769 dvss.n2663 dvss.n2662 3.43925
R21770 dvss.n3026 dvss.n3025 3.43925
R21771 dvss.n3017 dvss.n3016 3.43925
R21772 dvss.n2672 dvss.n2666 3.43925
R21773 dvss.n3445 dvss.n3444 3.43925
R21774 dvss.n3810 dvss.n3809 3.43925
R21775 dvss.n3792 dvss.n3791 3.43925
R21776 dvss.n4005 dvss.n3449 3.43925
R21777 dvss.n3478 dvss.n3448 3.43925
R21778 dvss.n4410 dvss.n4409 3.43925
R21779 dvss.n4412 dvss.n2404 3.43925
R21780 dvss.n4707 dvss.n4706 3.43925
R21781 dvss.n4711 dvss.n4710 3.43925
R21782 dvss.n5098 dvss.n1213 3.43925
R21783 dvss.n4926 dvss.n1212 3.43925
R21784 dvss.n2410 dvss.n2408 3.4105
R21785 dvss.n2657 dvss.n2656 3.4105
R21786 dvss.n2862 dvss.n2861 3.4105
R21787 dvss.n3024 dvss.n3023 3.4105
R21788 dvss.n2669 dvss.n2667 3.4105
R21789 dvss.n3439 dvss.n3438 3.4105
R21790 dvss.n3640 dvss.n3639 3.4105
R21791 dvss.n3808 dvss.n3807 3.4105
R21792 dvss.n3479 dvss.n3450 3.4105
R21793 dvss.n4004 dvss.n4003 3.4105
R21794 dvss.n4414 dvss.n4413 3.4105
R21795 dvss.n4293 dvss.n2406 3.4105
R21796 dvss.n4709 dvss.n4561 3.4105
R21797 dvss.n4708 dvss.n4562 3.4105
R21798 dvss.n4927 dvss.n1214 3.4105
R21799 dvss.n5097 dvss.n5096 3.4105
R21800 dvss.n4292 dvss.n4291 3.4105
R21801 dvss.n4292 dvss.n4008 3.4105
R21802 dvss.n4291 dvss.n4290 3.4105
R21803 dvss.n4169 dvss.n4008 3.4105
R21804 dvss.n4154 dvss.n4153 3.4105
R21805 dvss.n4164 dvss.n4009 3.4105
R21806 dvss.n2763 dvss.n2701 3.4019
R21807 dvss.n4471 dvss.n4470 3.4019
R21808 dvss.n2529 dvss.n2528 3.38874
R21809 dvss.n3552 dvss.n3533 3.38874
R21810 dvss.n5010 dvss.n5007 3.38874
R21811 dvss.n3622 dvss.n3620 3.37632
R21812 dvss.n1760 dvss 3.25474
R21813 dvss.n5123 dvss 3.25474
R21814 dvss.n5102 dvss.n5101 3.20904
R21815 dvss.n3582 dvss.n3522 3.2005
R21816 dvss.n4682 dvss.n4681 3.2005
R21817 dvss.n4664 dvss.n4608 3.2005
R21818 dvss.n2634 dvss.n2427 3.13241
R21819 dvss.n2683 dvss.n2681 3.13241
R21820 dvss.n3433 dvss.n2676 3.13241
R21821 dvss.n2750 dvss.n2749 3.13241
R21822 dvss.n2791 dvss.n2790 3.13241
R21823 dvss.n4436 dvss.n2390 3.13241
R21824 dvss.n4314 dvss.n4311 3.13241
R21825 dvss.n4135 dvss.n4134 3.13241
R21826 dvss.n4186 dvss.n4185 3.13241
R21827 dvss.n3387 dvss.n3350 3.09945
R21828 dvss.n2458 dvss.n2457 3.05586
R21829 dvss.n2882 dvss.n2881 3.05586
R21830 dvss.n2718 dvss.n2716 3.05586
R21831 dvss.n3669 dvss.n3667 3.05586
R21832 dvss.n3540 dvss.n3539 3.05586
R21833 dvss.n2338 dvss.n2337 3.05586
R21834 dvss.n4503 dvss.n4502 3.05586
R21835 dvss.n4062 dvss.n4061 3.05586
R21836 dvss.n2589 dvss.n2588 3.04861
R21837 dvss.n2610 dvss.n2577 3.04861
R21838 dvss.n3076 dvss.n3075 3.04861
R21839 dvss.n3364 dvss.n3363 3.04861
R21840 dvss.n3863 dvss.n3862 3.04861
R21841 dvss.n3927 dvss.n3925 3.04861
R21842 dvss.n4340 dvss.n4338 3.04861
R21843 dvss.n4628 dvss.n4626 3.04861
R21844 dvss.n5032 dvss.n5023 3.04861
R21845 dvss.n4221 dvss.n4220 3.04861
R21846 dvss.n2549 dvss.n2543 3.04861
R21847 dvss.n2722 dvss.n2721 3.04861
R21848 dvss.n4374 dvss.n4373 3.04861
R21849 dvss.n2487 dvss.n2486 3.01483
R21850 dvss.n4784 dvss.n4783 3.01483
R21851 dvss.n4815 dvss.n1236 3.01226
R21852 dvss.n4378 dvss.n4375 2.99624
R21853 dvss.n4604 dvss.n4603 2.99624
R21854 dvss.n6580 dvss.n6579 2.94679
R21855 dvss dvss.n6 2.94111
R21856 dvss.n4513 dvss.n4496 2.88804
R21857 dvss.n6640 dvss.n6639 2.87444
R21858 dvss.n2544 dvss.n2543 2.86855
R21859 dvss.n4374 dvss.n4320 2.86855
R21860 dvss.t1277 dvss.t40 2.86835
R21861 dvss.n2419 dvss.n2416 2.86484
R21862 dvss.n4672 dvss.n4604 2.86007
R21863 dvss.n2611 dvss.n2610 2.8567
R21864 dvss.n3247 dvss.n3246 2.84494
R21865 dvss.n6466 dvss.n6465 2.84494
R21866 dvss.n6672 dvss.n6671 2.84494
R21867 dvss.n716 dvss.n715 2.84494
R21868 dvss.n639 dvss.n638 2.84494
R21869 dvss.n5635 dvss.n5634 2.84494
R21870 dvss.n5688 dvss.n5687 2.84494
R21871 dvss.n1387 dvss.n1386 2.84494
R21872 dvss.n1975 dvss.n1974 2.84494
R21873 dvss.n1843 dvss.n1842 2.84494
R21874 dvss.n6962 dvss.n6961 2.84494
R21875 dvss.n6779 dvss.n6778 2.84494
R21876 dvss.n6026 dvss.n6025 2.84494
R21877 dvss.n6076 dvss.n6075 2.84494
R21878 dvss.n5885 dvss.n5884 2.84494
R21879 dvss.n5807 dvss.n5806 2.84494
R21880 dvss.n2120 dvss.n2119 2.84494
R21881 dvss.n2175 dvss.n2174 2.84494
R21882 dvss.n2225 dvss.n2224 2.84494
R21883 dvss.n5100 dvss.n1210 2.80662
R21884 dvss.n4496 dvss.n4495 2.79323
R21885 dvss.n2554 dvss.n2553 2.78311
R21886 dvss.n2428 dvss.n2427 2.7239
R21887 dvss.n2677 dvss.n2676 2.7239
R21888 dvss.n2749 dvss.n2704 2.7239
R21889 dvss.n2391 dvss.n2390 2.7239
R21890 dvss.n4134 dvss.n4133 2.7239
R21891 dvss.n4185 dvss.n4184 2.7239
R21892 dvss.n2166 dvss 2.71109
R21893 dvss.n883 dvss 2.71109
R21894 dvss.n5815 dvss 2.71109
R21895 dvss.n5899 dvss 2.71109
R21896 dvss.n1403 dvss 2.71109
R21897 dvss.n1452 dvss 2.71109
R21898 dvss.n985 dvss 2.71109
R21899 dvss.n802 dvss 2.71109
R21900 dvss.n293 dvss.n292 2.66717
R21901 dvss.n261 dvss.n256 2.66717
R21902 dvss.n2945 dvss.n2932 2.63579
R21903 dvss.n3044 dvss.n2852 2.63579
R21904 dvss.n3747 dvss.n3744 2.63579
R21905 dvss.n3683 dvss.n3682 2.63579
R21906 dvss.n3834 dvss.n3630 2.63579
R21907 dvss.n3872 dvss.n3871 2.63579
R21908 dvss.n3956 dvss.n3954 2.63579
R21909 dvss.n3545 dvss.n3544 2.63579
R21910 dvss.n3553 dvss.n3552 2.63579
R21911 dvss.n4427 dvss.n4426 2.63579
R21912 dvss.n4100 dvss.n4041 2.63579
R21913 dvss.n4273 dvss.n4272 2.63579
R21914 dvss.n4662 dvss.n4661 2.63064
R21915 dvss.n399 dvss.n394 2.63064
R21916 dvss.n3247 dvss 2.60791
R21917 dvss.n6466 dvss 2.60791
R21918 dvss.n6671 dvss 2.60791
R21919 dvss.n715 dvss 2.60791
R21920 dvss.n639 dvss 2.60791
R21921 dvss.n5634 dvss 2.60791
R21922 dvss.n5687 dvss 2.60791
R21923 dvss.n1387 dvss 2.60791
R21924 dvss.n1974 dvss 2.60791
R21925 dvss.n1842 dvss 2.60791
R21926 dvss.n6961 dvss 2.60791
R21927 dvss.n6779 dvss 2.60791
R21928 dvss.n6025 dvss 2.60791
R21929 dvss.n6075 dvss 2.60791
R21930 dvss.n5885 dvss 2.60791
R21931 dvss.n5806 dvss 2.60791
R21932 dvss.n2119 dvss 2.60791
R21933 dvss.n2174 dvss 2.60791
R21934 dvss.n2224 dvss 2.60791
R21935 dvss.n2894 dvss.n2893 2.55412
R21936 dvss.n3383 dvss.n3351 2.55412
R21937 dvss.n5003 dvss.t2121 2.50987
R21938 dvss.n2327 dvss.n2326 2.50679
R21939 dvss.n3514 dvss.n3512 2.50485
R21940 dvss.n1616 dvss 2.49542
R21941 dvss.n1710 dvss 2.49542
R21942 dvss.n2272 dvss 2.49542
R21943 dvss.n2279 dvss 2.49542
R21944 dvss.n2323 dvss.n1233 2.46192
R21945 dvss.n2685 dvss.n2684 2.45156
R21946 dvss.n426 dvss.n380 2.43615
R21947 dvss.n349 dvss.n344 2.4005
R21948 dvss.n3620 dvss.n3506 2.39171
R21949 dvss.n2542 dvss.n2540 2.38348
R21950 dvss.n2472 dvss.n2450 2.33701
R21951 dvss.n2475 dvss.n2450 2.33701
R21952 dvss.n2517 dvss.n2435 2.33701
R21953 dvss.n2520 dvss.n2435 2.33701
R21954 dvss.n2598 dvss.n2583 2.33701
R21955 dvss.n2595 dvss.n2583 2.33701
R21956 dvss.n2982 dvss.n2916 2.33701
R21957 dvss.n2906 dvss.n2873 2.33701
R21958 dvss.n3085 dvss.n3070 2.33701
R21959 dvss.n3082 dvss.n3070 2.33701
R21960 dvss.n2353 dvss.n2352 2.33701
R21961 dvss.n2352 dvss.n2330 2.33701
R21962 dvss.n4364 dvss.n4363 2.33701
R21963 dvss.n4363 dvss.n4362 2.33701
R21964 dvss.n4325 dvss.n4324 2.33701
R21965 dvss.n4777 dvss.n4528 2.33701
R21966 dvss.n4767 dvss.n4766 2.33701
R21967 dvss.n4766 dvss.n4765 2.33701
R21968 dvss.n4755 dvss.n4536 2.33701
R21969 dvss.n2898 dvss.n2876 2.33067
R21970 dvss.n3382 dvss.n3354 2.33067
R21971 dvss.n4478 dvss.n2367 2.32777
R21972 dvss.n2790 dvss.n2789 2.31539
R21973 dvss.n4671 dvss.n4670 2.31539
R21974 dvss.n332 dvss.n281 2.31161
R21975 dvss.n323 dvss.n310 2.31161
R21976 dvss.n6613 dvss.n250 2.31161
R21977 dvss.n6622 dvss.n246 2.31161
R21978 dvss.n438 dvss.n388 2.27995
R21979 dvss.n447 dvss.n384 2.27995
R21980 dvss.n3676 dvss.n3675 2.25932
R21981 dvss.n4447 dvss.n2381 2.25932
R21982 dvss.n4302 dvss.n4301 2.25932
R21983 dvss.n4159 dvss.n4157 2.25932
R21984 dvss.n4516 dvss.n4515 2.25312
R21985 dvss.n7050 dvss 2.21678
R21986 dvss.n4141 dvss.n4140 2.17922
R21987 dvss.n424 dvss.n422 2.17238
R21988 dvss.n3113 dvss.n3056 2.13383
R21989 dvss.n3835 dvss.n3832 2.13383
R21990 dvss.n4517 dvss.n4516 2.09505
R21991 dvss.n368 dvss.n367 2.0805
R21992 dvss.n6598 dvss.n371 2.0805
R21993 dvss.n2501 dvss.n2500 2.06919
R21994 dvss.n4108 dvss.n4037 2.03468
R21995 dvss.n2916 dvss.n2915 2.03225
R21996 dvss.n2902 dvss.n2873 2.03225
R21997 dvss.n4326 dvss.n4325 2.03225
R21998 dvss.n4528 dvss.n4526 2.03225
R21999 dvss.n4536 dvss.n4534 2.03225
R22000 dvss.n4702 dvss.n4701 2.01789
R22001 dvss.n4686 dvss.n4588 1.99413
R22002 dvss.n2496 dvss.n2442 1.98299
R22003 dvss.n2499 dvss.n2442 1.98299
R22004 dvss.n3598 dvss.n3516 1.98299
R22005 dvss.n3606 dvss.n3605 1.98299
R22006 dvss.n4618 dvss.n4617 1.98299
R22007 dvss.n4394 dvss.n4308 1.97497
R22008 dvss.n2546 dvss.n2545 1.96973
R22009 dvss.n2897 dvss.n2874 1.91571
R22010 dvss.n3380 dvss.n3379 1.91571
R22011 dvss.n2502 dvss.n2501 1.8968
R22012 dvss.n3693 dvss.n3692 1.8968
R22013 dvss.n4116 dvss.n4115 1.8968
R22014 dvss.n5100 dvss 1.89242
R22015 dvss.n2955 dvss.n2927 1.88285
R22016 dvss.n2799 dvss.n2686 1.88285
R22017 dvss.n3738 dvss.n3737 1.88285
R22018 dvss.n3788 dvss.n3642 1.88285
R22019 dvss.n3900 dvss.n3899 1.88285
R22020 dvss.n3878 dvss.n3852 1.88285
R22021 dvss.n3946 dvss.n3945 1.88285
R22022 dvss.n3954 dvss.n3953 1.88285
R22023 dvss.n4550 dvss.n4547 1.88285
R22024 dvss.n2757 dvss.n2755 1.88081
R22025 dvss.n6633 dvss.n6632 1.87648
R22026 dvss.n3231 dvss 1.84457
R22027 dvss dvss.n3230 1.84457
R22028 dvss.n3230 dvss 1.84457
R22029 dvss.n6937 dvss 1.84457
R22030 dvss dvss.n6936 1.84457
R22031 dvss.n6936 dvss 1.84457
R22032 dvss.n6683 dvss 1.84457
R22033 dvss dvss.n6682 1.84457
R22034 dvss.n6682 dvss 1.84457
R22035 dvss.n727 dvss 1.84457
R22036 dvss dvss.n726 1.84457
R22037 dvss.n726 dvss 1.84457
R22038 dvss.n6196 dvss 1.84457
R22039 dvss dvss.n6195 1.84457
R22040 dvss.n6195 dvss 1.84457
R22041 dvss.n1099 dvss 1.84457
R22042 dvss dvss.n1098 1.84457
R22043 dvss.n1098 dvss 1.84457
R22044 dvss.n5699 dvss 1.84457
R22045 dvss dvss.n5698 1.84457
R22046 dvss.n5698 dvss 1.84457
R22047 dvss.n2093 dvss 1.84457
R22048 dvss dvss.n2092 1.84457
R22049 dvss.n2092 dvss 1.84457
R22050 dvss.n1940 dvss 1.84457
R22051 dvss.n1923 dvss 1.84457
R22052 dvss.n1923 dvss 1.84457
R22053 dvss.n1828 dvss 1.84457
R22054 dvss.n1808 dvss 1.84457
R22055 dvss.n1808 dvss 1.84457
R22056 dvss.n6826 dvss 1.84457
R22057 dvss dvss.n6825 1.84457
R22058 dvss.n6825 dvss 1.84457
R22059 dvss.n6764 dvss 1.84457
R22060 dvss dvss.n6763 1.84457
R22061 dvss.n6763 dvss 1.84457
R22062 dvss.n6035 dvss 1.84457
R22063 dvss dvss.n6034 1.84457
R22064 dvss.n6034 dvss 1.84457
R22065 dvss.n6085 dvss 1.84457
R22066 dvss dvss.n6084 1.84457
R22067 dvss.n6084 dvss 1.84457
R22068 dvss.n5870 dvss 1.84457
R22069 dvss dvss.n5869 1.84457
R22070 dvss.n5869 dvss 1.84457
R22071 dvss.n5792 dvss 1.84457
R22072 dvss.n5778 dvss 1.84457
R22073 dvss.n5778 dvss 1.84457
R22074 dvss.n2129 dvss 1.84457
R22075 dvss dvss.n2128 1.84457
R22076 dvss.n2128 dvss 1.84457
R22077 dvss.n2184 dvss 1.84457
R22078 dvss dvss.n2183 1.84457
R22079 dvss.n2183 dvss 1.84457
R22080 dvss.n2234 dvss 1.84457
R22081 dvss dvss.n2233 1.84457
R22082 dvss.n2233 dvss 1.84457
R22083 dvss.n3102 dvss.n3064 1.82737
R22084 dvss.n2617 dvss.n2573 1.79071
R22085 dvss.n2964 dvss.n2963 1.79071
R22086 dvss.n4458 dvss.n2375 1.79071
R22087 dvss.n4132 dvss.n4131 1.77071
R22088 dvss.n4595 dvss.n4592 1.75392
R22089 dvss.n3599 dvss.n3598 1.72441
R22090 dvss.n3607 dvss.n3606 1.72441
R22091 dvss.n4619 dvss.n4618 1.72441
R22092 dvss.n7037 dvss.n7023 1.72109
R22093 dvss.n7024 dvss.n7017 1.72109
R22094 dvss.n5099 dvss.n1212 1.69188
R22095 dvss.n5099 dvss.n5098 1.69188
R22096 dvss.n4707 dvss.n1211 1.69188
R22097 dvss.n4710 dvss.n1211 1.69188
R22098 dvss.n4411 dvss.n4410 1.69188
R22099 dvss.n4412 dvss.n4411 1.69188
R22100 dvss.n4006 dvss.n3448 1.69188
R22101 dvss.n4006 dvss.n4005 1.69188
R22102 dvss.n3809 dvss.n3447 1.69188
R22103 dvss.n3791 dvss.n3447 1.69188
R22104 dvss.n3446 dvss.n2666 1.69188
R22105 dvss.n3446 dvss.n3445 1.69188
R22106 dvss.n3025 dvss.n2665 1.69188
R22107 dvss.n3016 dvss.n2665 1.69188
R22108 dvss.n2664 dvss.n2407 1.69188
R22109 dvss.n2664 dvss.n2663 1.69188
R22110 dvss.n4292 dvss.n4007 1.69188
R22111 dvss.n2553 dvss.n2552 1.6005
R22112 dvss.n6989 dvss.n6 1.5923
R22113 dvss.n437 dvss.n415 1.57858
R22114 dvss.n3120 dvss.n3119 1.50638
R22115 dvss.n3110 dvss.n3057 1.50638
R22116 dvss.n2809 dvss.n2806 1.50638
R22117 dvss.n2737 dvss.n2708 1.50638
R22118 dvss.n3671 dvss.n3670 1.50638
R22119 dvss.n3963 dvss.n3962 1.50638
R22120 dvss.n3972 dvss.n3971 1.50638
R22121 dvss.n4076 dvss.n4054 1.50638
R22122 dvss.n4174 dvss.n4173 1.50638
R22123 dvss.n6633 dvss.n241 1.50538
R22124 dvss.n2637 dvss.n2426 1.48166
R22125 dvss dvss.n241 1.47804
R22126 dvss dvss.n6633 1.47268
R22127 dvss.n322 dvss.n311 1.42272
R22128 dvss.n6624 dvss.n6623 1.42272
R22129 dvss.n449 dvss.n448 1.40324
R22130 dvss.n4379 dvss.n4378 1.3622
R22131 dvss.n7006 dvss.n6997 1.35909
R22132 dvss.n3214 dvss.n3190 1.34003
R22133 dvss.n3216 dvss.n3181 1.34003
R22134 dvss.n3229 dvss.n3181 1.34003
R22135 dvss.n6919 dvss.n54 1.34003
R22136 dvss.n6921 dvss.n37 1.34003
R22137 dvss.n6935 dvss.n37 1.34003
R22138 dvss.n6693 dvss.n151 1.34003
R22139 dvss.n6691 dvss.n153 1.34003
R22140 dvss.n6681 dvss.n153 1.34003
R22141 dvss.n737 dvss.n563 1.34003
R22142 dvss.n735 dvss.n565 1.34003
R22143 dvss.n725 dvss.n565 1.34003
R22144 dvss.n6178 dvss.n778 1.34003
R22145 dvss.n6180 dvss.n761 1.34003
R22146 dvss.n6194 dvss.n761 1.34003
R22147 dvss.n1086 dvss.n1084 1.34003
R22148 dvss.n1095 dvss.n1093 1.34003
R22149 dvss.n1097 dvss.n1095 1.34003
R22150 dvss.n5709 dvss.n917 1.34003
R22151 dvss.n5707 dvss.n919 1.34003
R22152 dvss.n5697 dvss.n919 1.34003
R22153 dvss.n2075 dvss.n1428 1.34003
R22154 dvss.n2077 dvss.n1411 1.34003
R22155 dvss.n2091 dvss.n1411 1.34003
R22156 dvss.n1909 dvss.n1908 1.34003
R22157 dvss.n1922 dvss.n1920 1.34003
R22158 dvss.n1924 dvss.n1922 1.34003
R22159 dvss.n1787 dvss.n1786 1.34003
R22160 dvss.n1807 dvss.n1805 1.34003
R22161 dvss.n1809 dvss.n1807 1.34003
R22162 dvss.n6843 dvss.n6842 1.34003
R22163 dvss.n6835 dvss.n6834 1.34003
R22164 dvss.n6834 dvss.n6833 1.34003
R22165 dvss.n6747 dvss.n108 1.34003
R22166 dvss.n6749 dvss.n99 1.34003
R22167 dvss.n6762 dvss.n99 1.34003
R22168 dvss.n6052 dvss.n6051 1.34003
R22169 dvss.n6044 dvss.n6043 1.34003
R22170 dvss.n6043 dvss.n6042 1.34003
R22171 dvss.n6102 dvss.n6101 1.34003
R22172 dvss.n6094 dvss.n6093 1.34003
R22173 dvss.n6093 dvss.n6092 1.34003
R22174 dvss.n5853 dvss.n837 1.34003
R22175 dvss.n5855 dvss.n828 1.34003
R22176 dvss.n5868 dvss.n828 1.34003
R22177 dvss.n5762 dvss.n5761 1.34003
R22178 dvss.n5777 dvss.n5775 1.34003
R22179 dvss.n5779 dvss.n5777 1.34003
R22180 dvss.n2146 dvss.n2145 1.34003
R22181 dvss.n2138 dvss.n2137 1.34003
R22182 dvss.n2137 dvss.n2136 1.34003
R22183 dvss.n2201 dvss.n2200 1.34003
R22184 dvss.n2193 dvss.n2192 1.34003
R22185 dvss.n2192 dvss.n2191 1.34003
R22186 dvss.n2251 dvss.n2250 1.34003
R22187 dvss.n2243 dvss.n2242 1.34003
R22188 dvss.n2242 dvss.n2241 1.34003
R22189 dvss.n2542 dvss.n2541 1.3283
R22190 dvss.n2725 dvss.n2712 1.32281
R22191 dvss.n2714 dvss.n2713 1.32281
R22192 dvss.n6597 dvss.n372 1.2805
R22193 dvss.n6588 dvss.n376 1.2805
R22194 dvss.n4678 dvss.n4677 1.27173
R22195 dvss.n2484 dvss.n2483 1.26739
R22196 dvss.n2648 dvss.n2419 1.25365
R22197 dvss.n2773 dvss.n2696 1.25365
R22198 dvss.n3608 dvss.n3512 1.25033
R22199 dvss.n4508 dvss.n4507 1.25033
R22200 dvss.n4931 dvss.n4923 1.23559
R22201 dvss.n5049 dvss.n5048 1.23559
R22202 dvss.n6989 dvss 1.23235
R22203 dvss.n2886 dvss.n2885 1.20723
R22204 dvss.n1210 dvss.n1209 1.20499
R22205 dvss.n3099 dvss.n3098 1.18311
R22206 dvss.n4718 dvss.n4717 1.18311
R22207 dvss.n4697 dvss.n4696 1.18311
R22208 dvss.n4866 dvss.n4865 1.18311
R22209 dvss.n4991 dvss.n4990 1.18311
R22210 dvss.n4978 dvss.n4977 1.18311
R22211 dvss.n4965 dvss.n4964 1.18311
R22212 dvss.n4940 dvss.n4939 1.18311
R22213 dvss.n5027 dvss.n5026 1.18311
R22214 dvss.n457 dvss.n380 1.16554
R22215 dvss.n4389 dvss.n4311 1.15795
R22216 dvss.n3582 dvss.n3581 1.14023
R22217 dvss.n4681 dvss.n4591 1.14023
R22218 dvss.n4662 dvss.n4608 1.14023
R22219 dvss.n3971 dvss.n3970 1.12991
R22220 dvss.n3545 dvss.n3534 1.12991
R22221 dvss.n4724 dvss.n4723 1.12991
R22222 dvss.n4575 dvss.n4574 1.12991
R22223 dvss.n4827 dvss.n1235 1.12991
R22224 dvss.n351 dvss.n345 1.12105
R22225 dvss.n7047 dvss.n6997 1.09648
R22226 dvss.n426 dvss.n425 1.09487
R22227 dvss.n401 dvss.n395 1.05227
R22228 dvss.n4439 dvss.n2389 1.0468
R22229 dvss.n290 dvss.n289 1.04213
R22230 dvss.n263 dvss.n257 1.04213
R22231 dvss.n1238 dvss.n1236 0.970649
R22232 dvss.n1237 dvss.n1235 0.970649
R22233 dvss.n2296 dvss.n1237 0.970649
R22234 dvss.n6589 dvss.n375 0.9605
R22235 dvss.n4376 dvss.n4375 0.956517
R22236 dvss.n4390 dvss.n4389 0.953691
R22237 dvss.n5033 dvss.n5022 0.952566
R22238 dvss.n4084 dvss.n4083 0.952566
R22239 dvss.n380 dvss.n242 0.934094
R22240 dvss.n4814 dvss.n4813 0.907477
R22241 dvss.n4813 dvss.n4812 0.907477
R22242 dvss.n4826 dvss.n4825 0.907477
R22243 dvss.n4051 dvss.n4050 0.899674
R22244 dvss.n4516 dvss.n4496 0.892621
R22245 dvss.n427 dvss.n426 0.886661
R22246 dvss.n4595 dvss.n4591 0.877212
R22247 dvss dvss.n3214 0.856314
R22248 dvss.n3216 dvss.n3215 0.856314
R22249 dvss dvss.n3229 0.856314
R22250 dvss dvss.n6919 0.856314
R22251 dvss.n6921 dvss.n6920 0.856314
R22252 dvss dvss.n6935 0.856314
R22253 dvss.n6693 dvss 0.856314
R22254 dvss.n6692 dvss.n6691 0.856314
R22255 dvss dvss.n6681 0.856314
R22256 dvss.n737 dvss 0.856314
R22257 dvss.n736 dvss.n735 0.856314
R22258 dvss dvss.n725 0.856314
R22259 dvss dvss.n6178 0.856314
R22260 dvss.n6180 dvss.n6179 0.856314
R22261 dvss dvss.n6194 0.856314
R22262 dvss dvss.n1086 0.856314
R22263 dvss.n1093 dvss.n1087 0.856314
R22264 dvss dvss.n1097 0.856314
R22265 dvss.n5709 dvss 0.856314
R22266 dvss.n5708 dvss.n5707 0.856314
R22267 dvss dvss.n5697 0.856314
R22268 dvss dvss.n2075 0.856314
R22269 dvss.n2077 dvss.n2076 0.856314
R22270 dvss dvss.n2091 0.856314
R22271 dvss.n1909 dvss 0.856314
R22272 dvss.n1920 dvss.n1478 0.856314
R22273 dvss.n1924 dvss 0.856314
R22274 dvss.n1786 dvss 0.856314
R22275 dvss.n1805 dvss.n1544 0.856314
R22276 dvss.n1809 dvss 0.856314
R22277 dvss.n6842 dvss 0.856314
R22278 dvss.n6835 dvss.n6803 0.856314
R22279 dvss.n6833 dvss 0.856314
R22280 dvss dvss.n6747 0.856314
R22281 dvss.n6749 dvss.n6748 0.856314
R22282 dvss dvss.n6762 0.856314
R22283 dvss.n6051 dvss 0.856314
R22284 dvss.n6044 dvss.n5961 0.856314
R22285 dvss.n6042 dvss 0.856314
R22286 dvss.n6101 dvss 0.856314
R22287 dvss.n6094 dvss.n5914 0.856314
R22288 dvss.n6092 dvss 0.856314
R22289 dvss dvss.n5853 0.856314
R22290 dvss.n5855 dvss.n5854 0.856314
R22291 dvss dvss.n5868 0.856314
R22292 dvss.n5762 dvss 0.856314
R22293 dvss.n5775 dvss.n865 0.856314
R22294 dvss.n5779 dvss 0.856314
R22295 dvss.n2145 dvss 0.856314
R22296 dvss.n2138 dvss.n1331 0.856314
R22297 dvss.n2136 dvss 0.856314
R22298 dvss.n2200 dvss 0.856314
R22299 dvss.n2193 dvss.n1300 0.856314
R22300 dvss.n2191 dvss 0.856314
R22301 dvss.n2250 dvss 0.856314
R22302 dvss.n2243 dvss.n1269 0.856314
R22303 dvss.n2241 dvss 0.856314
R22304 dvss.n3577 dvss.n3522 0.833377
R22305 dvss.n4682 dvss.n4590 0.833377
R22306 dvss.n4665 dvss.n4664 0.833377
R22307 dvss.n2898 dvss.n2897 0.830425
R22308 dvss.n3380 dvss.n3354 0.830425
R22309 dvss.n7052 dvss.n7051 0.827044
R22310 dvss.n6632 dvss.n242 0.808117
R22311 dvss.n3387 dvss.n3386 0.798505
R22312 dvss.n2664 dvss.n1210 0.792753
R22313 dvss.n1701 dvss.n5 0.789073
R22314 dvss.n425 dvss.n418 0.7755
R22315 dvss.n430 dvss.n429 0.7755
R22316 dvss.n2939 dvss.n2938 0.753441
R22317 dvss.n3031 dvss.n2856 0.753441
R22318 dvss.n2838 dvss.n2837 0.753441
R22319 dvss.n3998 dvss.n3997 0.753441
R22320 dvss.n4732 dvss.n4550 0.753441
R22321 dvss.n4253 dvss.n4252 0.753441
R22322 dvss.n4240 dvss.n4207 0.753441
R22323 dvss.n4231 dvss.n4230 0.753441
R22324 dvss.n2486 dvss.n2445 0.743162
R22325 dvss.n4783 dvss.n4782 0.743162
R22326 dvss.n3053 dvss.n3051 0.711611
R22327 dvss.n3105 dvss.n3060 0.711611
R22328 dvss.n3829 dvss.n3828 0.711611
R22329 dvss.n4112 dvss.n4111 0.711611
R22330 dvss.n333 dvss.n279 0.711611
R22331 dvss.n6612 dvss.n277 0.711611
R22332 dvss.n428 dvss.n427 0.705857
R22333 dvss.n3623 dvss.n3622 0.703797
R22334 dvss.n4599 dvss.n4598 0.696152
R22335 dvss.n6580 dvss.n457 0.692883
R22336 dvss.n3434 dvss.n2675 0.681351
R22337 dvss.n3572 dvss.n3571 0.681351
R22338 dvss.n3623 dvss.n3618 0.633467
R22339 dvss.n6992 dvss.t657 0.627052
R22340 dvss.n6990 dvss.t654 0.627052
R22341 dvss.n7026 dvss.t287 0.627052
R22342 dvss.n2893 dvss.n2876 0.606984
R22343 dvss.n3383 dvss.n3382 0.606984
R22344 dvss.n6991 dvss.n6990 0.5805
R22345 dvss.n6993 dvss.n6992 0.5805
R22346 dvss.n7030 dvss.n7029 0.5805
R22347 dvss.n7029 dvss.n7028 0.5805
R22348 dvss.n7028 dvss.n7027 0.5805
R22349 dvss.n7027 dvss.n7026 0.5805
R22350 dvss.n4818 dvss.n4817 0.561438
R22351 dvss.n7035 dvss.n6996 0.54848
R22352 dvss dvss.n6 0.543548
R22353 dvss.n2626 dvss.n2569 0.537563
R22354 dvss.n2976 dvss.n2918 0.537563
R22355 dvss.n2963 dvss.n2962 0.537563
R22356 dvss.n2757 dvss.n2756 0.537563
R22357 dvss.n2777 dvss.n2696 0.537563
R22358 dvss.n3342 dvss.n3340 0.537563
R22359 dvss.n3366 dvss.n3365 0.537563
R22360 dvss.n4352 dvss.n4329 0.537563
R22361 dvss.n4469 dvss.n4468 0.537563
R22362 dvss.n4467 dvss.n2371 0.537563
R22363 dvss.n4448 dvss.n2380 0.537563
R22364 dvss.n4737 dvss.n4543 0.537563
R22365 dvss.n4657 dvss.n4656 0.537563
R22366 dvss.n4873 dvss.n4863 0.537563
R22367 dvss.n4889 dvss.n4857 0.537563
R22368 dvss.n328 dvss.n327 0.533833
R22369 dvss.n6618 dvss.n6617 0.533833
R22370 dvss.n429 dvss.n422 0.529518
R22371 dvss.n3578 dvss.n3523 0.526527
R22372 dvss.n4686 dvss.n4685 0.526527
R22373 dvss.n4607 dvss.n4606 0.526527
R22374 dvss.n443 dvss.n442 0.526527
R22375 dvss.n4849 dvss.n4829 0.514786
R22376 dvss.n6603 dvss.n6602 0.4805
R22377 dvss.n3689 dvss.n3688 0.474574
R22378 dvss.n3692 dvss.n3657 0.474574
R22379 dvss.n4921 dvss.n4918 0.449623
R22380 dvss.n5056 dvss.n5055 0.449623
R22381 dvss.n4489 dvss.n4488 0.448052
R22382 dvss.n2302 dvss.n2301 0.429848
R22383 dvss.n4844 dvss.n4843 0.429848
R22384 dvss.n4831 dvss.n4830 0.429848
R22385 dvss.n4835 dvss.n4834 0.429848
R22386 dvss.n4839 dvss.n4838 0.429848
R22387 dvss.n2310 dvss.n2309 0.429848
R22388 dvss.n2316 dvss.n2315 0.429848
R22389 dvss.n2319 dvss.n2318 0.429848
R22390 dvss.n7010 dvss.n7009 0.427268
R22391 dvss.n4599 dvss.n4596 0.427167
R22392 dvss.n2556 dvss.n2537 0.417891
R22393 dvss.n3102 dvss.n3101 0.417891
R22394 dvss.n3098 dvss.n3097 0.417891
R22395 dvss.n4722 dvss.n4554 0.417891
R22396 dvss.n4717 dvss.n4716 0.417891
R22397 dvss.n4701 dvss.n4580 0.417891
R22398 dvss.n4696 dvss.n4695 0.417891
R22399 dvss.n4867 dvss.n4864 0.417891
R22400 dvss.n4995 dvss.n4897 0.417891
R22401 dvss.n4990 dvss.n4989 0.417891
R22402 dvss.n4982 dvss.n4902 0.417891
R22403 dvss.n4977 dvss.n4976 0.417891
R22404 dvss.n4969 dvss.n4907 0.417891
R22405 dvss.n4964 dvss.n4963 0.417891
R22406 dvss.n4944 dvss.n4916 0.417891
R22407 dvss.n4939 dvss.n4938 0.417891
R22408 dvss.n5031 dvss.n5024 0.417891
R22409 dvss.n2637 dvss.n2636 0.409011
R22410 dvss.n2631 dvss.n2428 0.409011
R22411 dvss.n3419 dvss.n3418 0.409011
R22412 dvss.n3413 dvss.n2685 0.409011
R22413 dvss.n2820 dvss.n2819 0.409011
R22414 dvss.n3430 dvss.n2677 0.409011
R22415 dvss.n2747 dvss.n2746 0.409011
R22416 dvss.n2753 dvss.n2704 0.409011
R22417 dvss.n2785 dvss.n2784 0.409011
R22418 dvss.n2789 dvss.n2788 0.409011
R22419 dvss.n2788 dvss.n2690 0.409011
R22420 dvss.n3567 dvss.n3526 0.409011
R22421 dvss.n4439 dvss.n4438 0.409011
R22422 dvss.n4694 dvss.n4583 0.409011
R22423 dvss.n4603 dvss.n4600 0.409011
R22424 dvss.n5021 dvss.n5019 0.409011
R22425 dvss.n4130 dvss.n4129 0.409011
R22426 dvss.n4133 dvss.n4025 0.409011
R22427 dvss.n4081 dvss.n4080 0.409011
R22428 dvss.n4140 dvss.n4026 0.409011
R22429 dvss.n4184 dvss.n4183 0.409011
R22430 dvss.n2894 dvss.n2892 0.383542
R22431 dvss.n3386 dvss.n3351 0.383542
R22432 dvss.n2824 dvss.n2823 0.376971
R22433 dvss.n2797 dvss.n2796 0.376971
R22434 dvss.n4568 dvss.n4567 0.376971
R22435 dvss.n5068 dvss.n5067 0.376971
R22436 dvss.n4175 dvss.n4174 0.376971
R22437 dvss.n2643 dvss.n2421 0.358542
R22438 dvss.n2972 dvss.n2971 0.358542
R22439 dvss.n3404 dvss.n3343 0.358542
R22440 dvss.n4484 dvss.n2328 0.358542
R22441 dvss.n4642 dvss.n4620 0.358542
R22442 dvss.n4638 dvss.n4637 0.358542
R22443 dvss.n4586 dvss.n4583 0.340926
R22444 dvss.n7013 dvss.n7000 0.312562
R22445 dvss.n2461 dvss.n2454 0.305262
R22446 dvss.n2477 dvss.n2447 0.305262
R22447 dvss.n2506 dvss.n2439 0.305262
R22448 dvss.n2522 dvss.n2433 0.305262
R22449 dvss.n2609 dvss.n2579 0.305262
R22450 dvss.n2590 dvss.n2585 0.305262
R22451 dvss.n2915 dvss.n2913 0.305262
R22452 dvss.n2977 dvss.n2917 0.305262
R22453 dvss.n2903 dvss.n2902 0.305262
R22454 dvss.n2908 dvss.n2871 0.305262
R22455 dvss.n3067 dvss.n3065 0.305262
R22456 dvss.n3077 dvss.n3072 0.305262
R22457 dvss.n2341 dvss.n2334 0.305262
R22458 dvss.n2360 dvss.n2359 0.305262
R22459 dvss.n4371 dvss.n4370 0.305262
R22460 dvss.n4357 dvss.n4326 0.305262
R22461 dvss.n4519 dvss.n4518 0.305262
R22462 dvss.n4520 dvss.n4492 0.305262
R22463 dvss.n4780 dvss.n4526 0.305262
R22464 dvss.n4772 dvss.n4529 0.305262
R22465 dvss.n4771 dvss.n4530 0.305262
R22466 dvss.n4760 dvss.n4759 0.305262
R22467 dvss.n4758 dvss.n4534 0.305262
R22468 dvss.n4750 dvss.n4537 0.305262
R22469 dvss.n7008 dvss.n7007 0.299742
R22470 dvss.n4515 dvss.n4514 0.298074
R22471 dvss.n6994 dvss.n6991 0.279444
R22472 dvss.n2684 dvss.n2683 0.27284
R22473 dvss.n4433 dvss.n2392 0.27284
R22474 dvss.n4749 dvss.n4748 0.269031
R22475 dvss.n6994 dvss.n6993 0.268206
R22476 dvss.n4678 dvss.n4592 0.263514
R22477 dvss.n4661 dvss.n4660 0.263514
R22478 dvss.n2485 dvss.n2484 0.262616
R22479 dvss.n2490 dvss.n2445 0.262616
R22480 dvss.n4525 dvss.n4493 0.262616
R22481 dvss.n4782 dvss.n4781 0.262616
R22482 dvss.n2491 dvss.n2444 0.259086
R22483 dvss.n2505 dvss.n2440 0.259086
R22484 dvss.n2887 dvss.n2886 0.259086
R22485 dvss.n3393 dvss.n3348 0.259086
R22486 dvss.n3389 dvss.n3388 0.259086
R22487 dvss.n3600 dvss.n3599 0.259086
R22488 dvss.n3608 dvss.n3607 0.259086
R22489 dvss.n4508 dvss.n4498 0.259086
R22490 dvss.n4616 dvss.n4614 0.259086
R22491 dvss.n4643 dvss.n4619 0.259086
R22492 dvss.n7014 dvss.n7013 0.254288
R22493 dvss.n425 dvss.n424 0.2505
R22494 dvss.n4849 dvss.n4848 0.246929
R22495 dvss.n5023 dvss.n5020 0.239726
R22496 dvss.n4660 dvss.n4611 0.230065
R22497 dvss.n2588 dvss 0.217246
R22498 dvss.n3075 dvss 0.217246
R22499 dvss.n2312 dvss.n2311 0.215174
R22500 dvss.n2311 dvss.n2310 0.215174
R22501 dvss.n2317 dvss.n2316 0.215174
R22502 dvss.n2318 dvss.n2317 0.215174
R22503 dvss.n2320 dvss.n2319 0.215174
R22504 dvss.n2321 dvss.n2320 0.215174
R22505 dvss.n2323 dvss.n2322 0.213463
R22506 dvss.n4818 dvss.n2303 0.209875
R22507 dvss.n2746 dvss.n2706 0.207909
R22508 dvss.n4394 dvss.n4393 0.204755
R22509 dvss.n4393 dvss.n4392 0.204755
R22510 dvss.n7051 dvss.n5 0.201543
R22511 dvss.n4515 dvss 0.199635
R22512 dvss.n4848 dvss.n4842 0.193435
R22513 dvss.n5101 dvss.n5 0.192025
R22514 dvss.n2901 dvss.n2874 0.192021
R22515 dvss.n3379 dvss.n3378 0.192021
R22516 dvss.n2303 dvss.n2302 0.188611
R22517 dvss.n4087 dvss.n4086 0.180304
R22518 dvss.n3862 dvss 0.17983
R22519 dvss.n4220 dvss 0.17983
R22520 dvss dvss.n2549 0.17983
R22521 dvss.n2721 dvss 0.17983
R22522 dvss.n2421 dvss.n2420 0.179521
R22523 dvss.n2615 dvss.n2575 0.179521
R22524 dvss.n3406 dvss.n3405 0.179521
R22525 dvss.n3587 dvss.n3520 0.179521
R22526 dvss.n3594 dvss.n3518 0.179521
R22527 dvss.n4456 dvss.n2377 0.179521
R22528 dvss.n4542 dvss.n4540 0.179521
R22529 dvss.n4655 dvss.n4654 0.179521
R22530 dvss.n4637 dvss.n4636 0.179521
R22531 dvss.n2577 dvss 0.179485
R22532 dvss.n3363 dvss 0.179485
R22533 dvss.n3925 dvss 0.179485
R22534 dvss.n4373 dvss 0.179485
R22535 dvss.n4338 dvss 0.179485
R22536 dvss.n4626 dvss 0.179485
R22537 dvss.n7038 dvss.n7032 0.179346
R22538 dvss.n7036 dvss.n7035 0.179346
R22539 dvss.n7046 dvss.n7045 0.179346
R22540 dvss.n7015 dvss.n7014 0.179346
R22541 dvss.n429 dvss.n428 0.176839
R22542 dvss.n7000 dvss.n6999 0.174082
R22543 dvss dvss.n2458 0.172576
R22544 dvss dvss.n2882 0.172576
R22545 dvss.n2716 dvss 0.172576
R22546 dvss.n3667 dvss 0.172576
R22547 dvss dvss.n3540 0.172576
R22548 dvss dvss.n2338 0.172576
R22549 dvss dvss.n4503 0.172576
R22550 dvss dvss.n4062 0.172576
R22551 dvss.n2665 dvss.n2664 0.1603
R22552 dvss.n3446 dvss.n2665 0.1603
R22553 dvss.n3447 dvss.n3446 0.1603
R22554 dvss.n4006 dvss.n3447 0.1603
R22555 dvss.n4292 dvss.n4006 0.1603
R22556 dvss.n4411 dvss.n4292 0.1603
R22557 dvss.n4411 dvss.n1211 0.1603
R22558 dvss.n5099 dvss.n1211 0.1603
R22559 dvss.n4846 dvss.n4844 0.152674
R22560 dvss.n4833 dvss.n4831 0.152674
R22561 dvss.n4834 dvss.n4833 0.152674
R22562 dvss.n4837 dvss.n4835 0.152674
R22563 dvss.n4838 dvss.n4837 0.152674
R22564 dvss.n4841 dvss.n4839 0.152674
R22565 dvss.n4842 dvss.n4841 0.152674
R22566 dvss.n4847 dvss.n4846 0.152674
R22567 dvss.n7014 dvss.n7010 0.145702
R22568 dvss dvss.n2577 0.14207
R22569 dvss.n2588 dvss 0.14207
R22570 dvss.n3075 dvss 0.14207
R22571 dvss.n3363 dvss 0.14207
R22572 dvss.n3925 dvss 0.14207
R22573 dvss.n4338 dvss 0.14207
R22574 dvss.n4626 dvss 0.14207
R22575 dvss.n4373 dvss 0.14207
R22576 dvss.n2549 dvss 0.141725
R22577 dvss.n2721 dvss 0.141725
R22578 dvss.n3862 dvss 0.141725
R22579 dvss dvss.n5023 0.141725
R22580 dvss.n4220 dvss 0.141725
R22581 dvss.n4719 dvss.n4557 0.13963
R22582 dvss.n2392 dvss.n2391 0.13667
R22583 dvss.n4080 dvss.n4053 0.13667
R22584 dvss.n2322 dvss.n2321 0.130935
R22585 dvss.n7035 dvss.n7034 0.129288
R22586 dvss dvss.n4087 0.120408
R22587 dvss.n2463 dvss.n2462 0.120292
R22588 dvss.n2463 dvss.n2453 0.120292
R22589 dvss.n2467 dvss.n2453 0.120292
R22590 dvss.n2468 dvss.n2467 0.120292
R22591 dvss.n2469 dvss.n2468 0.120292
R22592 dvss.n2469 dvss.n2451 0.120292
R22593 dvss.n2473 dvss.n2451 0.120292
R22594 dvss.n2474 dvss.n2473 0.120292
R22595 dvss.n2474 dvss.n2449 0.120292
R22596 dvss.n2479 dvss.n2449 0.120292
R22597 dvss.n2480 dvss.n2479 0.120292
R22598 dvss.n2488 dvss.n2446 0.120292
R22599 dvss.n2489 dvss.n2488 0.120292
R22600 dvss.n2493 dvss.n2492 0.120292
R22601 dvss.n2493 dvss.n2443 0.120292
R22602 dvss.n2497 dvss.n2443 0.120292
R22603 dvss.n2498 dvss.n2497 0.120292
R22604 dvss.n2498 dvss.n2441 0.120292
R22605 dvss.n2503 dvss.n2441 0.120292
R22606 dvss.n2504 dvss.n2503 0.120292
R22607 dvss.n2508 dvss.n2507 0.120292
R22608 dvss.n2508 dvss.n2438 0.120292
R22609 dvss.n2512 dvss.n2438 0.120292
R22610 dvss.n2513 dvss.n2512 0.120292
R22611 dvss.n2514 dvss.n2513 0.120292
R22612 dvss.n2514 dvss.n2436 0.120292
R22613 dvss.n2518 dvss.n2436 0.120292
R22614 dvss.n2519 dvss.n2518 0.120292
R22615 dvss.n2519 dvss.n2434 0.120292
R22616 dvss.n2524 dvss.n2434 0.120292
R22617 dvss.n2525 dvss.n2524 0.120292
R22618 dvss.n2530 dvss.n2430 0.120292
R22619 dvss.n2531 dvss.n2530 0.120292
R22620 dvss.n2560 dvss.n2534 0.120292
R22621 dvss.n2536 dvss.n2534 0.120292
R22622 dvss dvss.n2555 0.120292
R22623 dvss.n2650 dvss.n2649 0.120292
R22624 dvss.n2649 dvss.n2417 0.120292
R22625 dvss.n2645 dvss.n2644 0.120292
R22626 dvss.n2640 dvss.n2639 0.120292
R22627 dvss.n2638 dvss.n2424 0.120292
R22628 dvss.n2633 dvss.n2424 0.120292
R22629 dvss.n2633 dvss.n2632 0.120292
R22630 dvss.n2625 dvss.n2624 0.120292
R22631 dvss.n2624 dvss.n2570 0.120292
R22632 dvss.n2620 dvss.n2570 0.120292
R22633 dvss.n2620 dvss.n2619 0.120292
R22634 dvss.n2619 dvss.n2618 0.120292
R22635 dvss.n2618 dvss.n2572 0.120292
R22636 dvss.n2614 dvss.n2572 0.120292
R22637 dvss.n2614 dvss.n2613 0.120292
R22638 dvss.n2608 dvss.n2607 0.120292
R22639 dvss.n2607 dvss.n2580 0.120292
R22640 dvss.n2603 dvss.n2580 0.120292
R22641 dvss.n2603 dvss.n2602 0.120292
R22642 dvss.n2602 dvss.n2601 0.120292
R22643 dvss.n2601 dvss.n2582 0.120292
R22644 dvss.n2597 dvss.n2582 0.120292
R22645 dvss.n2597 dvss.n2596 0.120292
R22646 dvss.n2596 dvss.n2584 0.120292
R22647 dvss.n2592 dvss.n2584 0.120292
R22648 dvss.n2592 dvss.n2591 0.120292
R22649 dvss.n2889 dvss.n2878 0.120292
R22650 dvss.n2890 dvss.n2889 0.120292
R22651 dvss.n2891 dvss.n2890 0.120292
R22652 dvss.n2891 dvss.n2875 0.120292
R22653 dvss.n2899 dvss.n2875 0.120292
R22654 dvss.n2900 dvss.n2899 0.120292
R22655 dvss.n2905 dvss.n2904 0.120292
R22656 dvss.n2905 dvss.n2872 0.120292
R22657 dvss.n2910 dvss.n2872 0.120292
R22658 dvss.n2911 dvss.n2910 0.120292
R22659 dvss.n2984 dvss.n2983 0.120292
R22660 dvss.n2983 dvss.n2914 0.120292
R22661 dvss.n2979 dvss.n2914 0.120292
R22662 dvss.n2979 dvss.n2978 0.120292
R22663 dvss.n2975 dvss.n2974 0.120292
R22664 dvss.n2974 dvss.n2919 0.120292
R22665 dvss.n2968 dvss.n2919 0.120292
R22666 dvss.n2968 dvss.n2967 0.120292
R22667 dvss.n2967 dvss.n2966 0.120292
R22668 dvss.n2966 dvss.n2921 0.120292
R22669 dvss.n2960 dvss.n2959 0.120292
R22670 dvss.n2959 dvss.n2924 0.120292
R22671 dvss.n2954 dvss.n2924 0.120292
R22672 dvss.n2954 dvss.n2953 0.120292
R22673 dvss.n2953 dvss.n2928 0.120292
R22674 dvss.n2948 dvss.n2928 0.120292
R22675 dvss.n2948 dvss.n2947 0.120292
R22676 dvss.n2947 dvss.n2946 0.120292
R22677 dvss.n2946 dvss.n2930 0.120292
R22678 dvss.n2942 dvss.n2930 0.120292
R22679 dvss.n2942 dvss.n2941 0.120292
R22680 dvss.n2941 dvss.n2940 0.120292
R22681 dvss.n2940 dvss.n2934 0.120292
R22682 dvss.n2993 dvss.n2868 0.120292
R22683 dvss.n2998 dvss.n2868 0.120292
R22684 dvss.n2999 dvss.n2998 0.120292
R22685 dvss.n3000 dvss.n2999 0.120292
R22686 dvss.n3000 dvss.n2866 0.120292
R22687 dvss.n3006 dvss.n2866 0.120292
R22688 dvss.n3014 dvss.n2864 0.120292
R22689 dvss.n3032 dvss.n2857 0.120292
R22690 dvss.n3037 dvss.n3036 0.120292
R22691 dvss.n3038 dvss.n3037 0.120292
R22692 dvss.n3038 dvss.n2853 0.120292
R22693 dvss.n3042 dvss.n2853 0.120292
R22694 dvss.n3043 dvss.n3042 0.120292
R22695 dvss.n3043 dvss.n2850 0.120292
R22696 dvss.n3048 dvss.n2850 0.120292
R22697 dvss.n3121 dvss.n3050 0.120292
R22698 dvss.n3116 dvss.n3050 0.120292
R22699 dvss.n3116 dvss.n3115 0.120292
R22700 dvss.n3115 dvss.n3114 0.120292
R22701 dvss.n3114 dvss.n3052 0.120292
R22702 dvss.n3109 dvss.n3108 0.120292
R22703 dvss.n3108 dvss.n3058 0.120292
R22704 dvss.n3104 dvss.n3058 0.120292
R22705 dvss.n3103 dvss.n3061 0.120292
R22706 dvss.n3095 dvss.n3094 0.120292
R22707 dvss.n3094 dvss.n3066 0.120292
R22708 dvss.n3090 dvss.n3066 0.120292
R22709 dvss.n3090 dvss.n3089 0.120292
R22710 dvss.n3089 dvss.n3088 0.120292
R22711 dvss.n3088 dvss.n3069 0.120292
R22712 dvss.n3084 dvss.n3069 0.120292
R22713 dvss.n3084 dvss.n3083 0.120292
R22714 dvss.n3083 dvss.n3071 0.120292
R22715 dvss.n3079 dvss.n3071 0.120292
R22716 dvss.n3079 dvss.n3078 0.120292
R22717 dvss.n2735 dvss.n2734 0.120292
R22718 dvss.n2740 dvss.n2739 0.120292
R22719 dvss.n2745 dvss.n2705 0.120292
R22720 dvss.n2751 dvss.n2705 0.120292
R22721 dvss.n2752 dvss.n2751 0.120292
R22722 dvss.n2759 dvss.n2758 0.120292
R22723 dvss.n2760 dvss.n2759 0.120292
R22724 dvss.n2760 dvss.n2702 0.120292
R22725 dvss.n2764 dvss.n2702 0.120292
R22726 dvss.n2765 dvss.n2764 0.120292
R22727 dvss.n2765 dvss.n2699 0.120292
R22728 dvss.n2769 dvss.n2699 0.120292
R22729 dvss.n2770 dvss.n2769 0.120292
R22730 dvss.n2770 dvss.n2697 0.120292
R22731 dvss.n2775 dvss.n2697 0.120292
R22732 dvss.n2776 dvss.n2775 0.120292
R22733 dvss.n2781 dvss.n2695 0.120292
R22734 dvss.n2782 dvss.n2781 0.120292
R22735 dvss.n2783 dvss.n2691 0.120292
R22736 dvss.n2792 dvss.n2691 0.120292
R22737 dvss.n2793 dvss.n2792 0.120292
R22738 dvss.n2802 dvss.n2687 0.120292
R22739 dvss.n2803 dvss.n2802 0.120292
R22740 dvss.n2841 dvss.n2840 0.120292
R22741 dvss.n2840 dvss.n2807 0.120292
R22742 dvss.n2833 dvss.n2832 0.120292
R22743 dvss.n2832 dvss.n2814 0.120292
R22744 dvss.n2827 dvss.n2826 0.120292
R22745 dvss.n2826 dvss.n2816 0.120292
R22746 dvss.n3432 dvss.n3431 0.120292
R22747 dvss.n3426 dvss.n2679 0.120292
R22748 dvss.n3422 dvss.n2679 0.120292
R22749 dvss.n3416 dvss.n3415 0.120292
R22750 dvss.n3415 dvss.n3414 0.120292
R22751 dvss.n3409 dvss.n3408 0.120292
R22752 dvss.n3408 dvss.n3341 0.120292
R22753 dvss.n3403 dvss.n3402 0.120292
R22754 dvss.n3402 dvss.n3344 0.120292
R22755 dvss.n3398 dvss.n3344 0.120292
R22756 dvss.n3398 dvss.n3397 0.120292
R22757 dvss.n3397 dvss.n3347 0.120292
R22758 dvss.n3392 dvss.n3391 0.120292
R22759 dvss.n3391 dvss.n3349 0.120292
R22760 dvss.n3385 dvss.n3352 0.120292
R22761 dvss.n3385 dvss.n3384 0.120292
R22762 dvss.n3384 dvss.n3353 0.120292
R22763 dvss.n3377 dvss.n3353 0.120292
R22764 dvss.n3375 dvss.n3357 0.120292
R22765 dvss.n3369 dvss.n3368 0.120292
R22766 dvss.n3368 dvss.n3359 0.120292
R22767 dvss.n3679 dvss.n3678 0.120292
R22768 dvss.n3684 dvss.n3659 0.120292
R22769 dvss.n3685 dvss.n3684 0.120292
R22770 dvss.n3686 dvss.n3685 0.120292
R22771 dvss.n3686 dvss.n3655 0.120292
R22772 dvss.n3694 dvss.n3655 0.120292
R22773 dvss.n3695 dvss.n3694 0.120292
R22774 dvss.n3755 dvss.n3696 0.120292
R22775 dvss.n3751 dvss.n3696 0.120292
R22776 dvss.n3751 dvss.n3750 0.120292
R22777 dvss.n3750 dvss.n3749 0.120292
R22778 dvss.n3749 dvss.n3698 0.120292
R22779 dvss.n3742 dvss.n3698 0.120292
R22780 dvss.n3742 dvss.n3741 0.120292
R22781 dvss.n3741 dvss.n3740 0.120292
R22782 dvss.n3740 dvss.n3700 0.120292
R22783 dvss.n3733 dvss.n3700 0.120292
R22784 dvss.n3733 dvss.n3732 0.120292
R22785 dvss.n3732 dvss.n3731 0.120292
R22786 dvss.n3731 dvss.n3702 0.120292
R22787 dvss.n3727 dvss.n3702 0.120292
R22788 dvss.n3727 dvss.n3726 0.120292
R22789 dvss.n3726 dvss.n3725 0.120292
R22790 dvss.n3725 dvss.n3704 0.120292
R22791 dvss.n3720 dvss.n3704 0.120292
R22792 dvss.n3720 dvss.n3719 0.120292
R22793 dvss.n3714 dvss.n3713 0.120292
R22794 dvss.n3713 dvss.n3710 0.120292
R22795 dvss.n3710 dvss.n3709 0.120292
R22796 dvss.n3764 dvss.n3649 0.120292
R22797 dvss.n3771 dvss.n3649 0.120292
R22798 dvss.n3772 dvss.n3771 0.120292
R22799 dvss.n3773 dvss.n3772 0.120292
R22800 dvss.n3773 dvss.n3646 0.120292
R22801 dvss.n3781 dvss.n3646 0.120292
R22802 dvss.n3782 dvss.n3781 0.120292
R22803 dvss.n3783 dvss.n3782 0.120292
R22804 dvss.n3783 dvss.n3643 0.120292
R22805 dvss.n3789 dvss.n3643 0.120292
R22806 dvss.n3813 dvss.n3812 0.120292
R22807 dvss.n3813 dvss.n3635 0.120292
R22808 dvss.n3819 dvss.n3635 0.120292
R22809 dvss.n3820 dvss.n3819 0.120292
R22810 dvss.n3821 dvss.n3820 0.120292
R22811 dvss.n3825 dvss.n3824 0.120292
R22812 dvss.n3826 dvss.n3825 0.120292
R22813 dvss.n3826 dvss.n3631 0.120292
R22814 dvss.n3836 dvss.n3631 0.120292
R22815 dvss.n3837 dvss.n3836 0.120292
R22816 dvss.n3903 dvss.n3902 0.120292
R22817 dvss.n3902 dvss.n3901 0.120292
R22818 dvss.n3901 dvss.n3840 0.120292
R22819 dvss.n3842 dvss.n3840 0.120292
R22820 dvss.n3894 dvss.n3893 0.120292
R22821 dvss.n3893 dvss.n3845 0.120292
R22822 dvss.n3887 dvss.n3845 0.120292
R22823 dvss.n3887 dvss.n3886 0.120292
R22824 dvss.n3886 dvss.n3885 0.120292
R22825 dvss.n3885 dvss.n3847 0.120292
R22826 dvss.n3881 dvss.n3880 0.120292
R22827 dvss.n3879 dvss.n3850 0.120292
R22828 dvss.n3875 dvss.n3850 0.120292
R22829 dvss.n3875 dvss.n3874 0.120292
R22830 dvss.n3874 dvss.n3873 0.120292
R22831 dvss.n3873 dvss.n3855 0.120292
R22832 dvss.n3857 dvss.n3855 0.120292
R22833 dvss.n3867 dvss.n3857 0.120292
R22834 dvss.n3866 dvss.n3865 0.120292
R22835 dvss.n3542 dvss.n3541 0.120292
R22836 dvss.n3547 dvss.n3546 0.120292
R22837 dvss.n3557 dvss.n3530 0.120292
R22838 dvss.n3563 dvss.n3530 0.120292
R22839 dvss.n3564 dvss.n3563 0.120292
R22840 dvss.n3565 dvss.n3564 0.120292
R22841 dvss.n3569 dvss.n3524 0.120292
R22842 dvss.n3574 dvss.n3524 0.120292
R22843 dvss.n3575 dvss.n3574 0.120292
R22844 dvss.n3576 dvss.n3575 0.120292
R22845 dvss.n3591 dvss.n3590 0.120292
R22846 dvss.n3591 dvss.n3519 0.120292
R22847 dvss.n3595 dvss.n3519 0.120292
R22848 dvss.n3596 dvss.n3595 0.120292
R22849 dvss.n3602 dvss.n3601 0.120292
R22850 dvss.n3603 dvss.n3602 0.120292
R22851 dvss.n3603 dvss.n3513 0.120292
R22852 dvss.n3609 dvss.n3513 0.120292
R22853 dvss.n3614 dvss.n3613 0.120292
R22854 dvss.n3509 dvss.n3507 0.120292
R22855 dvss.n3624 dvss.n3507 0.120292
R22856 dvss.n3499 dvss.n3498 0.120292
R22857 dvss.n3495 dvss.n3494 0.120292
R22858 dvss.n3490 dvss.n3489 0.120292
R22859 dvss.n3489 dvss.n3488 0.120292
R22860 dvss.n3488 dvss.n3474 0.120292
R22861 dvss.n3996 dvss.n3995 0.120292
R22862 dvss.n3995 dvss.n3994 0.120292
R22863 dvss.n3994 dvss.n3456 0.120292
R22864 dvss.n3989 dvss.n3988 0.120292
R22865 dvss.n3988 dvss.n3458 0.120292
R22866 dvss.n3984 dvss.n3458 0.120292
R22867 dvss.n3984 dvss.n3983 0.120292
R22868 dvss.n3983 dvss.n3982 0.120292
R22869 dvss.n3982 dvss.n3463 0.120292
R22870 dvss.n3974 dvss.n3909 0.120292
R22871 dvss.n3968 dvss.n3967 0.120292
R22872 dvss.n3966 dvss.n3911 0.120292
R22873 dvss.n3960 dvss.n3911 0.120292
R22874 dvss.n3960 dvss.n3959 0.120292
R22875 dvss.n3959 dvss.n3958 0.120292
R22876 dvss.n3958 dvss.n3914 0.120292
R22877 dvss.n3950 dvss.n3914 0.120292
R22878 dvss.n3950 dvss.n3949 0.120292
R22879 dvss.n3949 dvss.n3948 0.120292
R22880 dvss.n3948 dvss.n3916 0.120292
R22881 dvss.n3942 dvss.n3916 0.120292
R22882 dvss.n3942 dvss.n3941 0.120292
R22883 dvss.n3941 dvss.n3940 0.120292
R22884 dvss.n3940 dvss.n3918 0.120292
R22885 dvss.n3936 dvss.n3918 0.120292
R22886 dvss.n3936 dvss.n3935 0.120292
R22887 dvss.n3931 dvss.n3930 0.120292
R22888 dvss.n3930 dvss.n3929 0.120292
R22889 dvss.n2343 dvss.n2342 0.120292
R22890 dvss.n2343 dvss.n2333 0.120292
R22891 dvss.n2347 dvss.n2333 0.120292
R22892 dvss.n2348 dvss.n2347 0.120292
R22893 dvss.n2349 dvss.n2348 0.120292
R22894 dvss.n2349 dvss.n2331 0.120292
R22895 dvss.n2354 dvss.n2331 0.120292
R22896 dvss.n2355 dvss.n2354 0.120292
R22897 dvss.n2356 dvss.n2355 0.120292
R22898 dvss.n2356 dvss.n2329 0.120292
R22899 dvss.n2361 dvss.n2329 0.120292
R22900 dvss.n4486 dvss.n4485 0.120292
R22901 dvss.n4485 dvss.n2363 0.120292
R22902 dvss.n4481 dvss.n2363 0.120292
R22903 dvss.n4481 dvss.n4480 0.120292
R22904 dvss.n4480 dvss.n4479 0.120292
R22905 dvss.n4479 dvss.n2365 0.120292
R22906 dvss.n4474 dvss.n2365 0.120292
R22907 dvss.n4474 dvss.n4473 0.120292
R22908 dvss.n4473 dvss.n4472 0.120292
R22909 dvss.n4472 dvss.n2369 0.120292
R22910 dvss.n4466 dvss.n4465 0.120292
R22911 dvss.n4465 dvss.n2372 0.120292
R22912 dvss.n4461 dvss.n2372 0.120292
R22913 dvss.n4461 dvss.n4460 0.120292
R22914 dvss.n4460 dvss.n4459 0.120292
R22915 dvss.n4459 dvss.n2374 0.120292
R22916 dvss.n4455 dvss.n2374 0.120292
R22917 dvss.n4455 dvss.n4454 0.120292
R22918 dvss.n4451 dvss.n4450 0.120292
R22919 dvss.n4446 dvss.n4445 0.120292
R22920 dvss.n4445 dvss.n2382 0.120292
R22921 dvss dvss.n2382 0.120292
R22922 dvss.n4440 dvss.n2387 0.120292
R22923 dvss.n4435 dvss.n4434 0.120292
R22924 dvss.n4430 dvss.n4429 0.120292
R22925 dvss.n4429 dvss.n2395 0.120292
R22926 dvss.n4424 dvss.n2395 0.120292
R22927 dvss.n4424 dvss.n4423 0.120292
R22928 dvss.n4423 dvss.n4422 0.120292
R22929 dvss.n4422 dvss.n2398 0.120292
R22930 dvss.n4407 dvss.n4298 0.120292
R22931 dvss.n4403 dvss.n4298 0.120292
R22932 dvss.n4403 dvss.n4402 0.120292
R22933 dvss.n4305 dvss.n4303 0.120292
R22934 dvss.n4397 dvss.n4305 0.120292
R22935 dvss.n4395 dvss.n4307 0.120292
R22936 dvss.n4388 dvss.n4307 0.120292
R22937 dvss.n4382 dvss.n4381 0.120292
R22938 dvss.n4381 dvss.n4318 0.120292
R22939 dvss.n4372 dvss.n4321 0.120292
R22940 dvss.n4367 dvss.n4321 0.120292
R22941 dvss.n4367 dvss.n4366 0.120292
R22942 dvss.n4366 dvss.n4365 0.120292
R22943 dvss.n4365 dvss.n4323 0.120292
R22944 dvss.n4360 dvss.n4323 0.120292
R22945 dvss.n4360 dvss.n4359 0.120292
R22946 dvss.n4359 dvss.n4358 0.120292
R22947 dvss.n4355 dvss.n4354 0.120292
R22948 dvss.n4354 dvss.n4353 0.120292
R22949 dvss.n4349 dvss.n4348 0.120292
R22950 dvss.n4343 dvss.n4336 0.120292
R22951 dvss.n4510 dvss.n4509 0.120292
R22952 dvss.n4510 dvss.n4497 0.120292
R22953 dvss.n4514 dvss.n4497 0.120292
R22954 dvss.n4522 dvss.n4494 0.120292
R22955 dvss.n4523 dvss.n4522 0.120292
R22956 dvss.n4786 dvss.n4785 0.120292
R22957 dvss.n4785 dvss.n4524 0.120292
R22958 dvss.n4779 dvss.n4778 0.120292
R22959 dvss.n4778 dvss.n4527 0.120292
R22960 dvss.n4774 dvss.n4527 0.120292
R22961 dvss.n4774 dvss.n4773 0.120292
R22962 dvss.n4770 dvss.n4769 0.120292
R22963 dvss.n4769 dvss.n4531 0.120292
R22964 dvss.n4764 dvss.n4531 0.120292
R22965 dvss.n4764 dvss.n4763 0.120292
R22966 dvss.n4763 dvss.n4762 0.120292
R22967 dvss.n4762 dvss.n4533 0.120292
R22968 dvss.n4757 dvss.n4756 0.120292
R22969 dvss.n4756 dvss.n4535 0.120292
R22970 dvss.n4752 dvss.n4535 0.120292
R22971 dvss.n4752 dvss.n4751 0.120292
R22972 dvss.n4746 dvss.n4745 0.120292
R22973 dvss.n4745 dvss.n4539 0.120292
R22974 dvss.n4740 dvss.n4539 0.120292
R22975 dvss.n4740 dvss.n4739 0.120292
R22976 dvss.n4739 dvss.n4738 0.120292
R22977 dvss.n4734 dvss.n4733 0.120292
R22978 dvss.n4733 dvss.n4548 0.120292
R22979 dvss.n4728 dvss.n4727 0.120292
R22980 dvss.n4727 dvss.n4553 0.120292
R22981 dvss.n4721 dvss.n4720 0.120292
R22982 dvss.n4720 dvss.n4555 0.120292
R22983 dvss.n4714 dvss.n4713 0.120292
R22984 dvss.n4700 dvss.n4699 0.120292
R22985 dvss.n4699 dvss.n4581 0.120292
R22986 dvss.n4693 dvss.n4692 0.120292
R22987 dvss.n4692 dvss.n4584 0.120292
R22988 dvss.n4688 dvss.n4584 0.120292
R22989 dvss.n4688 dvss.n4687 0.120292
R22990 dvss.n4687 dvss.n4589 0.120292
R22991 dvss.n4680 dvss.n4679 0.120292
R22992 dvss.n4674 dvss.n4673 0.120292
R22993 dvss.n4673 dvss.n4601 0.120292
R22994 dvss.n4668 dvss.n4601 0.120292
R22995 dvss.n4668 dvss.n4667 0.120292
R22996 dvss.n4658 dvss.n4613 0.120292
R22997 dvss.n4651 dvss.n4650 0.120292
R22998 dvss.n4650 dvss.n4615 0.120292
R22999 dvss.n4646 dvss.n4615 0.120292
R23000 dvss.n4646 dvss.n4645 0.120292
R23001 dvss.n4645 dvss.n4644 0.120292
R23002 dvss.n4641 dvss.n4640 0.120292
R23003 dvss.n4640 dvss.n4621 0.120292
R23004 dvss.n4633 dvss.n4632 0.120292
R23005 dvss.n4632 dvss.n4624 0.120292
R23006 dvss.n4870 dvss.n4869 0.120292
R23007 dvss.n4875 dvss.n4874 0.120292
R23008 dvss.n4875 dvss.n4862 0.120292
R23009 dvss.n4879 dvss.n4862 0.120292
R23010 dvss.n4880 dvss.n4879 0.120292
R23011 dvss.n4881 dvss.n4880 0.120292
R23012 dvss.n4881 dvss.n4860 0.120292
R23013 dvss.n4885 dvss.n4860 0.120292
R23014 dvss.n4886 dvss.n4885 0.120292
R23015 dvss.n4886 dvss.n4858 0.120292
R23016 dvss.n4891 dvss.n4858 0.120292
R23017 dvss.n4892 dvss.n4891 0.120292
R23018 dvss.n4999 dvss.n4894 0.120292
R23019 dvss.n4999 dvss.n4998 0.120292
R23020 dvss.n4998 dvss.n4997 0.120292
R23021 dvss.n4994 dvss.n4993 0.120292
R23022 dvss.n4993 dvss.n4898 0.120292
R23023 dvss.n4986 dvss.n4899 0.120292
R23024 dvss.n4986 dvss.n4985 0.120292
R23025 dvss.n4985 dvss.n4984 0.120292
R23026 dvss.n4981 dvss.n4980 0.120292
R23027 dvss.n4980 dvss.n4903 0.120292
R23028 dvss.n4973 dvss.n4904 0.120292
R23029 dvss.n4973 dvss.n4972 0.120292
R23030 dvss.n4972 dvss.n4971 0.120292
R23031 dvss.n4968 dvss.n4967 0.120292
R23032 dvss.n4967 dvss.n4908 0.120292
R23033 dvss.n4960 dvss.n4909 0.120292
R23034 dvss.n4960 dvss.n4959 0.120292
R23035 dvss.n4959 dvss.n4958 0.120292
R23036 dvss.n4955 dvss.n4954 0.120292
R23037 dvss.n4952 dvss.n4913 0.120292
R23038 dvss.n4948 dvss.n4913 0.120292
R23039 dvss.n4948 dvss.n4947 0.120292
R23040 dvss.n4947 dvss.n4946 0.120292
R23041 dvss.n4943 dvss.n4942 0.120292
R23042 dvss.n4942 dvss.n4917 0.120292
R23043 dvss.n4936 dvss.n4935 0.120292
R23044 dvss.n4935 dvss.n4934 0.120292
R23045 dvss.n4934 dvss.n4919 0.120292
R23046 dvss.n5090 dvss.n5089 0.120292
R23047 dvss.n5089 dvss.n1221 0.120292
R23048 dvss.n5084 dvss.n5083 0.120292
R23049 dvss.n5083 dvss.n1224 0.120292
R23050 dvss.n5078 dvss.n5077 0.120292
R23051 dvss.n5077 dvss.n1226 0.120292
R23052 dvss.n5073 dvss.n1226 0.120292
R23053 dvss.n5071 dvss.n5005 0.120292
R23054 dvss.n5066 dvss.n5005 0.120292
R23055 dvss.n5066 dvss.n5065 0.120292
R23056 dvss.n5065 dvss.n5064 0.120292
R23057 dvss.n5064 dvss.n5008 0.120292
R23058 dvss.n5060 dvss.n5059 0.120292
R23059 dvss.n5058 dvss.n5012 0.120292
R23060 dvss.n5052 dvss.n5012 0.120292
R23061 dvss.n5052 dvss.n5051 0.120292
R23062 dvss.n5051 dvss.n5050 0.120292
R23063 dvss.n5050 dvss.n5014 0.120292
R23064 dvss.n5044 dvss.n5014 0.120292
R23065 dvss.n5044 dvss.n5043 0.120292
R23066 dvss.n5043 dvss.n5042 0.120292
R23067 dvss.n5042 dvss.n5016 0.120292
R23068 dvss.n5037 dvss.n5036 0.120292
R23069 dvss.n5036 dvss.n5020 0.120292
R23070 dvss.n5030 dvss.n5029 0.120292
R23071 dvss.n5029 dvss.n5025 0.120292
R23072 dvss.n4068 dvss.n4067 0.120292
R23073 dvss.n4068 dvss.n4055 0.120292
R23074 dvss.n4074 dvss.n4055 0.120292
R23075 dvss.n4075 dvss.n4074 0.120292
R23076 dvss.n4079 dvss.n4052 0.120292
R23077 dvss.n4086 dvss.n4052 0.120292
R23078 dvss.n4047 dvss.n4045 0.120292
R23079 dvss.n4095 dvss.n4094 0.120292
R23080 dvss.n4096 dvss.n4095 0.120292
R23081 dvss.n4096 dvss.n4042 0.120292
R23082 dvss.n4102 dvss.n4042 0.120292
R23083 dvss.n4104 dvss.n4040 0.120292
R23084 dvss.n4040 dvss.n4038 0.120292
R23085 dvss.n4109 dvss.n4038 0.120292
R23086 dvss.n4110 dvss.n4109 0.120292
R23087 dvss.n4110 dvss.n4035 0.120292
R23088 dvss.n4118 dvss.n4035 0.120292
R23089 dvss.n4120 dvss.n4119 0.120292
R23090 dvss.n4120 dvss.n4033 0.120292
R23091 dvss.n4032 dvss.n4030 0.120292
R23092 dvss.n4126 dvss.n4030 0.120292
R23093 dvss.n4127 dvss.n4126 0.120292
R23094 dvss.n4128 dvss.n4027 0.120292
R23095 dvss.n4136 dvss.n4027 0.120292
R23096 dvss.n4137 dvss.n4136 0.120292
R23097 dvss.n4189 dvss.n4188 0.120292
R23098 dvss.n4188 dvss.n4138 0.120292
R23099 dvss.n4182 dvss.n4138 0.120292
R23100 dvss.n4180 dvss.n4143 0.120292
R23101 dvss.n4145 dvss.n4143 0.120292
R23102 dvss.n4146 dvss.n4145 0.120292
R23103 dvss.n4149 dvss.n4146 0.120292
R23104 dvss.n4172 dvss.n4149 0.120292
R23105 dvss.n4288 dvss.n4012 0.120292
R23106 dvss.n4283 dvss.n4012 0.120292
R23107 dvss.n4283 dvss.n4282 0.120292
R23108 dvss.n4278 dvss.n4018 0.120292
R23109 dvss.n4278 dvss.n4277 0.120292
R23110 dvss.n4277 dvss.n4276 0.120292
R23111 dvss.n4276 dvss.n4022 0.120292
R23112 dvss.n4270 dvss.n4269 0.120292
R23113 dvss.n4269 dvss.n4268 0.120292
R23114 dvss.n4263 dvss.n4197 0.120292
R23115 dvss.n4258 dvss.n4197 0.120292
R23116 dvss.n4251 dvss.n4250 0.120292
R23117 dvss.n4250 dvss.n4249 0.120292
R23118 dvss.n4249 dvss.n4203 0.120292
R23119 dvss.n4245 dvss.n4203 0.120292
R23120 dvss.n4245 dvss.n4244 0.120292
R23121 dvss.n4244 dvss.n4243 0.120292
R23122 dvss.n4243 dvss.n4205 0.120292
R23123 dvss.n4239 dvss.n4205 0.120292
R23124 dvss.n4239 dvss.n4238 0.120292
R23125 dvss.n4234 dvss.n4233 0.120292
R23126 dvss.n4233 dvss.n4232 0.120292
R23127 dvss.n4232 dvss.n4212 0.120292
R23128 dvss.n4215 dvss.n4212 0.120292
R23129 dvss.n4225 dvss.n4215 0.120292
R23130 dvss.n4224 dvss.n4223 0.120292
R23131 dvss.n290 dvss.n285 0.120292
R23132 dvss.n297 dvss.n285 0.120292
R23133 dvss.n298 dvss.n297 0.120292
R23134 dvss.n299 dvss.n298 0.120292
R23135 dvss.n299 dvss.n282 0.120292
R23136 dvss.n306 dvss.n282 0.120292
R23137 dvss.n307 dvss.n306 0.120292
R23138 dvss.n331 dvss.n307 0.120292
R23139 dvss.n331 dvss.n330 0.120292
R23140 dvss.n330 dvss.n308 0.120292
R23141 dvss.n325 dvss.n308 0.120292
R23142 dvss.n325 dvss.n324 0.120292
R23143 dvss.n321 dvss.n320 0.120292
R23144 dvss.n320 dvss.n312 0.120292
R23145 dvss.n316 dvss.n312 0.120292
R23146 dvss.n316 dvss.n315 0.120292
R23147 dvss.n402 dvss.n401 0.120292
R23148 dvss.n403 dvss.n402 0.120292
R23149 dvss.n403 dvss.n392 0.120292
R23150 dvss.n410 dvss.n392 0.120292
R23151 dvss.n411 dvss.n410 0.120292
R23152 dvss.n412 dvss.n411 0.120292
R23153 dvss.n412 dvss.n389 0.120292
R23154 dvss.n439 dvss.n389 0.120292
R23155 dvss.n440 dvss.n439 0.120292
R23156 dvss.n440 dvss.n385 0.120292
R23157 dvss.n445 dvss.n385 0.120292
R23158 dvss.n446 dvss.n445 0.120292
R23159 dvss.n451 dvss.n450 0.120292
R23160 dvss.n452 dvss.n451 0.120292
R23161 dvss.n452 dvss.n381 0.120292
R23162 dvss.n456 dvss.n381 0.120292
R23163 dvss.n264 dvss.n263 0.120292
R23164 dvss.n265 dvss.n264 0.120292
R23165 dvss.n265 dvss.n254 0.120292
R23166 dvss.n272 dvss.n254 0.120292
R23167 dvss.n273 dvss.n272 0.120292
R23168 dvss.n274 dvss.n273 0.120292
R23169 dvss.n274 dvss.n251 0.120292
R23170 dvss.n6614 dvss.n251 0.120292
R23171 dvss.n6615 dvss.n6614 0.120292
R23172 dvss.n6615 dvss.n247 0.120292
R23173 dvss.n6620 dvss.n247 0.120292
R23174 dvss.n6621 dvss.n6620 0.120292
R23175 dvss.n6626 dvss.n6625 0.120292
R23176 dvss.n6627 dvss.n6626 0.120292
R23177 dvss.n6627 dvss.n243 0.120292
R23178 dvss.n6631 dvss.n243 0.120292
R23179 dvss.n352 dvss.n351 0.120292
R23180 dvss.n353 dvss.n352 0.120292
R23181 dvss.n353 dvss.n342 0.120292
R23182 dvss.n360 dvss.n342 0.120292
R23183 dvss.n361 dvss.n360 0.120292
R23184 dvss.n362 dvss.n361 0.120292
R23185 dvss.n362 dvss.n339 0.120292
R23186 dvss.n369 dvss.n339 0.120292
R23187 dvss.n370 dvss.n369 0.120292
R23188 dvss.n6601 dvss.n370 0.120292
R23189 dvss.n6601 dvss.n6600 0.120292
R23190 dvss.n6600 dvss.n6599 0.120292
R23191 dvss.n6596 dvss.n6595 0.120292
R23192 dvss.n6595 dvss.n373 0.120292
R23193 dvss.n6591 dvss.n373 0.120292
R23194 dvss.n6591 dvss.n6590 0.120292
R23195 dvss.n6587 dvss.n6586 0.120292
R23196 dvss.n6586 dvss.n377 0.120292
R23197 dvss.n6582 dvss.n377 0.120292
R23198 dvss.n6582 dvss.n6581 0.120292
R23199 dvss.n2458 dvss 0.105238
R23200 dvss.n2882 dvss 0.105238
R23201 dvss.n2716 dvss 0.105238
R23202 dvss.n3667 dvss 0.105238
R23203 dvss.n3540 dvss 0.105238
R23204 dvss.n2338 dvss 0.105238
R23205 dvss.n4503 dvss 0.105238
R23206 dvss.n4062 dvss 0.105238
R23207 dvss.n7013 dvss.n7012 0.101043
R23208 dvss.n7007 dvss.n7006 0.100247
R23209 dvss.n2640 dvss 0.0994583
R23210 dvss.n2734 dvss 0.0994583
R23211 dvss.n2739 dvss 0.0994583
R23212 dvss.n7009 dvss.n7008 0.0989849
R23213 dvss.n2481 dvss 0.0981562
R23214 dvss.n2526 dvss 0.0981562
R23215 dvss dvss.n2430 0.0981562
R23216 dvss.n2422 dvss 0.0981562
R23217 dvss.n2912 dvss 0.0981562
R23218 dvss.n2975 dvss 0.0981562
R23219 dvss.n2960 dvss 0.0981562
R23220 dvss.n2729 dvss 0.0981562
R23221 dvss dvss.n2695 0.0981562
R23222 dvss dvss.n2687 0.0981562
R23223 dvss dvss.n3426 0.0981562
R23224 dvss.n3352 dvss 0.0981562
R23225 dvss dvss.n3375 0.0981562
R23226 dvss.n3673 dvss 0.0981562
R23227 dvss.n3715 dvss 0.0981562
R23228 dvss dvss.n3894 0.0981562
R23229 dvss.n3551 dvss 0.0981562
R23230 dvss.n3556 dvss 0.0981562
R23231 dvss.n3590 dvss 0.0981562
R23232 dvss.n3610 dvss 0.0981562
R23233 dvss dvss.n3509 0.0981562
R23234 dvss.n3626 dvss 0.0981562
R23235 dvss dvss.n3499 0.0981562
R23236 dvss.n3490 dvss 0.0981562
R23237 dvss.n3931 dvss 0.0981562
R23238 dvss.n2362 dvss 0.0981562
R23239 dvss.n4466 dvss 0.0981562
R23240 dvss.n4446 dvss 0.0981562
R23241 dvss dvss.n4430 0.0981562
R23242 dvss.n4355 dvss 0.0981562
R23243 dvss dvss.n4344 0.0981562
R23244 dvss.n4787 dvss 0.0981562
R23245 dvss.n4770 dvss 0.0981562
R23246 dvss.n4757 dvss 0.0981562
R23247 dvss.n4747 dvss 0.0981562
R23248 dvss.n4659 dvss 0.0981562
R23249 dvss.n4869 dvss 0.0981562
R23250 dvss.n4893 dvss 0.0981562
R23251 dvss dvss.n5084 0.0981562
R23252 dvss dvss.n4047 0.0981562
R23253 dvss.n4104 dvss 0.0981562
R23254 dvss dvss.n4180 0.0981562
R23255 dvss.n4251 dvss 0.0981562
R23256 dvss.n4234 dvss 0.0981562
R23257 dvss.n2993 dvss 0.0968542
R23258 dvss dvss.n2833 0.0968542
R23259 dvss.n3678 dvss 0.0968542
R23260 dvss dvss.n4349 0.0968542
R23261 dvss dvss.n4746 0.0968542
R23262 dvss dvss.n4728 0.0968542
R23263 dvss dvss.n4263 0.0968542
R23264 dvss.n2662 dvss.n2661 0.0950946
R23265 dvss.n2655 dvss.n2413 0.0950946
R23266 dvss.n3018 dvss.n3017 0.0950946
R23267 dvss.n3026 dvss.n2860 0.0950946
R23268 dvss.n3444 dvss.n3443 0.0950946
R23269 dvss.n3437 dvss.n2672 0.0950946
R23270 dvss.n3793 dvss.n3792 0.0950946
R23271 dvss.n3810 dvss.n3638 0.0950946
R23272 dvss.n3480 dvss.n3478 0.0950946
R23273 dvss.n4002 dvss.n3449 0.0950946
R23274 dvss.n4415 dvss.n2404 0.0950946
R23275 dvss.n4409 dvss.n4294 0.0950946
R23276 dvss.n4711 dvss.n4560 0.0950946
R23277 dvss.n4706 dvss.n4563 0.0950946
R23278 dvss.n4928 dvss.n4926 0.0950946
R23279 dvss.n5095 dvss.n1213 0.0950946
R23280 dvss.n4169 dvss.n4168 0.0950946
R23281 dvss.n4290 dvss.n4010 0.0950946
R23282 dvss.n2650 dvss.n2414 0.0916458
R23283 dvss.n3027 dvss.n2857 0.0916458
R23284 dvss.n3432 dvss.n2673 0.0916458
R23285 dvss.n3812 dvss.n3811 0.0916458
R23286 dvss.n3996 dvss.n3452 0.0916458
R23287 dvss.n4408 dvss.n4407 0.0916458
R23288 dvss.n5090 dvss.n1217 0.0916458
R23289 dvss.n4289 dvss.n4288 0.0916458
R23290 dvss.n4489 dvss.n2327 0.0900105
R23291 dvss.n7034 dvss.n6997 0.0888838
R23292 dvss.n2660 dvss.n2659 0.0838333
R23293 dvss.n3021 dvss.n3019 0.0838333
R23294 dvss.n4416 dvss.n2402 0.0838333
R23295 dvss.n4571 dvss.n4569 0.0838333
R23296 dvss.n4929 dvss.n4925 0.0838333
R23297 dvss.n4167 dvss.n4166 0.0838333
R23298 dvss.n7048 dvss.n6996 0.0808571
R23299 dvss.n2322 dvss.n2312 0.0793043
R23300 dvss.n4582 dvss.n4580 0.0700652
R23301 dvss.n2658 dvss.n2410 0.0680676
R23302 dvss.n2658 dvss.n2657 0.0680676
R23303 dvss.n3022 dvss.n2862 0.0680676
R23304 dvss.n3023 dvss.n3022 0.0680676
R23305 dvss.n3440 dvss.n2669 0.0680676
R23306 dvss.n3440 dvss.n3439 0.0680676
R23307 dvss.n3806 dvss.n3640 0.0680676
R23308 dvss.n3807 dvss.n3806 0.0680676
R23309 dvss.n3479 dvss.n3451 0.0680676
R23310 dvss.n4003 dvss.n3451 0.0680676
R23311 dvss.n4414 dvss.n2405 0.0680676
R23312 dvss.n4293 dvss.n2405 0.0680676
R23313 dvss.n4570 dvss.n4561 0.0680676
R23314 dvss.n4570 dvss.n4562 0.0680676
R23315 dvss.n4927 dvss.n1215 0.0680676
R23316 dvss.n5096 dvss.n1215 0.0680676
R23317 dvss.n4165 dvss.n4154 0.0680676
R23318 dvss.n4165 dvss.n4164 0.0680676
R23319 dvss dvss.n3333 0.067223
R23320 dvss.n3139 dvss 0.067223
R23321 dvss.n3140 dvss 0.067223
R23322 dvss.n3141 dvss 0.067223
R23323 dvss.n3142 dvss 0.067223
R23324 dvss.n3147 dvss 0.067223
R23325 dvss.n3148 dvss 0.067223
R23326 dvss.n3149 dvss 0.067223
R23327 dvss dvss.n3155 0.067223
R23328 dvss.n3268 dvss 0.067223
R23329 dvss.n3269 dvss 0.067223
R23330 dvss.n3284 dvss 0.067223
R23331 dvss.n3287 dvss 0.067223
R23332 dvss.n3288 dvss 0.067223
R23333 dvss.n3200 dvss 0.067223
R23334 dvss.n3203 dvss 0.067223
R23335 dvss dvss.n3202 0.067223
R23336 dvss.n3218 dvss 0.067223
R23337 dvss dvss.n3182 0.067223
R23338 dvss.n3243 dvss 0.067223
R23339 dvss.n3244 dvss 0.067223
R23340 dvss.n3257 dvss 0.067223
R23341 dvss.n3258 dvss 0.067223
R23342 dvss.n3261 dvss 0.067223
R23343 dvss dvss.n3260 0.067223
R23344 dvss dvss.n3259 0.067223
R23345 dvss.n6634 dvss 0.067223
R23346 dvss.n1208 dvss 0.067223
R23347 dvss.n5103 dvss 0.067223
R23348 dvss.n5104 dvss 0.067223
R23349 dvss.n5105 dvss 0.067223
R23350 dvss.n5106 dvss 0.067223
R23351 dvss.n5107 dvss 0.067223
R23352 dvss.n5108 dvss 0.067223
R23353 dvss.n5109 dvss 0.067223
R23354 dvss.n5110 dvss 0.067223
R23355 dvss.n5111 dvss 0.067223
R23356 dvss.n5119 dvss 0.067223
R23357 dvss.n5120 dvss 0.067223
R23358 dvss.n5129 dvss 0.067223
R23359 dvss.n5131 dvss 0.067223
R23360 dvss.n5139 dvss 0.067223
R23361 dvss.n5140 dvss 0.067223
R23362 dvss.n5141 dvss 0.067223
R23363 dvss.n5142 dvss 0.067223
R23364 dvss.n5143 dvss 0.067223
R23365 dvss.n5144 dvss 0.067223
R23366 dvss.n5145 dvss 0.067223
R23367 dvss.n5148 dvss 0.067223
R23368 dvss.n5151 dvss 0.067223
R23369 dvss.n5152 dvss 0.067223
R23370 dvss.n5166 dvss 0.067223
R23371 dvss.n5167 dvss 0.067223
R23372 dvss.n5168 dvss 0.067223
R23373 dvss.n5170 dvss 0.067223
R23374 dvss.n5178 dvss 0.067223
R23375 dvss.n5179 dvss 0.067223
R23376 dvss.n5180 dvss 0.067223
R23377 dvss.n5181 dvss 0.067223
R23378 dvss.n5182 dvss 0.067223
R23379 dvss.n5183 dvss 0.067223
R23380 dvss.n5184 dvss 0.067223
R23381 dvss.n5187 dvss 0.067223
R23382 dvss.n5190 dvss 0.067223
R23383 dvss.n5191 dvss 0.067223
R23384 dvss.n5205 dvss 0.067223
R23385 dvss.n5206 dvss 0.067223
R23386 dvss.n5207 dvss 0.067223
R23387 dvss.n5209 dvss 0.067223
R23388 dvss.n5217 dvss 0.067223
R23389 dvss.n5218 dvss 0.067223
R23390 dvss.n5219 dvss 0.067223
R23391 dvss.n5220 dvss 0.067223
R23392 dvss.n5221 dvss 0.067223
R23393 dvss.n5222 dvss 0.067223
R23394 dvss.n5223 dvss 0.067223
R23395 dvss.n5226 dvss 0.067223
R23396 dvss.n5229 dvss 0.067223
R23397 dvss.n5230 dvss 0.067223
R23398 dvss.n5244 dvss 0.067223
R23399 dvss.n5245 dvss 0.067223
R23400 dvss.n5246 dvss 0.067223
R23401 dvss.n5248 dvss 0.067223
R23402 dvss.n5256 dvss 0.067223
R23403 dvss.n5257 dvss 0.067223
R23404 dvss.n5258 dvss 0.067223
R23405 dvss.n5259 dvss 0.067223
R23406 dvss.n5260 dvss 0.067223
R23407 dvss.n5261 dvss 0.067223
R23408 dvss.n5262 dvss 0.067223
R23409 dvss.n5265 dvss 0.067223
R23410 dvss.n5268 dvss 0.067223
R23411 dvss.n5269 dvss 0.067223
R23412 dvss.n5283 dvss 0.067223
R23413 dvss.n5284 dvss 0.067223
R23414 dvss.n5286 dvss 0.067223
R23415 dvss.n5499 dvss 0.067223
R23416 dvss.n5507 dvss 0.067223
R23417 dvss dvss.n5506 0.067223
R23418 dvss.n5515 dvss 0.067223
R23419 dvss.n5516 dvss 0.067223
R23420 dvss.n5518 dvss 0.067223
R23421 dvss dvss.n5517 0.067223
R23422 dvss.n5526 dvss 0.067223
R23423 dvss.n1128 dvss 0.067223
R23424 dvss dvss.n1134 0.067223
R23425 dvss.n1135 dvss 0.067223
R23426 dvss.n5545 dvss 0.067223
R23427 dvss.n5546 dvss 0.067223
R23428 dvss.n5547 dvss 0.067223
R23429 dvss.n5553 dvss 0.067223
R23430 dvss.n5560 dvss 0.067223
R23431 dvss.n5566 dvss 0.067223
R23432 dvss.n5567 dvss 0.067223
R23433 dvss.n5568 dvss 0.067223
R23434 dvss.n5570 dvss 0.067223
R23435 dvss dvss.n5569 0.067223
R23436 dvss.n6212 dvss 0.067223
R23437 dvss dvss.n6216 0.067223
R23438 dvss dvss.n515 0.067223
R23439 dvss.n6235 dvss 0.067223
R23440 dvss.n6244 dvss 0.067223
R23441 dvss.n6245 dvss 0.067223
R23442 dvss.n6247 dvss 0.067223
R23443 dvss.n6256 dvss 0.067223
R23444 dvss dvss.n6262 0.067223
R23445 dvss.n6271 dvss 0.067223
R23446 dvss.n6272 dvss 0.067223
R23447 dvss.n6274 dvss 0.067223
R23448 dvss dvss.n6273 0.067223
R23449 dvss.n6283 dvss 0.067223
R23450 dvss.n6284 dvss 0.067223
R23451 dvss.n6296 dvss 0.067223
R23452 dvss dvss.n6304 0.067223
R23453 dvss dvss.n6303 0.067223
R23454 dvss.n6319 dvss 0.067223
R23455 dvss.n6320 dvss 0.067223
R23456 dvss.n6323 dvss 0.067223
R23457 dvss dvss.n6330 0.067223
R23458 dvss dvss.n6578 0.067223
R23459 dvss.n6575 dvss 0.067223
R23460 dvss dvss.n6574 0.067223
R23461 dvss dvss.n6573 0.067223
R23462 dvss.n464 dvss 0.067223
R23463 dvss.n6345 dvss 0.067223
R23464 dvss.n6564 dvss 0.067223
R23465 dvss.n232 dvss 0.067223
R23466 dvss.n6355 dvss 0.067223
R23467 dvss dvss.n6354 0.067223
R23468 dvss.n6365 dvss 0.067223
R23469 dvss.n6366 dvss 0.067223
R23470 dvss.n6367 dvss 0.067223
R23471 dvss.n6373 dvss 0.067223
R23472 dvss.n6380 dvss 0.067223
R23473 dvss.n6386 dvss 0.067223
R23474 dvss.n6387 dvss 0.067223
R23475 dvss.n6388 dvss 0.067223
R23476 dvss.n6389 dvss 0.067223
R23477 dvss.n6394 dvss 0.067223
R23478 dvss.n6395 dvss 0.067223
R23479 dvss.n6417 dvss 0.067223
R23480 dvss.n6404 dvss 0.067223
R23481 dvss.n6405 dvss 0.067223
R23482 dvss.n6426 dvss 0.067223
R23483 dvss.n6427 dvss 0.067223
R23484 dvss.n6428 dvss 0.067223
R23485 dvss dvss.n3178 0.0663784
R23486 dvss.n2411 dvss.n2409 0.0656042
R23487 dvss.n2654 dvss.n2412 0.0656042
R23488 dvss.n3015 dvss.n2863 0.0656042
R23489 dvss.n3020 dvss.n2859 0.0656042
R23490 dvss.n2670 dvss.n2668 0.0656042
R23491 dvss.n3436 dvss.n2671 0.0656042
R23492 dvss.n3795 dvss.n3790 0.0656042
R23493 dvss.n3482 dvss.n3475 0.0656042
R23494 dvss.n4296 dvss.n4295 0.0656042
R23495 dvss.n4712 dvss.n4559 0.0656042
R23496 dvss.n4930 dvss.n4924 0.0656042
R23497 dvss.n5094 dvss.n1216 0.0656042
R23498 dvss.n4170 dvss.n4152 0.0656042
R23499 dvss.n4163 dvss.n4155 0.0656042
R23500 dvss.n3277 dvss 0.0638446
R23501 dvss.n5159 dvss 0.0638446
R23502 dvss.n5198 dvss 0.0638446
R23503 dvss.n5237 dvss 0.0638446
R23504 dvss.n5276 dvss 0.0638446
R23505 dvss.n5533 dvss 0.0638446
R23506 dvss.n6228 dvss 0.0638446
R23507 dvss.n6298 dvss 0.0638446
R23508 dvss.n6347 dvss 0.0638446
R23509 dvss.n6419 dvss 0.0638446
R23510 dvss dvss.n3329 0.0613108
R23511 dvss.n5138 dvss 0.0613108
R23512 dvss.n5177 dvss 0.0613108
R23513 dvss.n5216 dvss 0.0613108
R23514 dvss.n5255 dvss 0.0613108
R23515 dvss.n5505 dvss 0.0613108
R23516 dvss.n5559 dvss 0.0613108
R23517 dvss.n6263 dvss 0.0613108
R23518 dvss dvss.n458 0.0613108
R23519 dvss.n6379 dvss 0.0613108
R23520 dvss.n2459 dvss 0.0603958
R23521 dvss.n2462 dvss 0.0603958
R23522 dvss dvss.n2446 0.0603958
R23523 dvss.n2492 dvss 0.0603958
R23524 dvss.n2507 dvss 0.0603958
R23525 dvss.n2532 dvss 0.0603958
R23526 dvss.n2562 dvss 0.0603958
R23527 dvss dvss.n2561 0.0603958
R23528 dvss dvss.n2560 0.0603958
R23529 dvss dvss.n2536 0.0603958
R23530 dvss.n2550 dvss 0.0603958
R23531 dvss dvss.n2548 0.0603958
R23532 dvss.n2645 dvss 0.0603958
R23533 dvss.n2639 dvss 0.0603958
R23534 dvss dvss.n2638 0.0603958
R23535 dvss.n2629 dvss 0.0603958
R23536 dvss dvss.n2628 0.0603958
R23537 dvss.n2625 dvss 0.0603958
R23538 dvss.n2608 dvss 0.0603958
R23539 dvss.n2883 dvss 0.0603958
R23540 dvss dvss.n2878 0.0603958
R23541 dvss.n2904 dvss 0.0603958
R23542 dvss.n2985 dvss 0.0603958
R23543 dvss dvss.n2984 0.0603958
R23544 dvss.n2991 dvss 0.0603958
R23545 dvss.n2992 dvss 0.0603958
R23546 dvss.n3007 dvss 0.0603958
R23547 dvss dvss.n3007 0.0603958
R23548 dvss.n3008 dvss 0.0603958
R23549 dvss dvss.n2864 0.0603958
R23550 dvss.n3033 dvss 0.0603958
R23551 dvss.n3036 dvss 0.0603958
R23552 dvss.n3049 dvss 0.0603958
R23553 dvss.n3122 dvss 0.0603958
R23554 dvss dvss.n3121 0.0603958
R23555 dvss.n3109 dvss 0.0603958
R23556 dvss dvss.n3103 0.0603958
R23557 dvss.n3096 dvss 0.0603958
R23558 dvss dvss.n3095 0.0603958
R23559 dvss.n2720 dvss 0.0603958
R23560 dvss.n2727 dvss 0.0603958
R23561 dvss.n2728 dvss 0.0603958
R23562 dvss.n2729 dvss 0.0603958
R23563 dvss.n2733 dvss 0.0603958
R23564 dvss.n2735 dvss 0.0603958
R23565 dvss.n2738 dvss 0.0603958
R23566 dvss.n2740 dvss 0.0603958
R23567 dvss.n2744 dvss 0.0603958
R23568 dvss.n2745 dvss 0.0603958
R23569 dvss.n2758 dvss 0.0603958
R23570 dvss.n2783 dvss 0.0603958
R23571 dvss dvss.n2803 0.0603958
R23572 dvss.n2804 dvss 0.0603958
R23573 dvss.n2842 dvss 0.0603958
R23574 dvss dvss.n2841 0.0603958
R23575 dvss.n2834 dvss 0.0603958
R23576 dvss.n2828 dvss 0.0603958
R23577 dvss dvss.n2827 0.0603958
R23578 dvss.n3428 dvss 0.0603958
R23579 dvss dvss.n3427 0.0603958
R23580 dvss.n3422 dvss 0.0603958
R23581 dvss dvss.n3421 0.0603958
R23582 dvss dvss.n3420 0.0603958
R23583 dvss.n3416 dvss 0.0603958
R23584 dvss.n3339 dvss 0.0603958
R23585 dvss.n3410 dvss 0.0603958
R23586 dvss dvss.n3409 0.0603958
R23587 dvss.n3403 dvss 0.0603958
R23588 dvss.n3392 dvss 0.0603958
R23589 dvss dvss.n3376 0.0603958
R23590 dvss dvss.n3357 0.0603958
R23591 dvss.n3370 dvss 0.0603958
R23592 dvss dvss.n3369 0.0603958
R23593 dvss.n3672 dvss 0.0603958
R23594 dvss.n3674 dvss 0.0603958
R23595 dvss dvss.n3679 0.0603958
R23596 dvss.n3680 dvss 0.0603958
R23597 dvss.n3680 dvss 0.0603958
R23598 dvss dvss.n3659 0.0603958
R23599 dvss.n3757 dvss 0.0603958
R23600 dvss dvss.n3756 0.0603958
R23601 dvss dvss.n3755 0.0603958
R23602 dvss dvss.n3718 0.0603958
R23603 dvss dvss.n3714 0.0603958
R23604 dvss.n3762 dvss 0.0603958
R23605 dvss.n3763 dvss 0.0603958
R23606 dvss.n3764 dvss 0.0603958
R23607 dvss.n3824 dvss 0.0603958
R23608 dvss.n3838 dvss 0.0603958
R23609 dvss.n3903 dvss 0.0603958
R23610 dvss.n3895 dvss 0.0603958
R23611 dvss.n3881 dvss 0.0603958
R23612 dvss dvss.n3879 0.0603958
R23613 dvss dvss.n3866 0.0603958
R23614 dvss.n3541 dvss 0.0603958
R23615 dvss.n3546 dvss 0.0603958
R23616 dvss.n3550 dvss 0.0603958
R23617 dvss.n3555 dvss 0.0603958
R23618 dvss dvss.n3556 0.0603958
R23619 dvss.n3557 dvss 0.0603958
R23620 dvss.n3568 dvss 0.0603958
R23621 dvss.n3569 dvss 0.0603958
R23622 dvss.n3583 dvss 0.0603958
R23623 dvss.n3584 dvss 0.0603958
R23624 dvss.n3589 dvss 0.0603958
R23625 dvss.n3596 dvss 0.0603958
R23626 dvss.n3601 dvss 0.0603958
R23627 dvss.n3613 dvss 0.0603958
R23628 dvss dvss.n3624 0.0603958
R23629 dvss.n3625 dvss 0.0603958
R23630 dvss dvss.n3505 0.0603958
R23631 dvss dvss.n3504 0.0603958
R23632 dvss dvss.n3503 0.0603958
R23633 dvss.n3503 dvss 0.0603958
R23634 dvss.n3500 dvss 0.0603958
R23635 dvss.n3495 dvss 0.0603958
R23636 dvss.n3494 dvss 0.0603958
R23637 dvss dvss.n3493 0.0603958
R23638 dvss.n3990 dvss 0.0603958
R23639 dvss.n3990 dvss 0.0603958
R23640 dvss dvss.n3989 0.0603958
R23641 dvss.n3976 dvss 0.0603958
R23642 dvss dvss.n3975 0.0603958
R23643 dvss dvss.n3974 0.0603958
R23644 dvss.n3968 dvss 0.0603958
R23645 dvss dvss.n3966 0.0603958
R23646 dvss dvss.n3934 0.0603958
R23647 dvss.n2339 dvss 0.0603958
R23648 dvss.n2342 dvss 0.0603958
R23649 dvss.n4486 dvss 0.0603958
R23650 dvss.n4451 dvss 0.0603958
R23651 dvss dvss.n4449 0.0603958
R23652 dvss dvss.n4441 0.0603958
R23653 dvss dvss.n4440 0.0603958
R23654 dvss dvss.n2387 0.0603958
R23655 dvss.n4435 dvss 0.0603958
R23656 dvss.n4431 dvss 0.0603958
R23657 dvss.n4417 dvss 0.0603958
R23658 dvss.n4303 dvss 0.0603958
R23659 dvss dvss.n4396 0.0603958
R23660 dvss dvss.n4395 0.0603958
R23661 dvss dvss.n4387 0.0603958
R23662 dvss.n4383 dvss 0.0603958
R23663 dvss dvss.n4382 0.0603958
R23664 dvss dvss.n4372 0.0603958
R23665 dvss.n4350 dvss 0.0603958
R23666 dvss.n4348 dvss 0.0603958
R23667 dvss.n4345 dvss 0.0603958
R23668 dvss.n4344 dvss 0.0603958
R23669 dvss dvss.n4343 0.0603958
R23670 dvss.n4504 dvss 0.0603958
R23671 dvss.n4505 dvss 0.0603958
R23672 dvss.n4509 dvss 0.0603958
R23673 dvss dvss.n4494 0.0603958
R23674 dvss dvss.n4786 0.0603958
R23675 dvss.n4779 dvss 0.0603958
R23676 dvss.n4544 dvss 0.0603958
R23677 dvss.n4734 dvss 0.0603958
R23678 dvss.n4729 dvss 0.0603958
R23679 dvss.n4721 dvss 0.0603958
R23680 dvss.n4714 dvss 0.0603958
R23681 dvss dvss.n4704 0.0603958
R23682 dvss.n4700 dvss 0.0603958
R23683 dvss.n4693 dvss 0.0603958
R23684 dvss.n4680 dvss 0.0603958
R23685 dvss.n4594 dvss 0.0603958
R23686 dvss.n4675 dvss 0.0603958
R23687 dvss dvss.n4674 0.0603958
R23688 dvss.n4667 dvss 0.0603958
R23689 dvss dvss.n4666 0.0603958
R23690 dvss.n4612 dvss 0.0603958
R23691 dvss dvss.n4658 0.0603958
R23692 dvss dvss.n4613 0.0603958
R23693 dvss.n4652 dvss 0.0603958
R23694 dvss dvss.n4651 0.0603958
R23695 dvss.n4641 dvss 0.0603958
R23696 dvss.n4634 dvss 0.0603958
R23697 dvss dvss.n4633 0.0603958
R23698 dvss dvss.n4870 0.0603958
R23699 dvss.n4871 dvss 0.0603958
R23700 dvss.n4874 dvss 0.0603958
R23701 dvss.n4894 dvss 0.0603958
R23702 dvss.n4994 dvss 0.0603958
R23703 dvss.n4899 dvss 0.0603958
R23704 dvss.n4981 dvss 0.0603958
R23705 dvss.n4904 dvss 0.0603958
R23706 dvss.n4968 dvss 0.0603958
R23707 dvss.n4909 dvss 0.0603958
R23708 dvss.n4955 dvss 0.0603958
R23709 dvss dvss.n4953 0.0603958
R23710 dvss dvss.n4952 0.0603958
R23711 dvss.n4943 dvss 0.0603958
R23712 dvss.n4936 dvss 0.0603958
R23713 dvss.n5085 dvss 0.0603958
R23714 dvss dvss.n1224 0.0603958
R23715 dvss.n5079 dvss 0.0603958
R23716 dvss dvss.n5078 0.0603958
R23717 dvss dvss.n5072 0.0603958
R23718 dvss dvss.n5071 0.0603958
R23719 dvss.n5060 dvss 0.0603958
R23720 dvss dvss.n5058 0.0603958
R23721 dvss.n5038 dvss 0.0603958
R23722 dvss dvss.n5037 0.0603958
R23723 dvss.n5030 dvss 0.0603958
R23724 dvss.n4063 dvss 0.0603958
R23725 dvss.n4066 dvss 0.0603958
R23726 dvss.n4067 dvss 0.0603958
R23727 dvss.n4078 dvss 0.0603958
R23728 dvss.n4079 dvss 0.0603958
R23729 dvss.n4088 dvss 0.0603958
R23730 dvss.n4089 dvss 0.0603958
R23731 dvss.n4094 dvss 0.0603958
R23732 dvss dvss.n4102 0.0603958
R23733 dvss.n4103 dvss 0.0603958
R23734 dvss dvss.n4118 0.0603958
R23735 dvss.n4119 dvss 0.0603958
R23736 dvss dvss.n4032 0.0603958
R23737 dvss.n4128 dvss 0.0603958
R23738 dvss.n4190 dvss 0.0603958
R23739 dvss dvss.n4189 0.0603958
R23740 dvss dvss.n4181 0.0603958
R23741 dvss dvss.n4171 0.0603958
R23742 dvss.n4018 dvss 0.0603958
R23743 dvss dvss.n4022 0.0603958
R23744 dvss.n4270 dvss 0.0603958
R23745 dvss.n4194 dvss 0.0603958
R23746 dvss.n4264 dvss 0.0603958
R23747 dvss.n4258 dvss 0.0603958
R23748 dvss dvss.n4257 0.0603958
R23749 dvss dvss.n4256 0.0603958
R23750 dvss.n4210 dvss 0.0603958
R23751 dvss.n4225 dvss 0.0603958
R23752 dvss dvss.n4224 0.0603958
R23753 dvss.n321 dvss 0.0603958
R23754 dvss.n450 dvss 0.0603958
R23755 dvss.n6625 dvss 0.0603958
R23756 dvss.n6596 dvss 0.0603958
R23757 dvss.n6587 dvss 0.0603958
R23758 dvss.n5101 dvss.n5100 0.058075
R23759 dvss.n2656 dvss.n2408 0.0574697
R23760 dvss.n3024 dvss.n2861 0.0574697
R23761 dvss.n3438 dvss.n2667 0.0574697
R23762 dvss.n3808 dvss.n3639 0.0574697
R23763 dvss.n4004 dvss.n3450 0.0574697
R23764 dvss.n4413 dvss.n2406 0.0574697
R23765 dvss.n4709 dvss.n4708 0.0574697
R23766 dvss.n5097 dvss.n1214 0.0574697
R23767 dvss.n4153 dvss.n4008 0.0574697
R23768 dvss.n4291 dvss.n4009 0.0574697
R23769 dvss.n2548 dvss.n2409 0.0551875
R23770 dvss.n2654 dvss.n2653 0.0551875
R23771 dvss.n3015 dvss.n3014 0.0551875
R23772 dvss.n3028 dvss.n2859 0.0551875
R23773 dvss.n2816 dvss.n2668 0.0551875
R23774 dvss.n3436 dvss.n3435 0.0551875
R23775 dvss.n3790 dvss.n3789 0.0551875
R23776 dvss.n3641 dvss.n3637 0.0551875
R23777 dvss.n3475 dvss.n3474 0.0551875
R23778 dvss.n4001 dvss.n4000 0.0551875
R23779 dvss.n2403 dvss.n2398 0.0551875
R23780 dvss.n4297 dvss.n4296 0.0551875
R23781 dvss.n4713 dvss.n4712 0.0551875
R23782 dvss.n4572 dvss.n4564 0.0551875
R23783 dvss.n4924 dvss.n4919 0.0551875
R23784 dvss.n5094 dvss.n5093 0.0551875
R23785 dvss.n4171 dvss.n4170 0.0551875
R23786 dvss.n4155 dvss.n4011 0.0551875
R23787 dvss dvss.n3212 0.0477973
R23788 dvss.n6993 dvss.t655 0.047052
R23789 dvss.n6992 dvss.t658 0.047052
R23790 dvss.n6990 dvss.t659 0.047052
R23791 dvss.n6991 dvss.t656 0.047052
R23792 dvss.n7026 dvss.t288 0.047052
R23793 dvss.n7027 dvss.t294 0.047052
R23794 dvss.n7028 dvss.t290 0.047052
R23795 dvss.n7029 dvss.t293 0.047052
R23796 dvss.n7030 dvss.t289 0.047052
R23797 dvss.n3282 dvss 0.0469527
R23798 dvss.n3172 dvss 0.0469527
R23799 dvss.n5117 dvss 0.0469527
R23800 dvss.n5164 dvss 0.0469527
R23801 dvss.n5203 dvss 0.0469527
R23802 dvss.n5242 dvss 0.0469527
R23803 dvss.n5281 dvss 0.0469527
R23804 dvss.n5538 dvss 0.0469527
R23805 dvss.n6232 dvss 0.0469527
R23806 dvss dvss.n474 0.0469527
R23807 dvss.n6556 dvss 0.0469527
R23808 dvss.n6424 dvss 0.0469527
R23809 dvss.n4848 dvss.n4847 0.0466957
R23810 dvss dvss.n3217 0.0461081
R23811 dvss dvss.n3232 0.0461081
R23812 dvss.n3273 dvss 0.0435743
R23813 dvss.n3275 dvss 0.0435743
R23814 dvss.n5155 dvss 0.0435743
R23815 dvss.n5157 dvss 0.0435743
R23816 dvss.n5194 dvss 0.0435743
R23817 dvss.n5196 dvss 0.0435743
R23818 dvss.n5233 dvss 0.0435743
R23819 dvss.n5235 dvss 0.0435743
R23820 dvss.n5272 dvss 0.0435743
R23821 dvss.n5274 dvss 0.0435743
R23822 dvss.n5528 dvss 0.0435743
R23823 dvss.n5531 dvss 0.0435743
R23824 dvss.n6213 dvss 0.0435743
R23825 dvss dvss.n512 0.0435743
R23826 dvss.n6285 dvss 0.0435743
R23827 dvss dvss.n483 0.0435743
R23828 dvss dvss.n6563 0.0435743
R23829 dvss.n6352 dvss 0.0435743
R23830 dvss.n6413 dvss 0.0435743
R23831 dvss dvss.n6415 0.0435743
R23832 dvss dvss.n3441 0.0421667
R23833 dvss.n3794 dvss 0.0421667
R23834 dvss.n3805 dvss 0.0421667
R23835 dvss.n3481 dvss 0.0421667
R23836 dvss dvss.n3477 0.0421667
R23837 dvss.n3249 dvss 0.0418851
R23838 dvss.n2661 dvss.n2410 0.0410405
R23839 dvss.n2657 dvss.n2655 0.0410405
R23840 dvss.n3018 dvss.n2862 0.0410405
R23841 dvss.n3023 dvss.n2860 0.0410405
R23842 dvss.n3443 dvss.n2669 0.0410405
R23843 dvss.n3439 dvss.n3437 0.0410405
R23844 dvss.n3793 dvss.n3640 0.0410405
R23845 dvss.n3807 dvss.n3638 0.0410405
R23846 dvss.n3480 dvss.n3479 0.0410405
R23847 dvss.n4003 dvss.n4002 0.0410405
R23848 dvss.n4415 dvss.n4414 0.0410405
R23849 dvss.n4294 dvss.n4293 0.0410405
R23850 dvss.n4561 dvss.n4560 0.0410405
R23851 dvss.n4563 dvss.n4562 0.0410405
R23852 dvss.n4928 dvss.n4927 0.0410405
R23853 dvss.n5096 dvss.n5095 0.0410405
R23854 dvss.n4168 dvss.n4154 0.0410405
R23855 dvss.n4164 dvss.n4010 0.0410405
R23856 dvss.n3131 dvss 0.0410405
R23857 dvss.n5130 dvss 0.0410405
R23858 dvss dvss.n5132 0.0410405
R23859 dvss.n5169 dvss 0.0410405
R23860 dvss dvss.n5171 0.0410405
R23861 dvss.n5208 dvss 0.0410405
R23862 dvss dvss.n5210 0.0410405
R23863 dvss.n5247 dvss 0.0410405
R23864 dvss dvss.n5249 0.0410405
R23865 dvss dvss.n5285 0.0410405
R23866 dvss dvss.n1148 0.0410405
R23867 dvss.n5548 dvss 0.0410405
R23868 dvss dvss.n5552 0.0410405
R23869 dvss dvss.n6246 0.0410405
R23870 dvss dvss.n499 0.0410405
R23871 dvss.n6331 dvss 0.0410405
R23872 dvss.n6326 dvss 0.0410405
R23873 dvss.n6368 dvss 0.0410405
R23874 dvss dvss.n6372 0.0410405
R23875 dvss.n5122 dvss 0.0385068
R23876 dvss.n7048 dvss.n7047 0.0362143
R23877 dvss.n5128 dvss 0.0351284
R23878 dvss.n3420 dvss 0.0343542
R23879 dvss dvss.n3673 0.0343542
R23880 dvss.n3715 dvss 0.0343542
R23881 dvss.n3880 dvss 0.0343542
R23882 dvss.n3865 dvss 0.0343542
R23883 dvss.n3542 dvss 0.0343542
R23884 dvss.n3967 dvss 0.0343542
R23885 dvss.n4450 dvss 0.0343542
R23886 dvss dvss.n4336 0.0343542
R23887 dvss.n4505 dvss 0.0343542
R23888 dvss.n4954 dvss 0.0343542
R23889 dvss.n5059 dvss 0.0343542
R23890 dvss dvss.n4066 0.0343542
R23891 dvss.n4223 dvss 0.0343542
R23892 dvss.n2481 dvss 0.0330521
R23893 dvss dvss.n2532 0.0330521
R23894 dvss.n2629 dvss 0.0330521
R23895 dvss dvss.n2912 0.0330521
R23896 dvss dvss.n2991 0.0330521
R23897 dvss.n3122 dvss 0.0330521
R23898 dvss dvss.n2744 0.0330521
R23899 dvss dvss.n2804 0.0330521
R23900 dvss dvss.n3339 0.0330521
R23901 dvss.n3757 dvss 0.0330521
R23902 dvss dvss.n3762 0.0330521
R23903 dvss dvss.n3838 0.0330521
R23904 dvss dvss.n3568 0.0330521
R23905 dvss.n3505 dvss 0.0330521
R23906 dvss.n3976 dvss 0.0330521
R23907 dvss dvss.n2362 0.0330521
R23908 dvss.n4441 dvss 0.0330521
R23909 dvss.n4383 dvss 0.0330521
R23910 dvss.n4787 dvss 0.0330521
R23911 dvss dvss.n4544 0.0330521
R23912 dvss dvss.n4893 0.0330521
R23913 dvss.n4953 dvss 0.0330521
R23914 dvss.n5072 dvss 0.0330521
R23915 dvss.n4190 dvss 0.0330521
R23916 dvss dvss.n4194 0.0330521
R23917 dvss dvss.n7056 0.0323548
R23918 dvss.n7053 dvss 0.0323548
R23919 dvss.n2286 dvss 0.0323548
R23920 dvss dvss.n2285 0.0323548
R23921 dvss dvss.n2284 0.0323548
R23922 dvss dvss.n2277 0.0323548
R23923 dvss.n2274 dvss 0.0323548
R23924 dvss dvss.n2269 0.0323548
R23925 dvss.n2266 dvss 0.0323548
R23926 dvss.n2259 dvss 0.0323548
R23927 dvss dvss.n2257 0.0323548
R23928 dvss.n2254 dvss 0.0323548
R23929 dvss dvss.n2253 0.0323548
R23930 dvss.n2245 dvss 0.0323548
R23931 dvss.n2236 dvss 0.0323548
R23932 dvss.n2228 dvss 0.0323548
R23933 dvss dvss.n2227 0.0323548
R23934 dvss.n2218 dvss 0.0323548
R23935 dvss dvss.n2217 0.0323548
R23936 dvss dvss.n2216 0.0323548
R23937 dvss.n2213 dvss 0.0323548
R23938 dvss dvss.n2212 0.0323548
R23939 dvss dvss.n2211 0.0323548
R23940 dvss dvss.n2207 0.0323548
R23941 dvss dvss.n2206 0.0323548
R23942 dvss.n2203 dvss 0.0323548
R23943 dvss.n2195 dvss 0.0323548
R23944 dvss.n2186 dvss 0.0323548
R23945 dvss.n2178 dvss 0.0323548
R23946 dvss dvss.n2177 0.0323548
R23947 dvss.n2168 dvss 0.0323548
R23948 dvss dvss.n2161 0.0323548
R23949 dvss.n2158 dvss 0.0323548
R23950 dvss dvss.n2157 0.0323548
R23951 dvss dvss.n2156 0.0323548
R23952 dvss dvss.n2152 0.0323548
R23953 dvss dvss.n2151 0.0323548
R23954 dvss.n2148 dvss 0.0323548
R23955 dvss.n2140 dvss 0.0323548
R23956 dvss.n2131 dvss 0.0323548
R23957 dvss.n2123 dvss 0.0323548
R23958 dvss dvss.n2122 0.0323548
R23959 dvss dvss.n1344 0.0323548
R23960 dvss.n5737 dvss 0.0323548
R23961 dvss.n5748 dvss 0.0323548
R23962 dvss dvss.n5747 0.0323548
R23963 dvss dvss.n5746 0.0323548
R23964 dvss dvss.n5742 0.0323548
R23965 dvss.n5757 dvss 0.0323548
R23966 dvss.n5758 dvss 0.0323548
R23967 dvss.n5772 dvss 0.0323548
R23968 dvss dvss.n5781 0.0323548
R23969 dvss.n5796 dvss 0.0323548
R23970 dvss dvss.n5795 0.0323548
R23971 dvss.n5817 dvss 0.0323548
R23972 dvss.n5827 dvss 0.0323548
R23973 dvss.n5828 dvss 0.0323548
R23974 dvss.n5830 dvss 0.0323548
R23975 dvss dvss.n5829 0.0323548
R23976 dvss.n5839 dvss 0.0323548
R23977 dvss.n5842 dvss 0.0323548
R23978 dvss dvss.n5841 0.0323548
R23979 dvss.n5857 dvss 0.0323548
R23980 dvss dvss.n829 0.0323548
R23981 dvss.n5881 dvss 0.0323548
R23982 dvss.n5882 dvss 0.0323548
R23983 dvss.n5895 dvss 0.0323548
R23984 dvss.n6115 dvss 0.0323548
R23985 dvss dvss.n6114 0.0323548
R23986 dvss dvss.n6113 0.0323548
R23987 dvss.n6110 dvss 0.0323548
R23988 dvss dvss.n6108 0.0323548
R23989 dvss.n6105 dvss 0.0323548
R23990 dvss dvss.n6104 0.0323548
R23991 dvss.n6096 dvss 0.0323548
R23992 dvss.n6087 dvss 0.0323548
R23993 dvss.n6079 dvss 0.0323548
R23994 dvss dvss.n6078 0.0323548
R23995 dvss.n6069 dvss 0.0323548
R23996 dvss dvss.n6068 0.0323548
R23997 dvss dvss.n6067 0.0323548
R23998 dvss.n6064 dvss 0.0323548
R23999 dvss dvss.n6063 0.0323548
R24000 dvss dvss.n6062 0.0323548
R24001 dvss dvss.n6058 0.0323548
R24002 dvss dvss.n6057 0.0323548
R24003 dvss.n6054 dvss 0.0323548
R24004 dvss.n6046 dvss 0.0323548
R24005 dvss.n6037 dvss 0.0323548
R24006 dvss.n6029 dvss 0.0323548
R24007 dvss dvss.n6028 0.0323548
R24008 dvss.n6019 dvss 0.0323548
R24009 dvss dvss.n6018 0.0323548
R24010 dvss.n6721 dvss 0.0323548
R24011 dvss.n6722 dvss 0.0323548
R24012 dvss.n6724 dvss 0.0323548
R24013 dvss dvss.n6723 0.0323548
R24014 dvss.n6733 dvss 0.0323548
R24015 dvss.n6736 dvss 0.0323548
R24016 dvss dvss.n6735 0.0323548
R24017 dvss.n6751 dvss 0.0323548
R24018 dvss dvss.n100 0.0323548
R24019 dvss.n6775 dvss 0.0323548
R24020 dvss.n6776 dvss 0.0323548
R24021 dvss.n6789 dvss 0.0323548
R24022 dvss.n6790 dvss 0.0323548
R24023 dvss.n6856 dvss 0.0323548
R24024 dvss dvss.n6855 0.0323548
R24025 dvss dvss.n6854 0.0323548
R24026 dvss.n6851 dvss 0.0323548
R24027 dvss dvss.n6849 0.0323548
R24028 dvss.n6846 dvss 0.0323548
R24029 dvss dvss.n6845 0.0323548
R24030 dvss.n6837 dvss 0.0323548
R24031 dvss.n6828 dvss 0.0323548
R24032 dvss.n6955 dvss 0.0323548
R24033 dvss.n6964 dvss 0.0323548
R24034 dvss.n6973 dvss 0.0323548
R24035 dvss.n6977 dvss 0.0323548
R24036 dvss dvss.n6976 0.0323548
R24037 dvss dvss.n6975 0.0323548
R24038 dvss dvss.n6974 0.0323548
R24039 dvss.n6988 dvss 0.0323548
R24040 dvss dvss.n2235 0.0319516
R24041 dvss dvss.n2185 0.0319516
R24042 dvss dvss.n2130 0.0319516
R24043 dvss.n5791 dvss 0.0319516
R24044 dvss dvss.n825 0.0319516
R24045 dvss dvss.n6086 0.0319516
R24046 dvss dvss.n6036 0.0319516
R24047 dvss dvss.n96 0.0319516
R24048 dvss dvss.n6827 0.0319516
R24049 dvss.n2459 dvss 0.03175
R24050 dvss.n2562 dvss 0.03175
R24051 dvss.n2628 dvss 0.03175
R24052 dvss.n2883 dvss 0.03175
R24053 dvss.n2985 dvss 0.03175
R24054 dvss.n3008 dvss 0.03175
R24055 dvss dvss.n3049 0.03175
R24056 dvss dvss.n2720 0.03175
R24057 dvss.n2842 dvss 0.03175
R24058 dvss.n2828 dvss 0.03175
R24059 dvss.n3421 dvss 0.03175
R24060 dvss.n3370 dvss 0.03175
R24061 dvss.n3756 dvss 0.03175
R24062 dvss dvss.n3763 0.03175
R24063 dvss.n3804 dvss 0.03175
R24064 dvss dvss.n3583 0.03175
R24065 dvss.n3504 dvss 0.03175
R24066 dvss.n3975 dvss 0.03175
R24067 dvss.n2339 dvss 0.03175
R24068 dvss.n4396 dvss 0.03175
R24069 dvss dvss.n4504 0.03175
R24070 dvss.n4666 dvss 0.03175
R24071 dvss.n4652 dvss 0.03175
R24072 dvss.n4871 dvss 0.03175
R24073 dvss.n5079 dvss 0.03175
R24074 dvss.n5038 dvss 0.03175
R24075 dvss.n4063 dvss 0.03175
R24076 dvss.n4257 dvss 0.03175
R24077 dvss.n5736 dvss.n884 0.0311452
R24078 dvss.n5816 dvss.n5811 0.0311452
R24079 dvss.n5901 dvss.n5900 0.0311452
R24080 dvss dvss.n3270 0.0300608
R24081 dvss dvss.n5147 0.0300608
R24082 dvss dvss.n5186 0.0300608
R24083 dvss dvss.n5225 0.0300608
R24084 dvss dvss.n5264 0.0300608
R24085 dvss dvss.n1127 0.0300608
R24086 dvss.n6217 dvss 0.0300608
R24087 dvss dvss.n6286 0.0300608
R24088 dvss dvss.n231 0.0300608
R24089 dvss dvss.n6397 0.0300608
R24090 dvss.n2167 dvss.n2162 0.0295323
R24091 dvss.n7025 dvss.n7024 0.029472
R24092 dvss.n7037 dvss.n7033 0.029472
R24093 dvss.n3450 dvss.n3448 0.0292489
R24094 dvss.n4005 dvss.n4004 0.0292489
R24095 dvss.n1214 dvss.n1212 0.0292489
R24096 dvss.n5098 dvss.n5097 0.0292489
R24097 dvss.n4710 dvss.n4709 0.0292489
R24098 dvss.n4708 dvss.n4707 0.0292489
R24099 dvss.n4413 dvss.n4412 0.0292489
R24100 dvss.n4410 dvss.n2406 0.0292489
R24101 dvss.n3791 dvss.n3639 0.0292489
R24102 dvss.n3809 dvss.n3808 0.0292489
R24103 dvss.n3445 dvss.n2667 0.0292489
R24104 dvss.n3438 dvss.n2666 0.0292489
R24105 dvss.n3016 dvss.n2861 0.0292489
R24106 dvss.n3025 dvss.n3024 0.0292489
R24107 dvss.n2663 dvss.n2408 0.0292489
R24108 dvss.n2656 dvss.n2407 0.0292489
R24109 dvss.n4009 dvss.n4007 0.0292489
R24110 dvss.n4153 dvss.n4007 0.0292489
R24111 dvss.n2653 dvss.n2414 0.0291458
R24112 dvss.n3028 dvss.n3027 0.0291458
R24113 dvss.n3435 dvss.n2673 0.0291458
R24114 dvss.n3811 dvss.n3637 0.0291458
R24115 dvss.n4000 dvss.n3452 0.0291458
R24116 dvss.n4408 dvss.n4297 0.0291458
R24117 dvss.n4705 dvss.n4564 0.0291458
R24118 dvss dvss.n4589 0.0291458
R24119 dvss.n5093 dvss.n1217 0.0291458
R24120 dvss dvss.n1221 0.0291458
R24121 dvss dvss.n5016 0.0291458
R24122 dvss.n4289 dvss.n4011 0.0291458
R24123 dvss.n1246 dvss 0.0287258
R24124 dvss.n1777 dvss 0.0282388
R24125 dvss.n1803 dvss 0.0282388
R24126 dvss.n1823 dvss 0.0282388
R24127 dvss.n1845 dvss 0.0282388
R24128 dvss dvss.n1856 0.0282388
R24129 dvss.n1866 dvss 0.0282388
R24130 dvss dvss.n1869 0.0282388
R24131 dvss.n1884 dvss 0.0282388
R24132 dvss dvss.n1883 0.0282388
R24133 dvss.n1892 dvss 0.0282388
R24134 dvss.n1918 dvss 0.0282388
R24135 dvss.n1937 dvss 0.0282388
R24136 dvss dvss.n1977 0.0282388
R24137 dvss.n1964 dvss 0.0282388
R24138 dvss.n2052 dvss 0.0282388
R24139 dvss.n2049 dvss 0.0282388
R24140 dvss dvss.n2048 0.0282388
R24141 dvss dvss.n2040 0.0282388
R24142 dvss.n2079 dvss 0.0282388
R24143 dvss dvss.n1413 0.0282388
R24144 dvss.n1384 dvss 0.0282388
R24145 dvss.n1399 dvss 0.0282388
R24146 dvss.n5724 dvss 0.0282388
R24147 dvss dvss.n5723 0.0282388
R24148 dvss dvss.n5722 0.0282388
R24149 dvss dvss.n5718 0.0282388
R24150 dvss.n996 dvss 0.0282388
R24151 dvss dvss.n5701 0.0282388
R24152 dvss dvss.n5690 0.0282388
R24153 dvss dvss.n987 0.0282388
R24154 dvss.n5675 dvss 0.0282388
R24155 dvss dvss.n5674 0.0282388
R24156 dvss dvss.n5673 0.0282388
R24157 dvss dvss.n956 0.0282388
R24158 dvss.n1091 dvss 0.0282388
R24159 dvss.n5648 dvss 0.0282388
R24160 dvss.n5637 dvss 0.0282388
R24161 dvss.n5624 dvss 0.0282388
R24162 dvss.n6155 dvss 0.0282388
R24163 dvss.n6152 dvss 0.0282388
R24164 dvss dvss.n6151 0.0282388
R24165 dvss dvss.n6143 0.0282388
R24166 dvss.n6182 dvss 0.0282388
R24167 dvss dvss.n763 0.0282388
R24168 dvss.n636 dvss 0.0282388
R24169 dvss dvss.n618 0.0282388
R24170 dvss dvss.n617 0.0282388
R24171 dvss.n752 dvss 0.0282388
R24172 dvss dvss.n751 0.0282388
R24173 dvss dvss.n750 0.0282388
R24174 dvss dvss.n746 0.0282388
R24175 dvss.n604 dvss 0.0282388
R24176 dvss dvss.n729 0.0282388
R24177 dvss dvss.n718 0.0282388
R24178 dvss.n705 dvss 0.0282388
R24179 dvss.n706 dvss 0.0282388
R24180 dvss.n6708 dvss 0.0282388
R24181 dvss dvss.n6707 0.0282388
R24182 dvss dvss.n6706 0.0282388
R24183 dvss dvss.n6702 0.0282388
R24184 dvss.n213 dvss 0.0282388
R24185 dvss dvss.n6685 0.0282388
R24186 dvss dvss.n6674 0.0282388
R24187 dvss.n6661 dvss 0.0282388
R24188 dvss.n6865 dvss 0.0282388
R24189 dvss.n6896 dvss 0.0282388
R24190 dvss.n6893 dvss 0.0282388
R24191 dvss dvss.n6892 0.0282388
R24192 dvss dvss.n6884 0.0282388
R24193 dvss.n6923 dvss 0.0282388
R24194 dvss dvss.n39 0.0282388
R24195 dvss.n6463 dvss 0.0282388
R24196 dvss.n6476 dvss 0.0282388
R24197 dvss.n6483 dvss 0.0282388
R24198 dvss.n6494 dvss 0.0282388
R24199 dvss.n6495 dvss 0.0282388
R24200 dvss.n6498 dvss 0.0282388
R24201 dvss.n1700 dvss 0.0278876
R24202 dvss dvss.n1600 0.0278876
R24203 dvss dvss.n1601 0.0278876
R24204 dvss dvss.n1602 0.0278876
R24205 dvss dvss.n1603 0.0278876
R24206 dvss dvss.n1606 0.0278876
R24207 dvss dvss.n1607 0.0278876
R24208 dvss.n1620 dvss 0.0278876
R24209 dvss.n1758 dvss 0.0278876
R24210 dvss.n1585 dvss 0.0278876
R24211 dvss.n1827 dvss 0.0278876
R24212 dvss.n1939 dvss 0.0278876
R24213 dvss dvss.n1355 0.0278876
R24214 dvss dvss.n5700 0.0278876
R24215 dvss.n1081 dvss 0.0278876
R24216 dvss dvss.n532 0.0278876
R24217 dvss dvss.n728 0.0278876
R24218 dvss dvss.n6684 0.0278876
R24219 dvss dvss.n30 0.0278876
R24220 dvss.n3211 dvss 0.027527
R24221 dvss dvss.n3227 0.027527
R24222 dvss.n2021 dvss.n1453 0.0271854
R24223 dvss.n1405 dvss.n1404 0.0271854
R24224 dvss.n986 dvss.n981 0.0271854
R24225 dvss.n6124 dvss.n803 0.0271854
R24226 dvss dvss.n3201 0.0258378
R24227 dvss.n3228 dvss 0.0258378
R24228 dvss.n1789 dvss 0.0257809
R24229 dvss.n1898 dvss 0.0257809
R24230 dvss.n2064 dvss 0.0257809
R24231 dvss dvss.n5714 0.0257809
R24232 dvss.n963 dvss 0.0257809
R24233 dvss.n6167 dvss 0.0257809
R24234 dvss dvss.n742 0.0257809
R24235 dvss dvss.n6698 0.0257809
R24236 dvss.n6908 dvss 0.0257809
R24237 dvss.n1709 dvss 0.0247275
R24238 dvss dvss.n2992 0.0239375
R24239 dvss dvss.n2807 0.0239375
R24240 dvss.n2834 dvss 0.0239375
R24241 dvss dvss.n3341 0.0239375
R24242 dvss.n3674 dvss 0.0239375
R24243 dvss.n3626 dvss 0.0239375
R24244 dvss.n4747 dvss 0.0239375
R24245 dvss.n4729 dvss 0.0239375
R24246 dvss.n4045 dvss 0.0239375
R24247 dvss.n4264 dvss 0.0239375
R24248 dvss dvss.n1701 0.0236742
R24249 dvss.n3271 dvss 0.0233041
R24250 dvss.n5153 dvss 0.0233041
R24251 dvss.n5192 dvss 0.0233041
R24252 dvss.n5231 dvss 0.0233041
R24253 dvss.n5270 dvss 0.0233041
R24254 dvss dvss.n1136 0.0233041
R24255 dvss.n6215 dvss 0.0233041
R24256 dvss dvss.n6287 0.0233041
R24257 dvss.n6560 dvss 0.0233041
R24258 dvss.n6411 dvss 0.0233041
R24259 dvss dvss.n2248 0.0230806
R24260 dvss dvss.n2198 0.0230806
R24261 dvss dvss.n2143 0.0230806
R24262 dvss dvss.n871 0.0230806
R24263 dvss dvss.n5851 0.0230806
R24264 dvss dvss.n6099 0.0230806
R24265 dvss dvss.n6049 0.0230806
R24266 dvss dvss.n6745 0.0230806
R24267 dvss dvss.n6840 0.0230806
R24268 dvss.n2271 dvss 0.0226774
R24269 dvss dvss.n2222 0.0226774
R24270 dvss dvss.n2172 0.0226774
R24271 dvss dvss.n2117 0.0226774
R24272 dvss.n5809 dvss 0.0226774
R24273 dvss.n819 dvss 0.0226774
R24274 dvss dvss.n6073 0.0226774
R24275 dvss dvss.n6023 0.0226774
R24276 dvss.n90 dvss 0.0226774
R24277 dvss dvss.n6959 0.0226774
R24278 dvss dvss.n2480 0.0226354
R24279 dvss.n2489 dvss 0.0226354
R24280 dvss.n2504 dvss 0.0226354
R24281 dvss dvss.n2525 0.0226354
R24282 dvss.n2526 dvss 0.0226354
R24283 dvss.n2561 dvss 0.0226354
R24284 dvss.n2555 dvss 0.0226354
R24285 dvss.n2550 dvss 0.0226354
R24286 dvss.n2644 dvss 0.0226354
R24287 dvss.n2632 dvss 0.0226354
R24288 dvss.n2613 dvss 0.0226354
R24289 dvss.n2591 dvss 0.0226354
R24290 dvss.n2900 dvss 0.0226354
R24291 dvss dvss.n2911 0.0226354
R24292 dvss.n2978 dvss 0.0226354
R24293 dvss dvss.n2921 0.0226354
R24294 dvss.n2934 dvss 0.0226354
R24295 dvss dvss.n3006 0.0226354
R24296 dvss dvss.n3032 0.0226354
R24297 dvss dvss.n3052 0.0226354
R24298 dvss.n3104 dvss 0.0226354
R24299 dvss dvss.n3061 0.0226354
R24300 dvss.n3096 dvss 0.0226354
R24301 dvss.n3078 dvss 0.0226354
R24302 dvss dvss.n2727 0.0226354
R24303 dvss dvss.n2728 0.0226354
R24304 dvss.n2752 dvss 0.0226354
R24305 dvss.n2776 dvss 0.0226354
R24306 dvss dvss.n2782 0.0226354
R24307 dvss dvss.n2793 0.0226354
R24308 dvss dvss.n2814 0.0226354
R24309 dvss.n3431 dvss 0.0226354
R24310 dvss.n3428 dvss 0.0226354
R24311 dvss.n3427 dvss 0.0226354
R24312 dvss.n3414 dvss 0.0226354
R24313 dvss.n3410 dvss 0.0226354
R24314 dvss dvss.n3347 0.0226354
R24315 dvss dvss.n3349 0.0226354
R24316 dvss.n3377 dvss 0.0226354
R24317 dvss.n3376 dvss 0.0226354
R24318 dvss dvss.n3359 0.0226354
R24319 dvss dvss.n3672 0.0226354
R24320 dvss dvss.n3695 0.0226354
R24321 dvss.n3719 dvss 0.0226354
R24322 dvss.n3718 dvss 0.0226354
R24323 dvss.n3709 dvss 0.0226354
R24324 dvss dvss.n3837 0.0226354
R24325 dvss.n3895 dvss 0.0226354
R24326 dvss dvss.n3847 0.0226354
R24327 dvss.n3867 dvss 0.0226354
R24328 dvss.n3547 dvss 0.0226354
R24329 dvss dvss.n3550 0.0226354
R24330 dvss.n3551 dvss 0.0226354
R24331 dvss dvss.n3555 0.0226354
R24332 dvss.n3565 dvss 0.0226354
R24333 dvss.n3576 dvss 0.0226354
R24334 dvss.n3584 dvss 0.0226354
R24335 dvss dvss.n3589 0.0226354
R24336 dvss dvss.n3609 0.0226354
R24337 dvss.n3610 dvss 0.0226354
R24338 dvss dvss.n3625 0.0226354
R24339 dvss.n3500 dvss 0.0226354
R24340 dvss.n3493 dvss 0.0226354
R24341 dvss.n3476 dvss 0.0226354
R24342 dvss.n3935 dvss 0.0226354
R24343 dvss.n3934 dvss 0.0226354
R24344 dvss.n3929 dvss 0.0226354
R24345 dvss dvss.n2361 0.0226354
R24346 dvss dvss.n2369 0.0226354
R24347 dvss.n4454 dvss 0.0226354
R24348 dvss.n4449 dvss 0.0226354
R24349 dvss.n4434 dvss 0.0226354
R24350 dvss.n4431 dvss 0.0226354
R24351 dvss.n4402 dvss 0.0226354
R24352 dvss.n4397 dvss 0.0226354
R24353 dvss.n4388 dvss 0.0226354
R24354 dvss.n4387 dvss 0.0226354
R24355 dvss dvss.n4318 0.0226354
R24356 dvss.n4358 dvss 0.0226354
R24357 dvss.n4350 dvss 0.0226354
R24358 dvss.n4345 dvss 0.0226354
R24359 dvss dvss.n4523 0.0226354
R24360 dvss dvss.n4524 0.0226354
R24361 dvss.n4773 dvss 0.0226354
R24362 dvss dvss.n4533 0.0226354
R24363 dvss.n4751 dvss 0.0226354
R24364 dvss.n4738 dvss 0.0226354
R24365 dvss dvss.n4548 0.0226354
R24366 dvss dvss.n4555 0.0226354
R24367 dvss.n4704 dvss 0.0226354
R24368 dvss dvss.n4581 0.0226354
R24369 dvss.n4679 dvss 0.0226354
R24370 dvss dvss.n4594 0.0226354
R24371 dvss.n4675 dvss 0.0226354
R24372 dvss dvss.n4612 0.0226354
R24373 dvss.n4659 dvss 0.0226354
R24374 dvss.n4644 dvss 0.0226354
R24375 dvss dvss.n4621 0.0226354
R24376 dvss.n4634 dvss 0.0226354
R24377 dvss dvss.n4624 0.0226354
R24378 dvss dvss.n4892 0.0226354
R24379 dvss.n4997 dvss 0.0226354
R24380 dvss dvss.n4898 0.0226354
R24381 dvss.n4984 dvss 0.0226354
R24382 dvss dvss.n4903 0.0226354
R24383 dvss.n4971 dvss 0.0226354
R24384 dvss dvss.n4908 0.0226354
R24385 dvss.n4958 dvss 0.0226354
R24386 dvss.n4946 dvss 0.0226354
R24387 dvss dvss.n4917 0.0226354
R24388 dvss.n5085 dvss 0.0226354
R24389 dvss.n5073 dvss 0.0226354
R24390 dvss dvss.n5008 0.0226354
R24391 dvss.n5025 dvss 0.0226354
R24392 dvss.n4075 dvss 0.0226354
R24393 dvss dvss.n4078 0.0226354
R24394 dvss dvss.n4088 0.0226354
R24395 dvss.n4089 dvss 0.0226354
R24396 dvss dvss.n4103 0.0226354
R24397 dvss.n4033 dvss 0.0226354
R24398 dvss dvss.n4127 0.0226354
R24399 dvss dvss.n4137 0.0226354
R24400 dvss.n4182 dvss 0.0226354
R24401 dvss.n4181 dvss 0.0226354
R24402 dvss.n4172 dvss 0.0226354
R24403 dvss.n4282 dvss 0.0226354
R24404 dvss.n4256 dvss 0.0226354
R24405 dvss.n4238 dvss 0.0226354
R24406 dvss dvss.n4210 0.0226354
R24407 dvss.n324 dvss 0.0226354
R24408 dvss.n315 dvss 0.0226354
R24409 dvss.n446 dvss 0.0226354
R24410 dvss dvss.n456 0.0226354
R24411 dvss.n6621 dvss 0.0226354
R24412 dvss dvss.n6631 0.0226354
R24413 dvss.n6599 dvss 0.0226354
R24414 dvss.n6590 dvss 0.0226354
R24415 dvss.n6581 dvss 0.0226354
R24416 dvss dvss.n2244 0.0222742
R24417 dvss.n2232 dvss 0.0222742
R24418 dvss dvss.n2194 0.0222742
R24419 dvss.n2182 dvss 0.0222742
R24420 dvss dvss.n2139 0.0222742
R24421 dvss.n2127 dvss 0.0222742
R24422 dvss.n5774 dvss 0.0222742
R24423 dvss.n5793 dvss 0.0222742
R24424 dvss dvss.n5856 0.0222742
R24425 dvss dvss.n5871 0.0222742
R24426 dvss dvss.n6095 0.0222742
R24427 dvss.n6083 dvss 0.0222742
R24428 dvss dvss.n6045 0.0222742
R24429 dvss.n6033 dvss 0.0222742
R24430 dvss dvss.n6750 0.0222742
R24431 dvss dvss.n6765 0.0222742
R24432 dvss dvss.n6836 0.0222742
R24433 dvss.n6824 dvss 0.0222742
R24434 dvss dvss.n2531 0.0213333
R24435 dvss dvss.n2417 0.0213333
R24436 dvss dvss.n2422 0.0213333
R24437 dvss.n3033 dvss 0.0213333
R24438 dvss dvss.n3048 0.0213333
R24439 dvss dvss.n2733 0.0213333
R24440 dvss dvss.n2738 0.0213333
R24441 dvss.n3821 dvss 0.0213333
R24442 dvss dvss.n3842 0.0213333
R24443 dvss dvss.n3614 0.0213333
R24444 dvss.n3498 dvss 0.0213333
R24445 dvss dvss.n3456 0.0213333
R24446 dvss dvss.n3463 0.0213333
R24447 dvss dvss.n3909 0.0213333
R24448 dvss dvss.n4553 0.0213333
R24449 dvss.n4573 dvss 0.0213333
R24450 dvss.n4268 dvss 0.0213333
R24451 dvss.n1281 dvss 0.0202581
R24452 dvss.n1312 dvss 0.0202581
R24453 dvss.n1343 dvss 0.0202581
R24454 dvss.n5804 dvss 0.0202581
R24455 dvss.n5887 dvss 0.0202581
R24456 dvss.n5942 dvss 0.0202581
R24457 dvss.n5973 dvss 0.0202581
R24458 dvss.n6781 dvss 0.0202581
R24459 dvss.n6958 dvss 0.0202581
R24460 dvss.n1800 dvss 0.0201629
R24461 dvss.n1911 dvss 0.0201629
R24462 dvss dvss.n2073 0.0201629
R24463 dvss.n995 dvss 0.0201629
R24464 dvss dvss.n1065 0.0201629
R24465 dvss dvss.n6176 0.0201629
R24466 dvss.n603 dvss 0.0201629
R24467 dvss.n212 dvss 0.0201629
R24468 dvss dvss.n6917 0.0201629
R24469 dvss.n4353 dvss 0.0200312
R24470 dvss.n2208 dvss 0.0198548
R24471 dvss.n2153 dvss 0.0198548
R24472 dvss.n5743 dvss 0.0198548
R24473 dvss.n5838 dvss 0.0198548
R24474 dvss dvss.n6109 0.0198548
R24475 dvss.n6059 dvss 0.0198548
R24476 dvss.n6732 dvss 0.0198548
R24477 dvss dvss.n6850 0.0198548
R24478 dvss dvss.n1509 0.0198118
R24479 dvss.n2024 dvss 0.0198118
R24480 dvss dvss.n895 0.0198118
R24481 dvss.n5679 dvss 0.0198118
R24482 dvss.n6127 dvss 0.0198118
R24483 dvss.n756 dvss 0.0198118
R24484 dvss dvss.n129 0.0198118
R24485 dvss.n6868 dvss 0.0198118
R24486 dvss.n6486 dvss 0.0198118
R24487 dvss.n1804 dvss 0.0194607
R24488 dvss.n1919 dvss 0.0194607
R24489 dvss dvss.n2078 0.0194607
R24490 dvss.n5706 dvss 0.0194607
R24491 dvss.n1092 dvss 0.0194607
R24492 dvss dvss.n6181 0.0194607
R24493 dvss.n734 dvss 0.0194607
R24494 dvss.n6690 dvss 0.0194607
R24495 dvss dvss.n6922 0.0194607
R24496 dvss.n7052 dvss.n4 0.0194516
R24497 dvss dvss.n2258 0.0194516
R24498 dvss dvss.n2280 0.0190484
R24499 dvss.n2660 dvss.n2411 0.0187292
R24500 dvss.n2659 dvss.n2412 0.0187292
R24501 dvss.n3019 dvss.n2863 0.0187292
R24502 dvss.n3021 dvss.n3020 0.0187292
R24503 dvss.n3442 dvss.n2670 0.0187292
R24504 dvss.n3441 dvss.n2671 0.0187292
R24505 dvss.n3795 dvss.n3794 0.0187292
R24506 dvss.n3805 dvss.n3804 0.0187292
R24507 dvss.n3482 dvss.n3481 0.0187292
R24508 dvss.n3477 dvss.n3476 0.0187292
R24509 dvss.n4417 dvss.n4416 0.0187292
R24510 dvss.n4295 dvss.n2402 0.0187292
R24511 dvss.n4569 dvss.n4559 0.0187292
R24512 dvss.n4573 dvss.n4571 0.0187292
R24513 dvss.n4930 dvss.n4929 0.0187292
R24514 dvss.n4925 dvss.n1216 0.0187292
R24515 dvss.n4167 dvss.n4152 0.0187292
R24516 dvss.n4166 dvss.n4163 0.0187292
R24517 dvss dvss.n2265 0.0186452
R24518 dvss dvss.n1533 0.0184073
R24519 dvss.n1942 dvss 0.0184073
R24520 dvss.n2095 dvss 0.0184073
R24521 dvss.n928 dvss 0.0184073
R24522 dvss dvss.n5644 0.0184073
R24523 dvss.n6198 dvss 0.0184073
R24524 dvss.n574 dvss 0.0184073
R24525 dvss.n162 dvss 0.0184073
R24526 dvss.n6939 dvss 0.0184073
R24527 dvss.n5127 dvss 0.0182365
R24528 dvss dvss.n1553 0.0173539
R24529 dvss dvss.n1882 0.0173539
R24530 dvss dvss.n1487 0.0173539
R24531 dvss dvss.n2047 0.0173539
R24532 dvss.n2061 dvss 0.0173539
R24533 dvss.n5719 dvss 0.0173539
R24534 dvss.n908 dvss 0.0173539
R24535 dvss.n968 dvss 0.0173539
R24536 dvss dvss.n957 0.0173539
R24537 dvss dvss.n6150 0.0173539
R24538 dvss.n6164 dvss 0.0173539
R24539 dvss.n747 dvss 0.0173539
R24540 dvss.n554 dvss 0.0173539
R24541 dvss.n6703 dvss 0.0173539
R24542 dvss.n142 dvss 0.0173539
R24543 dvss dvss.n6891 0.0173539
R24544 dvss.n6905 dvss 0.0173539
R24545 dvss dvss.n2262 0.0170323
R24546 dvss.n1588 dvss 0.0170028
R24547 dvss.n4816 dvss.n4815 0.0168445
R24548 dvss.n4828 dvss.n4827 0.0168445
R24549 dvss dvss.n1608 0.0166517
R24550 dvss dvss.n1711 0.0163006
R24551 dvss.n1861 dvss 0.0163006
R24552 dvss dvss.n1514 0.0163006
R24553 dvss.n1970 dvss 0.0163006
R24554 dvss dvss.n1972 0.0163006
R24555 dvss dvss.n1369 0.0163006
R24556 dvss.n1372 dvss 0.0163006
R24557 dvss.n5683 dvss 0.0163006
R24558 dvss dvss.n5685 0.0163006
R24559 dvss.n5630 dvss 0.0163006
R24560 dvss dvss.n5632 0.0163006
R24561 dvss dvss.n621 0.0163006
R24562 dvss.n623 dvss 0.0163006
R24563 dvss.n711 dvss 0.0163006
R24564 dvss dvss.n713 0.0163006
R24565 dvss.n6667 dvss 0.0163006
R24566 dvss dvss.n6669 0.0163006
R24567 dvss dvss.n6448 0.0163006
R24568 dvss.n6452 dvss 0.0163006
R24569 dvss.n1765 dvss 0.0159494
R24570 dvss.n4826 dvss.n1234 0.0157459
R24571 dvss.n4814 dvss.n2304 0.0157459
R24572 dvss.n3333 dvss 0.0148581
R24573 dvss.n3332 dvss 0.0148581
R24574 dvss.n3329 dvss 0.0148581
R24575 dvss dvss.n3139 0.0148581
R24576 dvss dvss.n3140 0.0148581
R24577 dvss dvss.n3141 0.0148581
R24578 dvss dvss.n3142 0.0148581
R24579 dvss dvss.n3147 0.0148581
R24580 dvss dvss.n3148 0.0148581
R24581 dvss dvss.n3149 0.0148581
R24582 dvss.n3273 dvss 0.0148581
R24583 dvss dvss.n3150 0.0148581
R24584 dvss.n3271 dvss 0.0148581
R24585 dvss.n3270 dvss 0.0148581
R24586 dvss dvss.n3155 0.0148581
R24587 dvss.n3275 dvss 0.0148581
R24588 dvss dvss.n3157 0.0148581
R24589 dvss dvss.n3268 0.0148581
R24590 dvss dvss.n3269 0.0148581
R24591 dvss.n3280 dvss 0.0148581
R24592 dvss dvss.n3284 0.0148581
R24593 dvss dvss.n3287 0.0148581
R24594 dvss.n3288 dvss 0.0148581
R24595 dvss dvss.n3200 0.0148581
R24596 dvss.n3203 dvss 0.0148581
R24597 dvss.n3202 dvss 0.0148581
R24598 dvss.n3201 dvss 0.0148581
R24599 dvss dvss.n3211 0.0148581
R24600 dvss.n3213 dvss 0.0148581
R24601 dvss.n3212 dvss 0.0148581
R24602 dvss.n3218 dvss 0.0148581
R24603 dvss.n3217 dvss 0.0148581
R24604 dvss.n3188 dvss 0.0148581
R24605 dvss.n3228 dvss 0.0148581
R24606 dvss.n3227 dvss 0.0148581
R24607 dvss.n3182 dvss 0.0148581
R24608 dvss.n3232 dvss 0.0148581
R24609 dvss.n3179 dvss 0.0148581
R24610 dvss dvss.n3243 0.0148581
R24611 dvss dvss.n3244 0.0148581
R24612 dvss.n3245 dvss 0.0148581
R24613 dvss.n3172 dvss 0.0148581
R24614 dvss.n3171 dvss 0.0148581
R24615 dvss dvss.n3257 0.0148581
R24616 dvss dvss.n3258 0.0148581
R24617 dvss.n3261 dvss 0.0148581
R24618 dvss.n3260 dvss 0.0148581
R24619 dvss.n3259 dvss 0.0148581
R24620 dvss.n6634 dvss 0.0148581
R24621 dvss dvss.n5103 0.0148581
R24622 dvss dvss.n5104 0.0148581
R24623 dvss dvss.n5105 0.0148581
R24624 dvss dvss.n5106 0.0148581
R24625 dvss dvss.n5107 0.0148581
R24626 dvss dvss.n5108 0.0148581
R24627 dvss dvss.n5109 0.0148581
R24628 dvss dvss.n5110 0.0148581
R24629 dvss dvss.n5111 0.0148581
R24630 dvss.n5112 dvss 0.0148581
R24631 dvss dvss.n5119 0.0148581
R24632 dvss dvss.n5120 0.0148581
R24633 dvss.n5122 dvss 0.0148581
R24634 dvss dvss.n5121 0.0148581
R24635 dvss dvss.n5121 0.0148581
R24636 dvss dvss.n5127 0.0148581
R24637 dvss dvss.n5128 0.0148581
R24638 dvss dvss.n5129 0.0148581
R24639 dvss dvss.n5130 0.0148581
R24640 dvss dvss.n5131 0.0148581
R24641 dvss.n5133 dvss 0.0148581
R24642 dvss dvss.n5138 0.0148581
R24643 dvss dvss.n5139 0.0148581
R24644 dvss dvss.n5140 0.0148581
R24645 dvss dvss.n5141 0.0148581
R24646 dvss dvss.n5142 0.0148581
R24647 dvss dvss.n5143 0.0148581
R24648 dvss dvss.n5144 0.0148581
R24649 dvss dvss.n5145 0.0148581
R24650 dvss.n5155 dvss 0.0148581
R24651 dvss dvss.n5146 0.0148581
R24652 dvss.n5153 dvss 0.0148581
R24653 dvss dvss.n5147 0.0148581
R24654 dvss dvss.n5148 0.0148581
R24655 dvss.n5157 dvss 0.0148581
R24656 dvss dvss.n5150 0.0148581
R24657 dvss dvss.n5151 0.0148581
R24658 dvss dvss.n5152 0.0148581
R24659 dvss.n5162 dvss 0.0148581
R24660 dvss dvss.n5166 0.0148581
R24661 dvss dvss.n5167 0.0148581
R24662 dvss dvss.n5168 0.0148581
R24663 dvss dvss.n5169 0.0148581
R24664 dvss dvss.n5170 0.0148581
R24665 dvss.n5172 dvss 0.0148581
R24666 dvss dvss.n5177 0.0148581
R24667 dvss dvss.n5178 0.0148581
R24668 dvss dvss.n5179 0.0148581
R24669 dvss dvss.n5180 0.0148581
R24670 dvss dvss.n5181 0.0148581
R24671 dvss dvss.n5182 0.0148581
R24672 dvss dvss.n5183 0.0148581
R24673 dvss dvss.n5184 0.0148581
R24674 dvss.n5194 dvss 0.0148581
R24675 dvss dvss.n5185 0.0148581
R24676 dvss.n5192 dvss 0.0148581
R24677 dvss dvss.n5186 0.0148581
R24678 dvss dvss.n5187 0.0148581
R24679 dvss.n5196 dvss 0.0148581
R24680 dvss dvss.n5189 0.0148581
R24681 dvss dvss.n5190 0.0148581
R24682 dvss dvss.n5191 0.0148581
R24683 dvss.n5201 dvss 0.0148581
R24684 dvss dvss.n5205 0.0148581
R24685 dvss dvss.n5206 0.0148581
R24686 dvss dvss.n5207 0.0148581
R24687 dvss dvss.n5208 0.0148581
R24688 dvss dvss.n5209 0.0148581
R24689 dvss.n5211 dvss 0.0148581
R24690 dvss dvss.n5216 0.0148581
R24691 dvss dvss.n5217 0.0148581
R24692 dvss dvss.n5218 0.0148581
R24693 dvss dvss.n5219 0.0148581
R24694 dvss dvss.n5220 0.0148581
R24695 dvss dvss.n5221 0.0148581
R24696 dvss dvss.n5222 0.0148581
R24697 dvss dvss.n5223 0.0148581
R24698 dvss.n5233 dvss 0.0148581
R24699 dvss dvss.n5224 0.0148581
R24700 dvss.n5231 dvss 0.0148581
R24701 dvss dvss.n5225 0.0148581
R24702 dvss dvss.n5226 0.0148581
R24703 dvss.n5235 dvss 0.0148581
R24704 dvss dvss.n5228 0.0148581
R24705 dvss dvss.n5229 0.0148581
R24706 dvss dvss.n5230 0.0148581
R24707 dvss.n5240 dvss 0.0148581
R24708 dvss dvss.n5244 0.0148581
R24709 dvss dvss.n5245 0.0148581
R24710 dvss dvss.n5246 0.0148581
R24711 dvss dvss.n5247 0.0148581
R24712 dvss dvss.n5248 0.0148581
R24713 dvss.n5250 dvss 0.0148581
R24714 dvss dvss.n5255 0.0148581
R24715 dvss dvss.n5256 0.0148581
R24716 dvss dvss.n5257 0.0148581
R24717 dvss dvss.n5258 0.0148581
R24718 dvss dvss.n5259 0.0148581
R24719 dvss dvss.n5260 0.0148581
R24720 dvss dvss.n5261 0.0148581
R24721 dvss dvss.n5262 0.0148581
R24722 dvss.n5272 dvss 0.0148581
R24723 dvss dvss.n5263 0.0148581
R24724 dvss.n5270 dvss 0.0148581
R24725 dvss dvss.n5264 0.0148581
R24726 dvss dvss.n5265 0.0148581
R24727 dvss.n5274 dvss 0.0148581
R24728 dvss dvss.n5267 0.0148581
R24729 dvss dvss.n5268 0.0148581
R24730 dvss dvss.n5269 0.0148581
R24731 dvss.n5279 dvss 0.0148581
R24732 dvss dvss.n5283 0.0148581
R24733 dvss dvss.n5284 0.0148581
R24734 dvss.n5286 dvss 0.0148581
R24735 dvss.n5285 dvss 0.0148581
R24736 dvss dvss.n5499 0.0148581
R24737 dvss.n5500 dvss 0.0148581
R24738 dvss dvss.n5505 0.0148581
R24739 dvss.n5507 dvss 0.0148581
R24740 dvss.n5506 dvss 0.0148581
R24741 dvss dvss.n5515 0.0148581
R24742 dvss dvss.n5516 0.0148581
R24743 dvss.n5518 dvss 0.0148581
R24744 dvss.n5517 dvss 0.0148581
R24745 dvss dvss.n5526 0.0148581
R24746 dvss.n5528 dvss 0.0148581
R24747 dvss.n5527 dvss 0.0148581
R24748 dvss.n1136 dvss 0.0148581
R24749 dvss dvss.n1127 0.0148581
R24750 dvss dvss.n1128 0.0148581
R24751 dvss.n5531 dvss 0.0148581
R24752 dvss.n5530 dvss 0.0148581
R24753 dvss dvss.n1134 0.0148581
R24754 dvss dvss.n1135 0.0148581
R24755 dvss.n5536 dvss 0.0148581
R24756 dvss dvss.n5545 0.0148581
R24757 dvss dvss.n5546 0.0148581
R24758 dvss dvss.n5547 0.0148581
R24759 dvss dvss.n5548 0.0148581
R24760 dvss dvss.n5553 0.0148581
R24761 dvss.n5554 dvss 0.0148581
R24762 dvss dvss.n5559 0.0148581
R24763 dvss dvss.n5560 0.0148581
R24764 dvss dvss.n5566 0.0148581
R24765 dvss dvss.n5567 0.0148581
R24766 dvss dvss.n5568 0.0148581
R24767 dvss.n5570 dvss 0.0148581
R24768 dvss.n5569 dvss 0.0148581
R24769 dvss dvss.n6212 0.0148581
R24770 dvss dvss.n6213 0.0148581
R24771 dvss dvss.n6214 0.0148581
R24772 dvss dvss.n6215 0.0148581
R24773 dvss.n6217 dvss 0.0148581
R24774 dvss.n6216 dvss 0.0148581
R24775 dvss dvss.n512 0.0148581
R24776 dvss.n516 dvss 0.0148581
R24777 dvss.n515 dvss 0.0148581
R24778 dvss.n6235 dvss 0.0148581
R24779 dvss.n6234 dvss 0.0148581
R24780 dvss dvss.n6244 0.0148581
R24781 dvss dvss.n6245 0.0148581
R24782 dvss.n6247 dvss 0.0148581
R24783 dvss.n6246 dvss 0.0148581
R24784 dvss dvss.n6256 0.0148581
R24785 dvss.n6257 dvss 0.0148581
R24786 dvss.n6263 dvss 0.0148581
R24787 dvss.n6262 dvss 0.0148581
R24788 dvss dvss.n6271 0.0148581
R24789 dvss dvss.n6272 0.0148581
R24790 dvss.n6274 dvss 0.0148581
R24791 dvss.n6273 dvss 0.0148581
R24792 dvss dvss.n6283 0.0148581
R24793 dvss dvss.n6284 0.0148581
R24794 dvss dvss.n6285 0.0148581
R24795 dvss.n6288 dvss 0.0148581
R24796 dvss.n6287 dvss 0.0148581
R24797 dvss.n6286 dvss 0.0148581
R24798 dvss dvss.n6296 0.0148581
R24799 dvss.n483 dvss 0.0148581
R24800 dvss.n6305 dvss 0.0148581
R24801 dvss.n6304 dvss 0.0148581
R24802 dvss.n6303 dvss 0.0148581
R24803 dvss.n6302 dvss 0.0148581
R24804 dvss dvss.n6319 0.0148581
R24805 dvss.n6320 dvss 0.0148581
R24806 dvss dvss.n6323 0.0148581
R24807 dvss.n6331 dvss 0.0148581
R24808 dvss.n6330 dvss 0.0148581
R24809 dvss.n6329 dvss 0.0148581
R24810 dvss.n6578 dvss 0.0148581
R24811 dvss.n6575 dvss 0.0148581
R24812 dvss.n6574 dvss 0.0148581
R24813 dvss.n6573 dvss 0.0148581
R24814 dvss dvss.n464 0.0148581
R24815 dvss dvss.n6345 0.0148581
R24816 dvss.n6564 dvss 0.0148581
R24817 dvss.n6563 dvss 0.0148581
R24818 dvss dvss.n6559 0.0148581
R24819 dvss.n6560 dvss 0.0148581
R24820 dvss dvss.n231 0.0148581
R24821 dvss dvss.n232 0.0148581
R24822 dvss dvss.n6352 0.0148581
R24823 dvss dvss.n6353 0.0148581
R24824 dvss.n6355 dvss 0.0148581
R24825 dvss.n6354 dvss 0.0148581
R24826 dvss dvss.n6349 0.0148581
R24827 dvss dvss.n6365 0.0148581
R24828 dvss dvss.n6366 0.0148581
R24829 dvss dvss.n6367 0.0148581
R24830 dvss dvss.n6368 0.0148581
R24831 dvss dvss.n6373 0.0148581
R24832 dvss.n6374 dvss 0.0148581
R24833 dvss dvss.n6379 0.0148581
R24834 dvss dvss.n6380 0.0148581
R24835 dvss dvss.n6386 0.0148581
R24836 dvss dvss.n6387 0.0148581
R24837 dvss dvss.n6388 0.0148581
R24838 dvss dvss.n6389 0.0148581
R24839 dvss dvss.n6394 0.0148581
R24840 dvss dvss.n6395 0.0148581
R24841 dvss.n6413 dvss 0.0148581
R24842 dvss dvss.n6396 0.0148581
R24843 dvss.n6411 dvss 0.0148581
R24844 dvss dvss.n6397 0.0148581
R24845 dvss dvss.n6417 0.0148581
R24846 dvss.n6415 dvss 0.0148581
R24847 dvss dvss.n6403 0.0148581
R24848 dvss dvss.n6404 0.0148581
R24849 dvss dvss.n6405 0.0148581
R24850 dvss.n6422 dvss 0.0148581
R24851 dvss dvss.n6426 0.0148581
R24852 dvss dvss.n6427 0.0148581
R24853 dvss.n6428 dvss 0.0148581
R24854 dvss.n1583 dvss 0.0145449
R24855 dvss.n3233 dvss 0.0140135
R24856 dvss dvss.n5118 0.0140135
R24857 dvss dvss.n7052 0.0134032
R24858 dvss.n1264 dvss 0.0134032
R24859 dvss dvss.n2239 0.0134032
R24860 dvss.n1296 dvss 0.0134032
R24861 dvss dvss.n2189 0.0134032
R24862 dvss.n1327 dvss 0.0134032
R24863 dvss dvss.n2134 0.0134032
R24864 dvss.n5764 dvss 0.0134032
R24865 dvss.n5782 dvss 0.0134032
R24866 dvss.n5850 dvss 0.0134032
R24867 dvss dvss.n5866 0.0134032
R24868 dvss.n5909 dvss 0.0134032
R24869 dvss dvss.n6090 0.0134032
R24870 dvss.n5957 dvss 0.0134032
R24871 dvss dvss.n6040 0.0134032
R24872 dvss.n6744 dvss 0.0134032
R24873 dvss dvss.n6760 0.0134032
R24874 dvss.n6798 dvss 0.0134032
R24875 dvss dvss.n6831 0.0134032
R24876 dvss.n1838 dvss 0.0127893
R24877 dvss.n1978 dvss 0.0127893
R24878 dvss.n1376 dvss 0.0127893
R24879 dvss.n5691 dvss 0.0127893
R24880 dvss dvss.n5640 0.0127893
R24881 dvss.n626 dvss 0.0127893
R24882 dvss.n719 dvss 0.0127893
R24883 dvss.n6675 dvss 0.0127893
R24884 dvss.n6456 dvss 0.0127893
R24885 dvss dvss.n2252 0.0125968
R24886 dvss.n2240 dvss 0.0125968
R24887 dvss dvss.n2202 0.0125968
R24888 dvss.n2190 dvss 0.0125968
R24889 dvss dvss.n2147 0.0125968
R24890 dvss.n2135 dvss 0.0125968
R24891 dvss.n5759 dvss 0.0125968
R24892 dvss.n5780 dvss 0.0125968
R24893 dvss dvss.n5840 0.0125968
R24894 dvss.n5867 dvss 0.0125968
R24895 dvss dvss.n6103 0.0125968
R24896 dvss.n6091 dvss 0.0125968
R24897 dvss dvss.n6053 0.0125968
R24898 dvss.n6041 dvss 0.0125968
R24899 dvss dvss.n6734 0.0125968
R24900 dvss.n6761 dvss 0.0125968
R24901 dvss dvss.n6844 0.0125968
R24902 dvss.n6832 dvss 0.0125968
R24903 dvss dvss.n3332 0.0123243
R24904 dvss.n5133 dvss 0.0123243
R24905 dvss.n5172 dvss 0.0123243
R24906 dvss.n5211 dvss 0.0123243
R24907 dvss.n5250 dvss 0.0123243
R24908 dvss.n5500 dvss 0.0123243
R24909 dvss.n5554 dvss 0.0123243
R24910 dvss.n6257 dvss 0.0123243
R24911 dvss dvss.n6329 0.0123243
R24912 dvss.n6374 dvss 0.0123243
R24913 dvss.n1784 dvss 0.011736
R24914 dvss dvss.n1543 0.011736
R24915 dvss dvss.n1905 0.011736
R24916 dvss dvss.n1477 0.011736
R24917 dvss.n2066 dvss 0.011736
R24918 dvss dvss.n2089 0.011736
R24919 dvss.n5711 dvss 0.011736
R24920 dvss.n5702 dvss 0.011736
R24921 dvss dvss.n1064 0.011736
R24922 dvss dvss.n1074 0.011736
R24923 dvss.n6169 dvss 0.011736
R24924 dvss dvss.n6192 0.011736
R24925 dvss.n739 dvss 0.011736
R24926 dvss.n730 dvss 0.011736
R24927 dvss.n6695 dvss 0.011736
R24928 dvss.n6686 dvss 0.011736
R24929 dvss.n6910 dvss 0.011736
R24930 dvss dvss.n6933 0.011736
R24931 dvss dvss.n3156 0.0114797
R24932 dvss dvss.n3283 0.0114797
R24933 dvss.n3245 dvss 0.0114797
R24934 dvss dvss.n5149 0.0114797
R24935 dvss dvss.n5165 0.0114797
R24936 dvss dvss.n5188 0.0114797
R24937 dvss dvss.n5204 0.0114797
R24938 dvss dvss.n5227 0.0114797
R24939 dvss dvss.n5243 0.0114797
R24940 dvss dvss.n5266 0.0114797
R24941 dvss dvss.n5282 0.0114797
R24942 dvss dvss.n1129 0.0114797
R24943 dvss dvss.n5539 0.0114797
R24944 dvss.n6227 dvss 0.0114797
R24945 dvss.n6231 dvss 0.0114797
R24946 dvss.n6297 dvss 0.0114797
R24947 dvss dvss.n6318 0.0114797
R24948 dvss dvss.n233 0.0114797
R24949 dvss.n6555 dvss 0.0114797
R24950 dvss.n6418 dvss 0.0114797
R24951 dvss dvss.n6425 0.0114797
R24952 dvss dvss.n1788 0.0110337
R24953 dvss dvss.n1810 0.0110337
R24954 dvss.n1906 dvss 0.0110337
R24955 dvss dvss.n1925 0.0110337
R24956 dvss.n2065 dvss 0.0110337
R24957 dvss.n2090 dvss 0.0110337
R24958 dvss.n915 dvss 0.0110337
R24959 dvss.n5696 dvss 0.0110337
R24960 dvss.n1082 dvss 0.0110337
R24961 dvss.n1096 dvss 0.0110337
R24962 dvss.n6168 dvss 0.0110337
R24963 dvss.n6193 dvss 0.0110337
R24964 dvss.n561 dvss 0.0110337
R24965 dvss.n724 dvss 0.0110337
R24966 dvss.n149 dvss 0.0110337
R24967 dvss.n6680 dvss 0.0110337
R24968 dvss.n6909 dvss 0.0110337
R24969 dvss.n6934 dvss 0.0110337
R24970 dvss dvss.n1830 0.00998034
R24971 dvss.n1944 dvss 0.00998034
R24972 dvss dvss.n2097 0.00998034
R24973 dvss.n940 dvss 0.00998034
R24974 dvss.n5641 dvss 0.00998034
R24975 dvss dvss.n6200 0.00998034
R24976 dvss.n586 dvss 0.00998034
R24977 dvss.n170 dvss 0.00998034
R24978 dvss dvss.n6941 0.00998034
R24979 dvss dvss.n3150 0.00979054
R24980 dvss dvss.n3157 0.00979054
R24981 dvss.n3248 dvss 0.00979054
R24982 dvss dvss.n5102 0.00979054
R24983 dvss dvss.n5146 0.00979054
R24984 dvss dvss.n5150 0.00979054
R24985 dvss dvss.n5185 0.00979054
R24986 dvss dvss.n5189 0.00979054
R24987 dvss dvss.n5224 0.00979054
R24988 dvss dvss.n5228 0.00979054
R24989 dvss dvss.n5263 0.00979054
R24990 dvss dvss.n5267 0.00979054
R24991 dvss dvss.n5527 0.00979054
R24992 dvss dvss.n5530 0.00979054
R24993 dvss.n6214 dvss 0.00979054
R24994 dvss.n516 dvss 0.00979054
R24995 dvss.n6288 dvss 0.00979054
R24996 dvss.n6305 dvss 0.00979054
R24997 dvss.n6559 dvss 0.00979054
R24998 dvss.n6353 dvss 0.00979054
R24999 dvss dvss.n6396 0.00979054
R25000 dvss dvss.n6403 0.00979054
R25001 dvss.n2263 dvss 0.00896774
R25002 dvss.n3330 dvss 0.00894595
R25003 dvss dvss.n5137 0.00894595
R25004 dvss dvss.n5176 0.00894595
R25005 dvss dvss.n5215 0.00894595
R25006 dvss dvss.n5254 0.00894595
R25007 dvss dvss.n5504 0.00894595
R25008 dvss dvss.n5558 0.00894595
R25009 dvss dvss.n6261 0.00894595
R25010 dvss.n6327 dvss 0.00894595
R25011 dvss dvss.n6378 0.00894595
R25012 dvss.n6579 dvss 0.00810135
R25013 dvss dvss.n5099 0.00755
R25014 dvss dvss.n1767 0.00752247
R25015 dvss.n7056 dvss 0.00735484
R25016 dvss.n7053 dvss 0.00735484
R25017 dvss dvss.n4 0.00735484
R25018 dvss.n2286 dvss 0.00735484
R25019 dvss.n2285 dvss 0.00735484
R25020 dvss.n2284 dvss 0.00735484
R25021 dvss.n2280 dvss 0.00735484
R25022 dvss.n2278 dvss 0.00735484
R25023 dvss.n2277 dvss 0.00735484
R25024 dvss.n2269 dvss 0.00735484
R25025 dvss.n2266 dvss 0.00735484
R25026 dvss.n2265 dvss 0.00735484
R25027 dvss.n1256 dvss 0.00735484
R25028 dvss dvss.n1256 0.00735484
R25029 dvss.n2263 dvss 0.00735484
R25030 dvss.n2262 dvss 0.00735484
R25031 dvss.n2259 dvss 0.00735484
R25032 dvss.n2258 dvss 0.00735484
R25033 dvss.n2257 dvss 0.00735484
R25034 dvss.n2254 dvss 0.00735484
R25035 dvss.n2253 dvss 0.00735484
R25036 dvss.n2252 dvss 0.00735484
R25037 dvss.n1264 dvss 0.00735484
R25038 dvss.n2249 dvss 0.00735484
R25039 dvss.n2248 dvss 0.00735484
R25040 dvss.n2245 dvss 0.00735484
R25041 dvss.n2244 dvss 0.00735484
R25042 dvss dvss.n1271 0.00735484
R25043 dvss.n2240 dvss 0.00735484
R25044 dvss.n2239 dvss 0.00735484
R25045 dvss.n2236 dvss 0.00735484
R25046 dvss.n2232 dvss 0.00735484
R25047 dvss.n2231 dvss 0.00735484
R25048 dvss.n2228 dvss 0.00735484
R25049 dvss.n2227 dvss 0.00735484
R25050 dvss.n2226 dvss 0.00735484
R25051 dvss.n2222 dvss 0.00735484
R25052 dvss.n2221 dvss 0.00735484
R25053 dvss.n2218 dvss 0.00735484
R25054 dvss.n2217 dvss 0.00735484
R25055 dvss.n2216 dvss 0.00735484
R25056 dvss.n2213 dvss 0.00735484
R25057 dvss.n2212 dvss 0.00735484
R25058 dvss.n2211 dvss 0.00735484
R25059 dvss.n2208 dvss 0.00735484
R25060 dvss.n2207 dvss 0.00735484
R25061 dvss.n2206 dvss 0.00735484
R25062 dvss.n2203 dvss 0.00735484
R25063 dvss.n2202 dvss 0.00735484
R25064 dvss dvss.n1296 0.00735484
R25065 dvss.n2199 dvss 0.00735484
R25066 dvss.n2198 dvss 0.00735484
R25067 dvss.n2195 dvss 0.00735484
R25068 dvss.n2194 dvss 0.00735484
R25069 dvss dvss.n1302 0.00735484
R25070 dvss.n2190 dvss 0.00735484
R25071 dvss.n2189 dvss 0.00735484
R25072 dvss.n2186 dvss 0.00735484
R25073 dvss.n2182 dvss 0.00735484
R25074 dvss.n2181 dvss 0.00735484
R25075 dvss.n2178 dvss 0.00735484
R25076 dvss.n2177 dvss 0.00735484
R25077 dvss.n2176 dvss 0.00735484
R25078 dvss.n2172 dvss 0.00735484
R25079 dvss.n2171 dvss 0.00735484
R25080 dvss.n2168 dvss 0.00735484
R25081 dvss.n2162 dvss 0.00735484
R25082 dvss.n2161 dvss 0.00735484
R25083 dvss.n2158 dvss 0.00735484
R25084 dvss.n2157 dvss 0.00735484
R25085 dvss.n2156 dvss 0.00735484
R25086 dvss.n2153 dvss 0.00735484
R25087 dvss.n2152 dvss 0.00735484
R25088 dvss.n2151 dvss 0.00735484
R25089 dvss.n2148 dvss 0.00735484
R25090 dvss.n2147 dvss 0.00735484
R25091 dvss dvss.n1327 0.00735484
R25092 dvss.n2144 dvss 0.00735484
R25093 dvss.n2143 dvss 0.00735484
R25094 dvss.n2140 dvss 0.00735484
R25095 dvss.n2139 dvss 0.00735484
R25096 dvss dvss.n1333 0.00735484
R25097 dvss.n2135 dvss 0.00735484
R25098 dvss.n2134 dvss 0.00735484
R25099 dvss.n2131 dvss 0.00735484
R25100 dvss.n2127 dvss 0.00735484
R25101 dvss.n2126 dvss 0.00735484
R25102 dvss.n2123 dvss 0.00735484
R25103 dvss.n2122 dvss 0.00735484
R25104 dvss.n2121 dvss 0.00735484
R25105 dvss.n2117 dvss 0.00735484
R25106 dvss.n2116 dvss 0.00735484
R25107 dvss.n1344 dvss 0.00735484
R25108 dvss dvss.n5736 0.00735484
R25109 dvss dvss.n5737 0.00735484
R25110 dvss.n5748 dvss 0.00735484
R25111 dvss.n5747 dvss 0.00735484
R25112 dvss.n5746 dvss 0.00735484
R25113 dvss.n5743 dvss 0.00735484
R25114 dvss.n5742 dvss 0.00735484
R25115 dvss dvss.n5757 0.00735484
R25116 dvss dvss.n5758 0.00735484
R25117 dvss.n5759 dvss 0.00735484
R25118 dvss.n5764 dvss 0.00735484
R25119 dvss.n5763 dvss 0.00735484
R25120 dvss.n871 dvss 0.00735484
R25121 dvss dvss.n5772 0.00735484
R25122 dvss.n5774 dvss 0.00735484
R25123 dvss.n5773 dvss 0.00735484
R25124 dvss dvss.n5780 0.00735484
R25125 dvss.n5782 dvss 0.00735484
R25126 dvss.n5781 dvss 0.00735484
R25127 dvss dvss.n5793 0.00735484
R25128 dvss dvss.n5794 0.00735484
R25129 dvss.n5796 dvss 0.00735484
R25130 dvss.n5795 dvss 0.00735484
R25131 dvss dvss.n853 0.00735484
R25132 dvss dvss.n5809 0.00735484
R25133 dvss dvss.n5810 0.00735484
R25134 dvss.n5817 dvss 0.00735484
R25135 dvss.n5811 dvss 0.00735484
R25136 dvss dvss.n5827 0.00735484
R25137 dvss dvss.n5828 0.00735484
R25138 dvss.n5830 dvss 0.00735484
R25139 dvss.n5829 dvss 0.00735484
R25140 dvss dvss.n5838 0.00735484
R25141 dvss dvss.n5839 0.00735484
R25142 dvss.n5842 dvss 0.00735484
R25143 dvss.n5841 dvss 0.00735484
R25144 dvss.n5840 dvss 0.00735484
R25145 dvss dvss.n5850 0.00735484
R25146 dvss.n5852 dvss 0.00735484
R25147 dvss.n5851 dvss 0.00735484
R25148 dvss.n5857 dvss 0.00735484
R25149 dvss.n5856 dvss 0.00735484
R25150 dvss.n835 dvss 0.00735484
R25151 dvss.n5867 dvss 0.00735484
R25152 dvss.n5866 dvss 0.00735484
R25153 dvss.n829 dvss 0.00735484
R25154 dvss.n5871 dvss 0.00735484
R25155 dvss.n826 dvss 0.00735484
R25156 dvss dvss.n5881 0.00735484
R25157 dvss dvss.n5882 0.00735484
R25158 dvss.n5883 dvss 0.00735484
R25159 dvss.n819 dvss 0.00735484
R25160 dvss.n818 dvss 0.00735484
R25161 dvss dvss.n5895 0.00735484
R25162 dvss dvss.n5901 0.00735484
R25163 dvss.n6115 dvss 0.00735484
R25164 dvss.n6114 dvss 0.00735484
R25165 dvss.n6113 dvss 0.00735484
R25166 dvss.n6110 dvss 0.00735484
R25167 dvss.n6109 dvss 0.00735484
R25168 dvss.n6108 dvss 0.00735484
R25169 dvss.n6105 dvss 0.00735484
R25170 dvss.n6104 dvss 0.00735484
R25171 dvss.n6103 dvss 0.00735484
R25172 dvss.n5909 dvss 0.00735484
R25173 dvss.n6100 dvss 0.00735484
R25174 dvss.n6099 dvss 0.00735484
R25175 dvss.n6096 dvss 0.00735484
R25176 dvss.n6095 dvss 0.00735484
R25177 dvss dvss.n5916 0.00735484
R25178 dvss.n6091 dvss 0.00735484
R25179 dvss.n6090 dvss 0.00735484
R25180 dvss.n6087 dvss 0.00735484
R25181 dvss.n6083 dvss 0.00735484
R25182 dvss.n6082 dvss 0.00735484
R25183 dvss.n6079 dvss 0.00735484
R25184 dvss.n6078 dvss 0.00735484
R25185 dvss.n6077 dvss 0.00735484
R25186 dvss.n6073 dvss 0.00735484
R25187 dvss.n6072 dvss 0.00735484
R25188 dvss.n6069 dvss 0.00735484
R25189 dvss.n6068 dvss 0.00735484
R25190 dvss.n6067 dvss 0.00735484
R25191 dvss.n6064 dvss 0.00735484
R25192 dvss.n6063 dvss 0.00735484
R25193 dvss.n6062 dvss 0.00735484
R25194 dvss.n6059 dvss 0.00735484
R25195 dvss.n6058 dvss 0.00735484
R25196 dvss.n6057 dvss 0.00735484
R25197 dvss.n6054 dvss 0.00735484
R25198 dvss.n6053 dvss 0.00735484
R25199 dvss dvss.n5957 0.00735484
R25200 dvss.n6050 dvss 0.00735484
R25201 dvss.n6049 dvss 0.00735484
R25202 dvss.n6046 dvss 0.00735484
R25203 dvss.n6045 dvss 0.00735484
R25204 dvss dvss.n5963 0.00735484
R25205 dvss.n6041 dvss 0.00735484
R25206 dvss.n6040 dvss 0.00735484
R25207 dvss.n6037 dvss 0.00735484
R25208 dvss.n6033 dvss 0.00735484
R25209 dvss.n6032 dvss 0.00735484
R25210 dvss.n6029 dvss 0.00735484
R25211 dvss.n6028 dvss 0.00735484
R25212 dvss.n6027 dvss 0.00735484
R25213 dvss.n6023 dvss 0.00735484
R25214 dvss.n6022 dvss 0.00735484
R25215 dvss.n6019 dvss 0.00735484
R25216 dvss.n6018 dvss 0.00735484
R25217 dvss dvss.n6721 0.00735484
R25218 dvss dvss.n6722 0.00735484
R25219 dvss.n6724 dvss 0.00735484
R25220 dvss.n6723 dvss 0.00735484
R25221 dvss dvss.n6732 0.00735484
R25222 dvss dvss.n6733 0.00735484
R25223 dvss.n6736 dvss 0.00735484
R25224 dvss.n6735 dvss 0.00735484
R25225 dvss.n6734 dvss 0.00735484
R25226 dvss dvss.n6744 0.00735484
R25227 dvss.n6746 dvss 0.00735484
R25228 dvss.n6745 dvss 0.00735484
R25229 dvss.n6751 dvss 0.00735484
R25230 dvss.n6750 dvss 0.00735484
R25231 dvss.n106 dvss 0.00735484
R25232 dvss.n6761 dvss 0.00735484
R25233 dvss.n6760 dvss 0.00735484
R25234 dvss.n100 dvss 0.00735484
R25235 dvss.n6765 dvss 0.00735484
R25236 dvss.n97 dvss 0.00735484
R25237 dvss dvss.n6775 0.00735484
R25238 dvss dvss.n6776 0.00735484
R25239 dvss.n6777 dvss 0.00735484
R25240 dvss.n90 dvss 0.00735484
R25241 dvss.n89 dvss 0.00735484
R25242 dvss dvss.n6789 0.00735484
R25243 dvss dvss.n6790 0.00735484
R25244 dvss.n6856 dvss 0.00735484
R25245 dvss.n6855 dvss 0.00735484
R25246 dvss.n6854 dvss 0.00735484
R25247 dvss.n6851 dvss 0.00735484
R25248 dvss.n6850 dvss 0.00735484
R25249 dvss.n6849 dvss 0.00735484
R25250 dvss.n6846 dvss 0.00735484
R25251 dvss.n6845 dvss 0.00735484
R25252 dvss.n6844 dvss 0.00735484
R25253 dvss.n6798 dvss 0.00735484
R25254 dvss.n6841 dvss 0.00735484
R25255 dvss.n6840 dvss 0.00735484
R25256 dvss.n6837 dvss 0.00735484
R25257 dvss.n6836 dvss 0.00735484
R25258 dvss dvss.n6805 0.00735484
R25259 dvss.n6832 dvss 0.00735484
R25260 dvss.n6831 dvss 0.00735484
R25261 dvss.n6828 dvss 0.00735484
R25262 dvss.n6824 dvss 0.00735484
R25263 dvss dvss.n6954 0.00735484
R25264 dvss dvss.n6955 0.00735484
R25265 dvss.n6964 dvss 0.00735484
R25266 dvss.n6963 dvss 0.00735484
R25267 dvss.n6959 dvss 0.00735484
R25268 dvss dvss.n6972 0.00735484
R25269 dvss dvss.n6973 0.00735484
R25270 dvss.n6977 dvss 0.00735484
R25271 dvss.n6976 dvss 0.00735484
R25272 dvss.n6975 dvss 0.00735484
R25273 dvss.n6974 dvss 0.00735484
R25274 dvss dvss.n6988 0.00735484
R25275 dvss dvss.n3188 0.00725676
R25276 dvss dvss.n3179 0.00725676
R25277 dvss.n6579 dvss.n458 0.00725676
R25278 dvss dvss.n2278 0.00695161
R25279 dvss dvss.n1275 0.00695161
R25280 dvss dvss.n1306 0.00695161
R25281 dvss dvss.n1337 0.00695161
R25282 dvss.n5790 dvss 0.00695161
R25283 dvss.n5872 dvss 0.00695161
R25284 dvss dvss.n5936 0.00695161
R25285 dvss dvss.n5967 0.00695161
R25286 dvss.n6766 dvss 0.00695161
R25287 dvss dvss.n6823 0.00695161
R25288 dvss.n2274 dvss.n2273 0.00654839
R25289 dvss.n1711 dvss 0.0064691
R25290 dvss.n1588 dvss 0.0064691
R25291 dvss dvss.n1777 0.0064691
R25292 dvss.n1778 dvss 0.0064691
R25293 dvss.n1789 dvss 0.0064691
R25294 dvss.n1788 dvss 0.0064691
R25295 dvss dvss.n1784 0.0064691
R25296 dvss.n1785 dvss 0.0064691
R25297 dvss.n1800 dvss 0.0064691
R25298 dvss dvss.n1803 0.0064691
R25299 dvss.n1804 dvss 0.0064691
R25300 dvss.n1811 dvss 0.0064691
R25301 dvss.n1810 dvss 0.0064691
R25302 dvss.n1543 dvss 0.0064691
R25303 dvss.n1823 dvss 0.0064691
R25304 dvss.n1831 dvss 0.0064691
R25305 dvss.n1830 dvss 0.0064691
R25306 dvss dvss.n1838 0.0064691
R25307 dvss.n1845 dvss 0.0064691
R25308 dvss.n1844 dvss 0.0064691
R25309 dvss.n1857 dvss 0.0064691
R25310 dvss.n1856 dvss 0.0064691
R25311 dvss.n1866 dvss 0.0064691
R25312 dvss.n1865 dvss 0.0064691
R25313 dvss.n1869 dvss 0.0064691
R25314 dvss.n1884 dvss 0.0064691
R25315 dvss.n1883 dvss 0.0064691
R25316 dvss.n1882 dvss 0.0064691
R25317 dvss dvss.n1892 0.0064691
R25318 dvss.n1893 dvss 0.0064691
R25319 dvss.n1898 dvss 0.0064691
R25320 dvss.n1906 dvss 0.0064691
R25321 dvss.n1905 dvss 0.0064691
R25322 dvss dvss.n1910 0.0064691
R25323 dvss.n1911 dvss 0.0064691
R25324 dvss dvss.n1918 0.0064691
R25325 dvss.n1919 dvss 0.0064691
R25326 dvss.n1926 dvss 0.0064691
R25327 dvss.n1925 dvss 0.0064691
R25328 dvss.n1477 dvss 0.0064691
R25329 dvss dvss.n1937 0.0064691
R25330 dvss.n1981 dvss 0.0064691
R25331 dvss dvss.n1944 0.0064691
R25332 dvss.n1978 dvss 0.0064691
R25333 dvss.n1977 dvss 0.0064691
R25334 dvss.n1976 dvss 0.0064691
R25335 dvss.n1967 dvss 0.0064691
R25336 dvss.n1964 dvss 0.0064691
R25337 dvss dvss.n2021 0.0064691
R25338 dvss.n2022 dvss 0.0064691
R25339 dvss.n2052 dvss 0.0064691
R25340 dvss.n2049 dvss 0.0064691
R25341 dvss.n2048 dvss 0.0064691
R25342 dvss.n2047 dvss 0.0064691
R25343 dvss.n2040 dvss 0.0064691
R25344 dvss.n2039 dvss 0.0064691
R25345 dvss dvss.n2064 0.0064691
R25346 dvss dvss.n2065 0.0064691
R25347 dvss.n2066 dvss 0.0064691
R25348 dvss.n2074 dvss 0.0064691
R25349 dvss.n2073 dvss 0.0064691
R25350 dvss.n2079 dvss 0.0064691
R25351 dvss.n2078 dvss 0.0064691
R25352 dvss.n1426 dvss 0.0064691
R25353 dvss.n2090 dvss 0.0064691
R25354 dvss.n2089 dvss 0.0064691
R25355 dvss.n1413 dvss 0.0064691
R25356 dvss.n2098 dvss 0.0064691
R25357 dvss.n2097 dvss 0.0064691
R25358 dvss.n1376 dvss 0.0064691
R25359 dvss dvss.n1384 0.0064691
R25360 dvss.n1385 dvss 0.0064691
R25361 dvss.n1373 dvss 0.0064691
R25362 dvss dvss.n1399 0.0064691
R25363 dvss dvss.n1405 0.0064691
R25364 dvss.n1406 dvss 0.0064691
R25365 dvss.n5724 dvss 0.0064691
R25366 dvss.n5723 dvss 0.0064691
R25367 dvss.n5722 dvss 0.0064691
R25368 dvss.n5719 dvss 0.0064691
R25369 dvss.n5718 dvss 0.0064691
R25370 dvss.n5717 dvss 0.0064691
R25371 dvss.n5714 dvss 0.0064691
R25372 dvss.n915 dvss 0.0064691
R25373 dvss.n5711 dvss 0.0064691
R25374 dvss.n5710 dvss 0.0064691
R25375 dvss dvss.n995 0.0064691
R25376 dvss.n996 dvss 0.0064691
R25377 dvss.n5706 dvss 0.0064691
R25378 dvss.n5705 dvss 0.0064691
R25379 dvss.n5696 dvss 0.0064691
R25380 dvss.n5702 dvss 0.0064691
R25381 dvss.n5701 dvss 0.0064691
R25382 dvss.n5694 dvss 0.0064691
R25383 dvss.n940 dvss 0.0064691
R25384 dvss.n5691 dvss 0.0064691
R25385 dvss.n5690 dvss 0.0064691
R25386 dvss.n5689 dvss 0.0064691
R25387 dvss.n1044 dvss 0.0064691
R25388 dvss.n987 dvss 0.0064691
R25389 dvss.n981 dvss 0.0064691
R25390 dvss dvss.n943 0.0064691
R25391 dvss.n5675 dvss 0.0064691
R25392 dvss.n5674 dvss 0.0064691
R25393 dvss.n5673 dvss 0.0064691
R25394 dvss.n968 dvss 0.0064691
R25395 dvss dvss.n956 0.0064691
R25396 dvss.n958 dvss 0.0064691
R25397 dvss dvss.n963 0.0064691
R25398 dvss.n1082 dvss 0.0064691
R25399 dvss dvss.n1064 0.0064691
R25400 dvss.n1085 dvss 0.0064691
R25401 dvss dvss.n1065 0.0064691
R25402 dvss dvss.n1091 0.0064691
R25403 dvss.n1092 dvss 0.0064691
R25404 dvss dvss.n1073 0.0064691
R25405 dvss.n1096 dvss 0.0064691
R25406 dvss dvss.n1074 0.0064691
R25407 dvss.n5648 dvss 0.0064691
R25408 dvss.n1114 dvss 0.0064691
R25409 dvss.n5641 dvss 0.0064691
R25410 dvss.n5640 dvss 0.0064691
R25411 dvss.n5637 dvss 0.0064691
R25412 dvss.n5636 dvss 0.0064691
R25413 dvss.n5627 dvss 0.0064691
R25414 dvss.n5624 dvss 0.0064691
R25415 dvss dvss.n6124 0.0064691
R25416 dvss.n6125 dvss 0.0064691
R25417 dvss.n6155 dvss 0.0064691
R25418 dvss.n6152 dvss 0.0064691
R25419 dvss.n6151 dvss 0.0064691
R25420 dvss.n6150 dvss 0.0064691
R25421 dvss.n6143 dvss 0.0064691
R25422 dvss.n6142 dvss 0.0064691
R25423 dvss dvss.n6167 0.0064691
R25424 dvss dvss.n6168 0.0064691
R25425 dvss.n6169 dvss 0.0064691
R25426 dvss.n6177 dvss 0.0064691
R25427 dvss.n6176 dvss 0.0064691
R25428 dvss.n6182 dvss 0.0064691
R25429 dvss.n6181 dvss 0.0064691
R25430 dvss.n776 dvss 0.0064691
R25431 dvss.n6193 dvss 0.0064691
R25432 dvss.n6192 dvss 0.0064691
R25433 dvss.n763 dvss 0.0064691
R25434 dvss.n6201 dvss 0.0064691
R25435 dvss.n6200 dvss 0.0064691
R25436 dvss.n626 dvss 0.0064691
R25437 dvss dvss.n636 0.0064691
R25438 dvss.n637 dvss 0.0064691
R25439 dvss.n644 dvss 0.0064691
R25440 dvss.n618 dvss 0.0064691
R25441 dvss.n617 dvss 0.0064691
R25442 dvss dvss.n538 0.0064691
R25443 dvss.n752 dvss 0.0064691
R25444 dvss.n751 dvss 0.0064691
R25445 dvss.n750 dvss 0.0064691
R25446 dvss.n747 dvss 0.0064691
R25447 dvss.n746 dvss 0.0064691
R25448 dvss.n745 dvss 0.0064691
R25449 dvss.n742 dvss 0.0064691
R25450 dvss.n561 dvss 0.0064691
R25451 dvss.n739 dvss 0.0064691
R25452 dvss.n738 dvss 0.0064691
R25453 dvss dvss.n603 0.0064691
R25454 dvss.n604 dvss 0.0064691
R25455 dvss.n734 dvss 0.0064691
R25456 dvss.n733 dvss 0.0064691
R25457 dvss.n724 dvss 0.0064691
R25458 dvss.n730 dvss 0.0064691
R25459 dvss.n729 dvss 0.0064691
R25460 dvss.n722 dvss 0.0064691
R25461 dvss.n586 dvss 0.0064691
R25462 dvss.n719 dvss 0.0064691
R25463 dvss.n718 dvss 0.0064691
R25464 dvss.n717 dvss 0.0064691
R25465 dvss.n595 dvss 0.0064691
R25466 dvss dvss.n705 0.0064691
R25467 dvss dvss.n706 0.0064691
R25468 dvss.n707 dvss 0.0064691
R25469 dvss.n6708 dvss 0.0064691
R25470 dvss.n6707 dvss 0.0064691
R25471 dvss.n6706 dvss 0.0064691
R25472 dvss.n6703 dvss 0.0064691
R25473 dvss.n6702 dvss 0.0064691
R25474 dvss.n6701 dvss 0.0064691
R25475 dvss.n6698 dvss 0.0064691
R25476 dvss.n149 dvss 0.0064691
R25477 dvss.n6695 dvss 0.0064691
R25478 dvss.n6694 dvss 0.0064691
R25479 dvss dvss.n212 0.0064691
R25480 dvss.n213 dvss 0.0064691
R25481 dvss.n6690 dvss 0.0064691
R25482 dvss.n6689 dvss 0.0064691
R25483 dvss.n6680 dvss 0.0064691
R25484 dvss.n6686 dvss 0.0064691
R25485 dvss.n6685 dvss 0.0064691
R25486 dvss.n6678 dvss 0.0064691
R25487 dvss dvss.n170 0.0064691
R25488 dvss.n6675 dvss 0.0064691
R25489 dvss.n6674 dvss 0.0064691
R25490 dvss.n6673 dvss 0.0064691
R25491 dvss.n6664 dvss 0.0064691
R25492 dvss.n6661 dvss 0.0064691
R25493 dvss dvss.n6865 0.0064691
R25494 dvss.n6866 dvss 0.0064691
R25495 dvss.n6896 dvss 0.0064691
R25496 dvss.n6893 dvss 0.0064691
R25497 dvss.n6892 dvss 0.0064691
R25498 dvss.n6891 dvss 0.0064691
R25499 dvss.n6884 dvss 0.0064691
R25500 dvss.n6883 dvss 0.0064691
R25501 dvss dvss.n6908 0.0064691
R25502 dvss dvss.n6909 0.0064691
R25503 dvss.n6910 dvss 0.0064691
R25504 dvss.n6918 dvss 0.0064691
R25505 dvss.n6917 dvss 0.0064691
R25506 dvss.n6923 dvss 0.0064691
R25507 dvss.n6922 dvss 0.0064691
R25508 dvss.n52 dvss 0.0064691
R25509 dvss.n6934 dvss 0.0064691
R25510 dvss.n6933 dvss 0.0064691
R25511 dvss.n39 dvss 0.0064691
R25512 dvss.n6942 dvss 0.0064691
R25513 dvss.n6941 dvss 0.0064691
R25514 dvss.n6456 dvss 0.0064691
R25515 dvss dvss.n6463 0.0064691
R25516 dvss.n6464 dvss 0.0064691
R25517 dvss dvss.n6475 0.0064691
R25518 dvss.n6476 dvss 0.0064691
R25519 dvss dvss.n6483 0.0064691
R25520 dvss.n6484 dvss 0.0064691
R25521 dvss dvss.n6494 0.0064691
R25522 dvss.n6495 dvss 0.0064691
R25523 dvss.n6498 dvss 0.0064691
R25524 dvss.n3330 dvss.n3131 0.00641216
R25525 dvss.n5137 dvss.n5132 0.00641216
R25526 dvss.n5176 dvss.n5171 0.00641216
R25527 dvss.n5215 dvss.n5210 0.00641216
R25528 dvss.n5254 dvss.n5249 0.00641216
R25529 dvss.n5504 dvss.n1148 0.00641216
R25530 dvss.n5558 dvss.n5552 0.00641216
R25531 dvss.n6261 dvss.n499 0.00641216
R25532 dvss.n6327 dvss.n6326 0.00641216
R25533 dvss.n6378 dvss.n6372 0.00641216
R25534 dvss dvss.n1699 0.00611798
R25535 dvss.n1702 dvss 0.00611798
R25536 dvss.n1704 dvss 0.00611798
R25537 dvss.n1705 dvss 0.00611798
R25538 dvss.n1706 dvss 0.00611798
R25539 dvss.n1707 dvss 0.00611798
R25540 dvss dvss.n1708 0.00611798
R25541 dvss dvss.n1605 0.00611798
R25542 dvss.n1713 dvss 0.00611798
R25543 dvss.n1714 dvss 0.00611798
R25544 dvss.n1621 dvss 0.00611798
R25545 dvss dvss.n1759 0.00611798
R25546 dvss.n1764 dvss 0.00611798
R25547 dvss dvss.n1563 0.00611798
R25548 dvss.n1768 dvss 0.00611798
R25549 dvss dvss.n1564 0.00611798
R25550 dvss dvss.n1584 0.00611798
R25551 dvss dvss.n1587 0.00611798
R25552 dvss.n1826 dvss 0.00611798
R25553 dvss.n1938 dvss 0.00611798
R25554 dvss.n2101 dvss 0.00611798
R25555 dvss dvss.n927 0.00611798
R25556 dvss.n5645 dvss 0.00611798
R25557 dvss.n6204 dvss 0.00611798
R25558 dvss dvss.n573 0.00611798
R25559 dvss dvss.n161 0.00611798
R25560 dvss.n6945 dvss 0.00611798
R25561 dvss dvss.n2226 0.00574194
R25562 dvss dvss.n2176 0.00574194
R25563 dvss dvss.n2121 0.00574194
R25564 dvss dvss.n853 0.00574194
R25565 dvss.n5883 dvss 0.00574194
R25566 dvss dvss.n6077 0.00574194
R25567 dvss dvss.n6027 0.00574194
R25568 dvss.n6777 dvss 0.00574194
R25569 dvss dvss.n6963 0.00574194
R25570 dvss dvss.n3641 0.00570833
R25571 dvss.n4001 dvss 0.00570833
R25572 dvss.n2403 dvss 0.00570833
R25573 dvss dvss.n4572 0.00570833
R25574 dvss.n3213 dvss 0.00556757
R25575 dvss.n3249 dvss.n3248 0.00556757
R25576 dvss.n5102 dvss.n1208 0.00556757
R25577 dvss.n5112 dvss 0.00556757
R25578 dvss.n1618 dvss.n1617 0.00541573
R25579 dvss.n1778 dvss 0.00541573
R25580 dvss dvss.n1829 0.00541573
R25581 dvss.n1893 dvss 0.00541573
R25582 dvss.n1941 dvss 0.00541573
R25583 dvss dvss.n2039 0.00541573
R25584 dvss.n2094 dvss 0.00541573
R25585 dvss dvss.n5717 0.00541573
R25586 dvss.n5695 dvss 0.00541573
R25587 dvss.n958 dvss 0.00541573
R25588 dvss dvss.n1100 0.00541573
R25589 dvss dvss.n6142 0.00541573
R25590 dvss.n6197 dvss 0.00541573
R25591 dvss dvss.n745 0.00541573
R25592 dvss.n723 dvss 0.00541573
R25593 dvss dvss.n6701 0.00541573
R25594 dvss.n6679 dvss 0.00541573
R25595 dvss dvss.n6883 0.00541573
R25596 dvss.n6938 dvss 0.00541573
R25597 dvss dvss.n1844 0.00506461
R25598 dvss.n1870 dvss 0.00506461
R25599 dvss dvss.n1976 0.00506461
R25600 dvss.n2025 dvss 0.00506461
R25601 dvss.n1385 dvss 0.00506461
R25602 dvss.n5727 dvss 0.00506461
R25603 dvss dvss.n5689 0.00506461
R25604 dvss.n5678 dvss 0.00506461
R25605 dvss dvss.n5636 0.00506461
R25606 dvss.n6128 dvss 0.00506461
R25607 dvss.n637 dvss 0.00506461
R25608 dvss.n755 dvss 0.00506461
R25609 dvss dvss.n717 0.00506461
R25610 dvss.n6711 dvss 0.00506461
R25611 dvss dvss.n6673 0.00506461
R25612 dvss.n6869 dvss 0.00506461
R25613 dvss.n6464 dvss 0.00506461
R25614 dvss.n6487 dvss 0.00506461
R25615 dvss.n2223 dvss 0.00493548
R25616 dvss.n2173 dvss 0.00493548
R25617 dvss.n2118 dvss 0.00493548
R25618 dvss.n5805 dvss 0.00493548
R25619 dvss.n5886 dvss 0.00493548
R25620 dvss.n6074 dvss 0.00493548
R25621 dvss.n6024 dvss 0.00493548
R25622 dvss.n6780 dvss 0.00493548
R25623 dvss.n6960 dvss 0.00493548
R25624 dvss.n1701 dvss.n1599 0.00471348
R25625 dvss.n2281 dvss.n1246 0.00412903
R25626 dvss.n2271 dvss.n2270 0.00412903
R25627 dvss dvss.n1782 0.00401124
R25628 dvss.n1839 dvss.n1514 0.00401124
R25629 dvss dvss.n1897 0.00401124
R25630 dvss.n1972 dvss.n1968 0.00401124
R25631 dvss.n1435 dvss 0.00401124
R25632 dvss.n1374 dvss.n1372 0.00401124
R25633 dvss.n5715 dvss 0.00401124
R25634 dvss.n5685 dvss.n939 0.00401124
R25635 dvss dvss.n962 0.00401124
R25636 dvss.n5632 dvss.n5628 0.00401124
R25637 dvss.n785 dvss 0.00401124
R25638 dvss.n624 dvss.n623 0.00401124
R25639 dvss.n743 dvss 0.00401124
R25640 dvss.n713 dvss.n585 0.00401124
R25641 dvss.n6699 dvss 0.00401124
R25642 dvss.n6669 dvss.n6665 0.00401124
R25643 dvss.n61 dvss 0.00401124
R25644 dvss.n6453 dvss.n6452 0.00401124
R25645 dvss.n3277 dvss.n3156 0.00387838
R25646 dvss.n3283 dvss.n3282 0.00387838
R25647 dvss.n5159 dvss.n5149 0.00387838
R25648 dvss.n5165 dvss.n5164 0.00387838
R25649 dvss.n5198 dvss.n5188 0.00387838
R25650 dvss.n5204 dvss.n5203 0.00387838
R25651 dvss.n5237 dvss.n5227 0.00387838
R25652 dvss.n5243 dvss.n5242 0.00387838
R25653 dvss.n5276 dvss.n5266 0.00387838
R25654 dvss.n5282 dvss.n5281 0.00387838
R25655 dvss.n5533 dvss.n1129 0.00387838
R25656 dvss.n5539 dvss.n5538 0.00387838
R25657 dvss.n6228 dvss.n6227 0.00387838
R25658 dvss.n6232 dvss.n6231 0.00387838
R25659 dvss.n6298 dvss.n6297 0.00387838
R25660 dvss.n6318 dvss.n474 0.00387838
R25661 dvss.n6347 dvss.n233 0.00387838
R25662 dvss.n6556 dvss.n6555 0.00387838
R25663 dvss.n6419 dvss.n6418 0.00387838
R25664 dvss.n6425 dvss.n6424 0.00387838
R25665 dvss.n2281 dvss 0.00372581
R25666 dvss.n2270 dvss 0.00372581
R25667 dvss.n1271 dvss 0.00372581
R25668 dvss dvss.n2231 0.00372581
R25669 dvss.n1302 dvss 0.00372581
R25670 dvss dvss.n2181 0.00372581
R25671 dvss.n1333 dvss 0.00372581
R25672 dvss dvss.n2126 0.00372581
R25673 dvss dvss.n5773 0.00372581
R25674 dvss.n5794 dvss 0.00372581
R25675 dvss dvss.n835 0.00372581
R25676 dvss dvss.n826 0.00372581
R25677 dvss.n5916 dvss 0.00372581
R25678 dvss dvss.n6082 0.00372581
R25679 dvss.n5963 dvss 0.00372581
R25680 dvss dvss.n6032 0.00372581
R25681 dvss dvss.n106 0.00372581
R25682 dvss dvss.n97 0.00372581
R25683 dvss.n6805 dvss 0.00372581
R25684 dvss.n6954 dvss 0.00372581
R25685 dvss.n1709 dvss.n1604 0.00366011
R25686 dvss.n1735 dvss.n1608 0.00366011
R25687 dvss dvss.n2167 0.00332258
R25688 dvss.n1613 dvss 0.00330899
R25689 dvss.n1811 dvss 0.00330899
R25690 dvss.n1831 dvss 0.00330899
R25691 dvss.n1926 dvss 0.00330899
R25692 dvss.n1981 dvss 0.00330899
R25693 dvss dvss.n1426 0.00330899
R25694 dvss.n2098 dvss 0.00330899
R25695 dvss dvss.n5705 0.00330899
R25696 dvss dvss.n5694 0.00330899
R25697 dvss dvss.n1073 0.00330899
R25698 dvss.n1114 dvss 0.00330899
R25699 dvss dvss.n776 0.00330899
R25700 dvss.n6201 dvss 0.00330899
R25701 dvss dvss.n733 0.00330899
R25702 dvss dvss.n722 0.00330899
R25703 dvss dvss.n6689 0.00330899
R25704 dvss dvss.n6678 0.00330899
R25705 dvss dvss.n52 0.00330899
R25706 dvss.n6942 dvss 0.00330899
R25707 dvss.n3442 dvss 0.00310417
R25708 dvss.n4705 dvss 0.00310417
R25709 dvss.n3280 dvss 0.00303378
R25710 dvss.n5162 dvss 0.00303378
R25711 dvss.n5201 dvss 0.00303378
R25712 dvss.n5240 dvss 0.00303378
R25713 dvss.n5279 dvss 0.00303378
R25714 dvss.n5536 dvss 0.00303378
R25715 dvss dvss.n6234 0.00303378
R25716 dvss dvss.n6302 0.00303378
R25717 dvss dvss.n6349 0.00303378
R25718 dvss.n6422 dvss 0.00303378
R25719 dvss.n1712 dvss 0.00295787
R25720 dvss.n1734 dvss 0.00295787
R25721 dvss.n1782 dvss.n1553 0.00295787
R25722 dvss.n1517 dvss 0.00295787
R25723 dvss.n1839 dvss 0.00295787
R25724 dvss.n1897 dvss.n1487 0.00295787
R25725 dvss.n1973 dvss 0.00295787
R25726 dvss.n1968 dvss 0.00295787
R25727 dvss.n2061 dvss.n1435 0.00295787
R25728 dvss.n1388 dvss 0.00295787
R25729 dvss.n1374 dvss 0.00295787
R25730 dvss.n5715 dvss.n908 0.00295787
R25731 dvss.n5686 dvss 0.00295787
R25732 dvss dvss.n939 0.00295787
R25733 dvss.n962 dvss.n957 0.00295787
R25734 dvss.n5633 dvss 0.00295787
R25735 dvss.n5628 dvss 0.00295787
R25736 dvss.n6164 dvss.n785 0.00295787
R25737 dvss.n640 dvss 0.00295787
R25738 dvss.n624 dvss 0.00295787
R25739 dvss.n743 dvss.n554 0.00295787
R25740 dvss.n714 dvss 0.00295787
R25741 dvss dvss.n585 0.00295787
R25742 dvss.n6699 dvss.n142 0.00295787
R25743 dvss.n6670 dvss 0.00295787
R25744 dvss.n6665 dvss 0.00295787
R25745 dvss.n6905 dvss.n61 0.00295787
R25746 dvss.n6467 dvss 0.00295787
R25747 dvss.n6453 dvss 0.00295787
R25748 dvss.n2249 dvss 0.00291935
R25749 dvss.n2223 dvss.n1281 0.00291935
R25750 dvss.n2199 dvss 0.00291935
R25751 dvss.n2173 dvss.n1312 0.00291935
R25752 dvss.n2144 dvss 0.00291935
R25753 dvss.n2118 dvss.n1343 0.00291935
R25754 dvss dvss.n5763 0.00291935
R25755 dvss.n5805 dvss.n5804 0.00291935
R25756 dvss.n5852 dvss 0.00291935
R25757 dvss.n5887 dvss.n5886 0.00291935
R25758 dvss.n6100 dvss 0.00291935
R25759 dvss.n6074 dvss.n5942 0.00291935
R25760 dvss.n6050 dvss 0.00291935
R25761 dvss.n6024 dvss.n5973 0.00291935
R25762 dvss.n6746 dvss 0.00291935
R25763 dvss.n6781 dvss.n6780 0.00291935
R25764 dvss.n6841 dvss 0.00291935
R25765 dvss.n6960 dvss.n6958 0.00291935
R25766 dvss dvss.n1613 0.00260674
R25767 dvss.n1785 dvss 0.00260674
R25768 dvss.n1860 dvss.n1517 0.00260674
R25769 dvss.n1910 dvss 0.00260674
R25770 dvss.n1973 dvss.n1948 0.00260674
R25771 dvss.n2074 dvss 0.00260674
R25772 dvss.n1389 dvss.n1388 0.00260674
R25773 dvss dvss.n5710 0.00260674
R25774 dvss.n5686 dvss.n938 0.00260674
R25775 dvss.n1085 dvss 0.00260674
R25776 dvss.n5633 dvss.n1108 0.00260674
R25777 dvss.n6177 dvss 0.00260674
R25778 dvss.n641 dvss.n640 0.00260674
R25779 dvss dvss.n738 0.00260674
R25780 dvss.n714 dvss.n584 0.00260674
R25781 dvss dvss.n6694 0.00260674
R25782 dvss.n6670 dvss.n175 0.00260674
R25783 dvss.n6918 dvss 0.00260674
R25784 dvss.n6468 dvss.n6467 0.00260674
R25785 dvss.n1861 dvss.n1860 0.00190449
R25786 dvss.n1870 dvss.n1509 0.00190449
R25787 dvss.n1970 dvss.n1948 0.00190449
R25788 dvss.n2025 dvss.n2024 0.00190449
R25789 dvss.n1389 dvss.n1369 0.00190449
R25790 dvss.n5727 dvss.n895 0.00190449
R25791 dvss.n5683 dvss.n938 0.00190449
R25792 dvss.n5679 dvss.n5678 0.00190449
R25793 dvss.n5630 dvss.n1108 0.00190449
R25794 dvss.n6128 dvss.n6127 0.00190449
R25795 dvss.n641 dvss.n621 0.00190449
R25796 dvss.n756 dvss.n755 0.00190449
R25797 dvss.n711 dvss.n584 0.00190449
R25798 dvss.n6711 dvss.n129 0.00190449
R25799 dvss.n6667 dvss.n175 0.00190449
R25800 dvss.n6869 dvss.n6868 0.00190449
R25801 dvss.n6468 dvss.n6448 0.00190449
R25802 dvss.n6487 dvss.n6486 0.00190449
R25803 dvss dvss.n884 0.00170968
R25804 dvss dvss.n5816 0.00170968
R25805 dvss.n5900 dvss 0.00170968
R25806 dvss.n1829 dvss.n1533 0.00155337
R25807 dvss dvss.n1865 0.00155337
R25808 dvss.n1942 dvss.n1941 0.00155337
R25809 dvss dvss.n1453 0.00155337
R25810 dvss.n2022 dvss 0.00155337
R25811 dvss.n2095 dvss.n2094 0.00155337
R25812 dvss.n1404 dvss 0.00155337
R25813 dvss.n1406 dvss 0.00155337
R25814 dvss.n5695 dvss.n928 0.00155337
R25815 dvss dvss.n986 0.00155337
R25816 dvss dvss.n943 0.00155337
R25817 dvss.n5644 dvss.n1100 0.00155337
R25818 dvss dvss.n803 0.00155337
R25819 dvss.n6125 dvss 0.00155337
R25820 dvss.n6198 dvss.n6197 0.00155337
R25821 dvss dvss.n538 0.00155337
R25822 dvss.n723 dvss.n574 0.00155337
R25823 dvss.n707 dvss 0.00155337
R25824 dvss.n6679 dvss.n162 0.00155337
R25825 dvss.n6866 dvss 0.00155337
R25826 dvss.n6939 dvss.n6938 0.00155337
R25827 dvss.n6484 dvss 0.00155337
R25828 dvss.n3233 dvss.n3178 0.00134459
R25829 dvss dvss.n3171 0.00134459
R25830 dvss.n5118 dvss.n5117 0.00134459
R25831 dvss.n2273 dvss 0.00130645
R25832 dvss.n1617 dvss 0.00120225
R25833 dvss.n2235 dvss.n1275 0.000903226
R25834 dvss dvss.n2221 0.000903226
R25835 dvss.n2185 dvss.n1306 0.000903226
R25836 dvss dvss.n2171 0.000903226
R25837 dvss.n2130 dvss.n1337 0.000903226
R25838 dvss dvss.n2116 0.000903226
R25839 dvss.n5791 dvss.n5790 0.000903226
R25840 dvss.n5810 dvss 0.000903226
R25841 dvss.n5872 dvss.n825 0.000903226
R25842 dvss dvss.n818 0.000903226
R25843 dvss.n6086 dvss.n5936 0.000903226
R25844 dvss dvss.n6072 0.000903226
R25845 dvss.n6036 dvss.n5967 0.000903226
R25846 dvss dvss.n6022 0.000903226
R25847 dvss.n6766 dvss.n96 0.000903226
R25848 dvss dvss.n89 0.000903226
R25849 dvss.n6827 dvss.n6823 0.000903226
R25850 dvss.n6972 dvss 0.000903226
R25851 dvss.n1702 dvss.n1700 0.000851124
R25852 dvss.n1704 dvss.n1599 0.000851124
R25853 dvss.n1705 dvss.n1600 0.000851124
R25854 dvss.n1706 dvss.n1601 0.000851124
R25855 dvss.n1707 dvss.n1602 0.000851124
R25856 dvss.n1708 dvss.n1603 0.000851124
R25857 dvss.n1712 dvss.n1604 0.000851124
R25858 dvss.n1713 dvss.n1605 0.000851124
R25859 dvss.n1714 dvss.n1606 0.000851124
R25860 dvss.n1618 dvss.n1607 0.000851124
R25861 dvss.n1735 dvss.n1734 0.000851124
R25862 dvss.n1621 dvss.n1620 0.000851124
R25863 dvss.n1759 dvss.n1758 0.000851124
R25864 dvss.n1765 dvss.n1764 0.000851124
R25865 dvss.n1768 dvss.n1563 0.000851124
R25866 dvss.n1767 dvss.n1564 0.000851124
R25867 dvss.n1584 dvss.n1583 0.000851124
R25868 dvss.n1587 dvss.n1585 0.000851124
R25869 dvss.n1827 dvss.n1826 0.000851124
R25870 dvss.n1857 dvss 0.000851124
R25871 dvss.n1939 dvss.n1938 0.000851124
R25872 dvss dvss.n1967 0.000851124
R25873 dvss.n2101 dvss.n1355 0.000851124
R25874 dvss dvss.n1373 0.000851124
R25875 dvss.n5700 dvss.n927 0.000851124
R25876 dvss.n1044 dvss 0.000851124
R25877 dvss.n5645 dvss.n1081 0.000851124
R25878 dvss dvss.n5627 0.000851124
R25879 dvss.n6204 dvss.n532 0.000851124
R25880 dvss.n644 dvss 0.000851124
R25881 dvss.n728 dvss.n573 0.000851124
R25882 dvss.n595 dvss 0.000851124
R25883 dvss.n6684 dvss.n161 0.000851124
R25884 dvss dvss.n6664 0.000851124
R25885 dvss.n6945 dvss.n30 0.000851124
R25886 dvss.n6475 dvss 0.000851124
R25887 porb.n2 porb.n0 243.458
R25888 porb.n2 porb.n1 205.059
R25889 porb.n4 porb.n3 205.059
R25890 porb.n6 porb.n5 205.059
R25891 porb.n8 porb.n7 205.059
R25892 porb.n10 porb.n9 205.059
R25893 porb.n12 porb.n11 205.059
R25894 porb.n14 porb.n13 205.059
R25895 porb.n17 porb.n15 133.534
R25896 porb.n17 porb.n16 99.1759
R25897 porb.n19 porb.n18 99.1759
R25898 porb.n21 porb.n20 99.1759
R25899 porb.n23 porb.n22 99.1759
R25900 porb.n25 porb.n24 99.1759
R25901 porb.n27 porb.n26 99.1759
R25902 porb porb.n28 97.4305
R25903 porb.n4 porb.n2 38.4005
R25904 porb.n6 porb.n4 38.4005
R25905 porb.n8 porb.n6 38.4005
R25906 porb.n10 porb.n8 38.4005
R25907 porb.n12 porb.n10 38.4005
R25908 porb.n14 porb.n12 38.4005
R25909 porb.n19 porb.n17 34.3584
R25910 porb.n21 porb.n19 34.3584
R25911 porb.n23 porb.n21 34.3584
R25912 porb.n25 porb.n23 34.3584
R25913 porb.n27 porb.n25 34.3584
R25914 porb.n29 porb.n27 34.3584
R25915 porb.n30 porb 32.1105
R25916 porb.n13 porb.t25 26.5955
R25917 porb.n13 porb.t23 26.5955
R25918 porb.n0 porb.t29 26.5955
R25919 porb.n0 porb.t18 26.5955
R25920 porb.n1 porb.t17 26.5955
R25921 porb.n1 porb.t31 26.5955
R25922 porb.n3 porb.t30 26.5955
R25923 porb.n3 porb.t19 26.5955
R25924 porb.n5 porb.t28 26.5955
R25925 porb.n5 porb.t24 26.5955
R25926 porb.n7 porb.t16 26.5955
R25927 porb.n7 porb.t22 26.5955
R25928 porb.n9 porb.t21 26.5955
R25929 porb.n9 porb.t27 26.5955
R25930 porb.n11 porb.t20 26.5955
R25931 porb.n11 porb.t26 26.5955
R25932 porb.n28 porb.t5 24.9236
R25933 porb.n28 porb.t3 24.9236
R25934 porb.n15 porb.t9 24.9236
R25935 porb.n15 porb.t14 24.9236
R25936 porb.n16 porb.t13 24.9236
R25937 porb.n16 porb.t11 24.9236
R25938 porb.n18 porb.t10 24.9236
R25939 porb.n18 porb.t15 24.9236
R25940 porb.n20 porb.t8 24.9236
R25941 porb.n20 porb.t4 24.9236
R25942 porb.n22 porb.t12 24.9236
R25943 porb.n22 porb.t2 24.9236
R25944 porb.n24 porb.t1 24.9236
R25945 porb.n24 porb.t7 24.9236
R25946 porb.n26 porb.t0 24.9236
R25947 porb.n26 porb.t6 24.9236
R25948 porb porb.n14 18.4247
R25949 porb.n30 porb.n29 8.33989
R25950 porb porb.n30 3.10353
R25951 porb.n29 porb 1.74595
R25952 vbg_1v2.n55 vbg_1v2.t20 384.709
R25953 vbg_1v2.n54 vbg_1v2.t20 384.709
R25954 vbg_1v2.n65 vbg_1v2.t8 384.226
R25955 vbg_1v2.t8 vbg_1v2.n50 384.226
R25956 vbg_1v2.n64 vbg_1v2.t2 384.226
R25957 vbg_1v2.t2 vbg_1v2.n63 384.226
R25958 vbg_1v2.t9 vbg_1v2.n51 384.226
R25959 vbg_1v2.n62 vbg_1v2.t9 384.226
R25960 vbg_1v2.t5 vbg_1v2.n60 384.226
R25961 vbg_1v2.n61 vbg_1v2.t5 384.226
R25962 vbg_1v2.n59 vbg_1v2.t32 384.226
R25963 vbg_1v2.t32 vbg_1v2.n52 384.226
R25964 vbg_1v2.n58 vbg_1v2.t22 384.226
R25965 vbg_1v2.t22 vbg_1v2.n57 384.226
R25966 vbg_1v2.t18 vbg_1v2.n53 384.226
R25967 vbg_1v2.n56 vbg_1v2.t18 384.226
R25968 vbg_1v2.t23 vbg_1v2.n54 384.226
R25969 vbg_1v2.n55 vbg_1v2.t23 384.226
R25970 vbg_1v2.t28 vbg_1v2.n66 384.226
R25971 vbg_1v2.n67 vbg_1v2.t28 384.226
R25972 vbg_1v2.n1 vbg_1v2.n0 92.8573
R25973 vbg_1v2.n49 vbg_1v2.n48 48.1045
R25974 vbg_1v2 vbg_1v2.n17 18.13
R25975 vbg_1v2.n0 vbg_1v2.t0 16.5305
R25976 vbg_1v2.n0 vbg_1v2.t1 16.5305
R25977 vbg_1v2.n47 vbg_1v2.t11 14.8978
R25978 vbg_1v2.n46 vbg_1v2.t11 14.8978
R25979 vbg_1v2.n43 vbg_1v2.t33 14.8978
R25980 vbg_1v2.n42 vbg_1v2.t33 14.8978
R25981 vbg_1v2.n39 vbg_1v2.t26 14.8978
R25982 vbg_1v2.n38 vbg_1v2.t26 14.8978
R25983 vbg_1v2.n35 vbg_1v2.t13 14.8978
R25984 vbg_1v2.n34 vbg_1v2.t13 14.8978
R25985 vbg_1v2.n31 vbg_1v2.t38 14.8978
R25986 vbg_1v2.n30 vbg_1v2.t38 14.8978
R25987 vbg_1v2.n27 vbg_1v2.t14 14.8978
R25988 vbg_1v2.n26 vbg_1v2.t14 14.8978
R25989 vbg_1v2.n23 vbg_1v2.t39 14.8978
R25990 vbg_1v2.n22 vbg_1v2.t39 14.8978
R25991 vbg_1v2.n19 vbg_1v2.t27 14.8978
R25992 vbg_1v2.t27 vbg_1v2.n18 14.8978
R25993 vbg_1v2.t4 vbg_1v2.n46 12.9902
R25994 vbg_1v2.n47 vbg_1v2.t4 12.9902
R25995 vbg_1v2.t29 vbg_1v2.n42 12.9902
R25996 vbg_1v2.n43 vbg_1v2.t29 12.9902
R25997 vbg_1v2.t17 vbg_1v2.n38 12.9902
R25998 vbg_1v2.n39 vbg_1v2.t17 12.9902
R25999 vbg_1v2.t6 vbg_1v2.n34 12.9902
R26000 vbg_1v2.n35 vbg_1v2.t6 12.9902
R26001 vbg_1v2.t30 vbg_1v2.n30 12.9902
R26002 vbg_1v2.n31 vbg_1v2.t30 12.9902
R26003 vbg_1v2.t7 vbg_1v2.n26 12.9902
R26004 vbg_1v2.n27 vbg_1v2.t7 12.9902
R26005 vbg_1v2.t31 vbg_1v2.n22 12.9902
R26006 vbg_1v2.n23 vbg_1v2.t31 12.9902
R26007 vbg_1v2.t19 vbg_1v2.n18 12.9902
R26008 vbg_1v2.n19 vbg_1v2.t19 12.9902
R26009 vbg_1v2.n17 vbg_1v2.n1 12.0156
R26010 vbg_1v2.n9 vbg_1v2.t25 9.72783
R26011 vbg_1v2.n2 vbg_1v2.t16 9.65028
R26012 vbg_1v2.n16 vbg_1v2.n8 8.96563
R26013 vbg_1v2.n15 vbg_1v2.t40 8.73727
R26014 vbg_1v2.n14 vbg_1v2.t21 8.73727
R26015 vbg_1v2.n13 vbg_1v2.t41 8.73727
R26016 vbg_1v2.n12 vbg_1v2.t10 8.73727
R26017 vbg_1v2.n11 vbg_1v2.t42 8.73727
R26018 vbg_1v2.n10 vbg_1v2.t24 8.73727
R26019 vbg_1v2.n9 vbg_1v2.t43 8.73727
R26020 vbg_1v2.n8 vbg_1v2.t34 8.65985
R26021 vbg_1v2.n7 vbg_1v2.t12 8.65985
R26022 vbg_1v2.n6 vbg_1v2.t35 8.65985
R26023 vbg_1v2.n5 vbg_1v2.t3 8.65985
R26024 vbg_1v2.n4 vbg_1v2.t36 8.65985
R26025 vbg_1v2.n3 vbg_1v2.t15 8.65985
R26026 vbg_1v2.n2 vbg_1v2.t37 8.65985
R26027 vbg_1v2.n16 vbg_1v2.n15 5.98511
R26028 vbg_1v2.n1 vbg_1v2 5.30666
R26029 vbg_1v2.n20 vbg_1v2.n18 5.24569
R26030 vbg_1v2.n20 vbg_1v2.n19 4.5005
R26031 vbg_1v2.n22 vbg_1v2.n21 4.5005
R26032 vbg_1v2.n24 vbg_1v2.n23 4.5005
R26033 vbg_1v2.n26 vbg_1v2.n25 4.5005
R26034 vbg_1v2.n28 vbg_1v2.n27 4.5005
R26035 vbg_1v2.n30 vbg_1v2.n29 4.5005
R26036 vbg_1v2.n32 vbg_1v2.n31 4.5005
R26037 vbg_1v2.n34 vbg_1v2.n33 4.5005
R26038 vbg_1v2.n36 vbg_1v2.n35 4.5005
R26039 vbg_1v2.n38 vbg_1v2.n37 4.5005
R26040 vbg_1v2.n40 vbg_1v2.n39 4.5005
R26041 vbg_1v2.n42 vbg_1v2.n41 4.5005
R26042 vbg_1v2.n44 vbg_1v2.n43 4.5005
R26043 vbg_1v2.n46 vbg_1v2.n45 4.5005
R26044 vbg_1v2.n48 vbg_1v2.n47 4.5005
R26045 vbg_1v2.n66 vbg_1v2.n49 4.5005
R26046 vbg_1v2.n68 vbg_1v2.n67 4.5005
R26047 vbg_1v2.n17 vbg_1v2.n16 4.39202
R26048 vbg_1v2.n68 vbg_1v2.n49 2.63992
R26049 vbg_1v2.n15 vbg_1v2.n14 0.99106
R26050 vbg_1v2.n14 vbg_1v2.n13 0.99106
R26051 vbg_1v2.n13 vbg_1v2.n12 0.99106
R26052 vbg_1v2.n12 vbg_1v2.n11 0.99106
R26053 vbg_1v2.n11 vbg_1v2.n10 0.99106
R26054 vbg_1v2.n10 vbg_1v2.n9 0.99106
R26055 vbg_1v2.n8 vbg_1v2.n7 0.99093
R26056 vbg_1v2.n7 vbg_1v2.n6 0.99093
R26057 vbg_1v2.n6 vbg_1v2.n5 0.99093
R26058 vbg_1v2.n5 vbg_1v2.n4 0.99093
R26059 vbg_1v2.n4 vbg_1v2.n3 0.99093
R26060 vbg_1v2.n3 vbg_1v2.n2 0.99093
R26061 vbg_1v2.n48 vbg_1v2.n45 0.745692
R26062 vbg_1v2.n44 vbg_1v2.n41 0.745692
R26063 vbg_1v2.n40 vbg_1v2.n37 0.745692
R26064 vbg_1v2.n36 vbg_1v2.n33 0.745692
R26065 vbg_1v2.n32 vbg_1v2.n29 0.745692
R26066 vbg_1v2.n28 vbg_1v2.n25 0.745692
R26067 vbg_1v2.n24 vbg_1v2.n21 0.745692
R26068 vbg_1v2.n56 vbg_1v2.n55 0.484196
R26069 vbg_1v2.n57 vbg_1v2.n56 0.484196
R26070 vbg_1v2.n57 vbg_1v2.n52 0.484196
R26071 vbg_1v2.n61 vbg_1v2.n52 0.484196
R26072 vbg_1v2.n62 vbg_1v2.n61 0.484196
R26073 vbg_1v2.n63 vbg_1v2.n62 0.484196
R26074 vbg_1v2.n63 vbg_1v2.n50 0.484196
R26075 vbg_1v2.n54 vbg_1v2.n53 0.484196
R26076 vbg_1v2.n58 vbg_1v2.n53 0.484196
R26077 vbg_1v2.n59 vbg_1v2.n58 0.484196
R26078 vbg_1v2.n60 vbg_1v2.n59 0.484196
R26079 vbg_1v2.n60 vbg_1v2.n51 0.484196
R26080 vbg_1v2.n64 vbg_1v2.n51 0.484196
R26081 vbg_1v2.n65 vbg_1v2.n64 0.484196
R26082 vbg_1v2.n67 vbg_1v2.n50 0.459739
R26083 vbg_1v2.n66 vbg_1v2.n65 0.459739
R26084 vbg_1v2.n45 vbg_1v2.n44 0.260115
R26085 vbg_1v2.n41 vbg_1v2.n40 0.260115
R26086 vbg_1v2.n37 vbg_1v2.n36 0.260115
R26087 vbg_1v2.n33 vbg_1v2.n32 0.260115
R26088 vbg_1v2.n29 vbg_1v2.n28 0.260115
R26089 vbg_1v2.n25 vbg_1v2.n24 0.260115
R26090 vbg_1v2.n21 vbg_1v2.n20 0.260115
R26091 vbg_1v2 vbg_1v2.n68 0.063
R26092 por_dig_0.clknet_1_1__leaf_osc_ck.n48 por_dig_0.clknet_1_1__leaf_osc_ck.n46 333.392
R26093 por_dig_0.clknet_1_1__leaf_osc_ck.n54 por_dig_0.clknet_1_1__leaf_osc_ck.n42 301.392
R26094 por_dig_0.clknet_1_1__leaf_osc_ck.n53 por_dig_0.clknet_1_1__leaf_osc_ck.n43 301.392
R26095 por_dig_0.clknet_1_1__leaf_osc_ck.n52 por_dig_0.clknet_1_1__leaf_osc_ck.n44 301.392
R26096 por_dig_0.clknet_1_1__leaf_osc_ck.n51 por_dig_0.clknet_1_1__leaf_osc_ck.n45 301.392
R26097 por_dig_0.clknet_1_1__leaf_osc_ck.n48 por_dig_0.clknet_1_1__leaf_osc_ck.n47 301.392
R26098 por_dig_0.clknet_1_1__leaf_osc_ck.n50 por_dig_0.clknet_1_1__leaf_osc_ck.n49 301.392
R26099 por_dig_0.clknet_1_1__leaf_osc_ck.n55 por_dig_0.clknet_1_1__leaf_osc_ck.n41 297.863
R26100 por_dig_0.clknet_1_1__leaf_osc_ck.n18 por_dig_0.clknet_1_1__leaf_osc_ck.t34 294.557
R26101 por_dig_0.clknet_1_1__leaf_osc_ck.n14 por_dig_0.clknet_1_1__leaf_osc_ck.t41 294.557
R26102 por_dig_0.clknet_1_1__leaf_osc_ck.n12 por_dig_0.clknet_1_1__leaf_osc_ck.t35 294.557
R26103 por_dig_0.clknet_1_1__leaf_osc_ck.n10 por_dig_0.clknet_1_1__leaf_osc_ck.t49 294.557
R26104 por_dig_0.clknet_1_1__leaf_osc_ck.n33 por_dig_0.clknet_1_1__leaf_osc_ck.t42 294.557
R26105 por_dig_0.clknet_1_1__leaf_osc_ck.n29 por_dig_0.clknet_1_1__leaf_osc_ck.t45 294.557
R26106 por_dig_0.clknet_1_1__leaf_osc_ck.n21 por_dig_0.clknet_1_1__leaf_osc_ck.t37 294.557
R26107 por_dig_0.clknet_1_1__leaf_osc_ck.n25 por_dig_0.clknet_1_1__leaf_osc_ck.t38 294.557
R26108 por_dig_0.clknet_1_1__leaf_osc_ck.n23 por_dig_0.clknet_1_1__leaf_osc_ck.t48 294.557
R26109 por_dig_0.clknet_1_1__leaf_osc_ck.n2 por_dig_0.clknet_1_1__leaf_osc_ck.n0 248.638
R26110 por_dig_0.clknet_1_1__leaf_osc_ck.n18 por_dig_0.clknet_1_1__leaf_osc_ck.t39 211.01
R26111 por_dig_0.clknet_1_1__leaf_osc_ck.n14 por_dig_0.clknet_1_1__leaf_osc_ck.t32 211.01
R26112 por_dig_0.clknet_1_1__leaf_osc_ck.n12 por_dig_0.clknet_1_1__leaf_osc_ck.t40 211.01
R26113 por_dig_0.clknet_1_1__leaf_osc_ck.n10 por_dig_0.clknet_1_1__leaf_osc_ck.t36 211.01
R26114 por_dig_0.clknet_1_1__leaf_osc_ck.n33 por_dig_0.clknet_1_1__leaf_osc_ck.t47 211.01
R26115 por_dig_0.clknet_1_1__leaf_osc_ck.n29 por_dig_0.clknet_1_1__leaf_osc_ck.t46 211.01
R26116 por_dig_0.clknet_1_1__leaf_osc_ck.n21 por_dig_0.clknet_1_1__leaf_osc_ck.t43 211.01
R26117 por_dig_0.clknet_1_1__leaf_osc_ck.n25 por_dig_0.clknet_1_1__leaf_osc_ck.t44 211.01
R26118 por_dig_0.clknet_1_1__leaf_osc_ck.n23 por_dig_0.clknet_1_1__leaf_osc_ck.t33 211.01
R26119 por_dig_0.clknet_1_1__leaf_osc_ck.n2 por_dig_0.clknet_1_1__leaf_osc_ck.n1 203.463
R26120 por_dig_0.clknet_1_1__leaf_osc_ck.n4 por_dig_0.clknet_1_1__leaf_osc_ck.n3 203.463
R26121 por_dig_0.clknet_1_1__leaf_osc_ck.n8 por_dig_0.clknet_1_1__leaf_osc_ck.n7 203.463
R26122 por_dig_0.clknet_1_1__leaf_osc_ck.n40 por_dig_0.clknet_1_1__leaf_osc_ck.n39 203.463
R26123 por_dig_0.clknet_1_1__leaf_osc_ck.n6 por_dig_0.clknet_1_1__leaf_osc_ck.n5 202.456
R26124 por_dig_0.clknet_1_1__leaf_osc_ck por_dig_0.clknet_1_1__leaf_osc_ck.n57 199.607
R26125 por_dig_0.clknet_1_1__leaf_osc_ck.n37 por_dig_0.clknet_1_1__leaf_osc_ck.n9 188.201
R26126 por_dig_0.clknet_1_1__leaf_osc_ck por_dig_0.clknet_1_1__leaf_osc_ck.n21 156.207
R26127 por_dig_0.clknet_1_1__leaf_osc_ck.n19 por_dig_0.clknet_1_1__leaf_osc_ck.n18 153.097
R26128 por_dig_0.clknet_1_1__leaf_osc_ck.n11 por_dig_0.clknet_1_1__leaf_osc_ck.n10 153.097
R26129 por_dig_0.clknet_1_1__leaf_osc_ck.n34 por_dig_0.clknet_1_1__leaf_osc_ck.n33 153.097
R26130 por_dig_0.clknet_1_1__leaf_osc_ck.n26 por_dig_0.clknet_1_1__leaf_osc_ck.n25 153.097
R26131 por_dig_0.clknet_1_1__leaf_osc_ck.n15 por_dig_0.clknet_1_1__leaf_osc_ck.n14 152
R26132 por_dig_0.clknet_1_1__leaf_osc_ck.n13 por_dig_0.clknet_1_1__leaf_osc_ck.n12 152
R26133 por_dig_0.clknet_1_1__leaf_osc_ck.n30 por_dig_0.clknet_1_1__leaf_osc_ck.n29 152
R26134 por_dig_0.clknet_1_1__leaf_osc_ck.n24 por_dig_0.clknet_1_1__leaf_osc_ck.n23 152
R26135 por_dig_0.clknet_1_1__leaf_osc_ck.n4 por_dig_0.clknet_1_1__leaf_osc_ck.n2 45.177
R26136 por_dig_0.clknet_1_1__leaf_osc_ck.n38 por_dig_0.clknet_1_1__leaf_osc_ck.n8 45.177
R26137 por_dig_0.clknet_1_1__leaf_osc_ck.n40 por_dig_0.clknet_1_1__leaf_osc_ck.n38 45.177
R26138 por_dig_0.clknet_1_1__leaf_osc_ck.n6 por_dig_0.clknet_1_1__leaf_osc_ck.n4 44.0476
R26139 por_dig_0.clknet_1_1__leaf_osc_ck.n8 por_dig_0.clknet_1_1__leaf_osc_ck.n6 44.0476
R26140 por_dig_0.clknet_1_1__leaf_osc_ck.n0 por_dig_0.clknet_1_1__leaf_osc_ck.t8 40.0005
R26141 por_dig_0.clknet_1_1__leaf_osc_ck.n0 por_dig_0.clknet_1_1__leaf_osc_ck.t14 40.0005
R26142 por_dig_0.clknet_1_1__leaf_osc_ck.n1 por_dig_0.clknet_1_1__leaf_osc_ck.t11 40.0005
R26143 por_dig_0.clknet_1_1__leaf_osc_ck.n1 por_dig_0.clknet_1_1__leaf_osc_ck.t0 40.0005
R26144 por_dig_0.clknet_1_1__leaf_osc_ck.n3 por_dig_0.clknet_1_1__leaf_osc_ck.t13 40.0005
R26145 por_dig_0.clknet_1_1__leaf_osc_ck.n3 por_dig_0.clknet_1_1__leaf_osc_ck.t4 40.0005
R26146 por_dig_0.clknet_1_1__leaf_osc_ck.n5 por_dig_0.clknet_1_1__leaf_osc_ck.t1 40.0005
R26147 por_dig_0.clknet_1_1__leaf_osc_ck.n5 por_dig_0.clknet_1_1__leaf_osc_ck.t6 40.0005
R26148 por_dig_0.clknet_1_1__leaf_osc_ck.n7 por_dig_0.clknet_1_1__leaf_osc_ck.t2 40.0005
R26149 por_dig_0.clknet_1_1__leaf_osc_ck.n7 por_dig_0.clknet_1_1__leaf_osc_ck.t7 40.0005
R26150 por_dig_0.clknet_1_1__leaf_osc_ck.n9 por_dig_0.clknet_1_1__leaf_osc_ck.t3 40.0005
R26151 por_dig_0.clknet_1_1__leaf_osc_ck.n9 por_dig_0.clknet_1_1__leaf_osc_ck.t9 40.0005
R26152 por_dig_0.clknet_1_1__leaf_osc_ck.n39 por_dig_0.clknet_1_1__leaf_osc_ck.t5 40.0005
R26153 por_dig_0.clknet_1_1__leaf_osc_ck.n39 por_dig_0.clknet_1_1__leaf_osc_ck.t10 40.0005
R26154 por_dig_0.clknet_1_1__leaf_osc_ck.n57 por_dig_0.clknet_1_1__leaf_osc_ck.t12 40.0005
R26155 por_dig_0.clknet_1_1__leaf_osc_ck.n57 por_dig_0.clknet_1_1__leaf_osc_ck.t15 40.0005
R26156 por_dig_0.clknet_1_1__leaf_osc_ck.n54 por_dig_0.clknet_1_1__leaf_osc_ck.n53 32.0005
R26157 por_dig_0.clknet_1_1__leaf_osc_ck.n53 por_dig_0.clknet_1_1__leaf_osc_ck.n52 32.0005
R26158 por_dig_0.clknet_1_1__leaf_osc_ck.n50 por_dig_0.clknet_1_1__leaf_osc_ck.n48 32.0005
R26159 por_dig_0.clknet_1_1__leaf_osc_ck.n51 por_dig_0.clknet_1_1__leaf_osc_ck.n50 32.0005
R26160 por_dig_0.clknet_1_1__leaf_osc_ck.n52 por_dig_0.clknet_1_1__leaf_osc_ck.n51 31.2005
R26161 por_dig_0.clknet_1_1__leaf_osc_ck.n42 por_dig_0.clknet_1_1__leaf_osc_ck.t23 27.5805
R26162 por_dig_0.clknet_1_1__leaf_osc_ck.n42 por_dig_0.clknet_1_1__leaf_osc_ck.t28 27.5805
R26163 por_dig_0.clknet_1_1__leaf_osc_ck.n41 por_dig_0.clknet_1_1__leaf_osc_ck.t30 27.5805
R26164 por_dig_0.clknet_1_1__leaf_osc_ck.n41 por_dig_0.clknet_1_1__leaf_osc_ck.t17 27.5805
R26165 por_dig_0.clknet_1_1__leaf_osc_ck.n43 por_dig_0.clknet_1_1__leaf_osc_ck.t21 27.5805
R26166 por_dig_0.clknet_1_1__leaf_osc_ck.n43 por_dig_0.clknet_1_1__leaf_osc_ck.t27 27.5805
R26167 por_dig_0.clknet_1_1__leaf_osc_ck.n44 por_dig_0.clknet_1_1__leaf_osc_ck.t20 27.5805
R26168 por_dig_0.clknet_1_1__leaf_osc_ck.n44 por_dig_0.clknet_1_1__leaf_osc_ck.t25 27.5805
R26169 por_dig_0.clknet_1_1__leaf_osc_ck.n45 por_dig_0.clknet_1_1__leaf_osc_ck.t19 27.5805
R26170 por_dig_0.clknet_1_1__leaf_osc_ck.n45 por_dig_0.clknet_1_1__leaf_osc_ck.t24 27.5805
R26171 por_dig_0.clknet_1_1__leaf_osc_ck.n46 por_dig_0.clknet_1_1__leaf_osc_ck.t26 27.5805
R26172 por_dig_0.clknet_1_1__leaf_osc_ck.n46 por_dig_0.clknet_1_1__leaf_osc_ck.t16 27.5805
R26173 por_dig_0.clknet_1_1__leaf_osc_ck.n47 por_dig_0.clknet_1_1__leaf_osc_ck.t29 27.5805
R26174 por_dig_0.clknet_1_1__leaf_osc_ck.n47 por_dig_0.clknet_1_1__leaf_osc_ck.t18 27.5805
R26175 por_dig_0.clknet_1_1__leaf_osc_ck.n49 por_dig_0.clknet_1_1__leaf_osc_ck.t31 27.5805
R26176 por_dig_0.clknet_1_1__leaf_osc_ck.n49 por_dig_0.clknet_1_1__leaf_osc_ck.t22 27.5805
R26177 por_dig_0.clknet_1_1__leaf_osc_ck.n27 por_dig_0.clknet_1_1__leaf_osc_ck 25.5892
R26178 por_dig_0.clknet_1_1__leaf_osc_ck.n32 por_dig_0.clknet_1_1__leaf_osc_ck.n28 21.6653
R26179 por_dig_0.clknet_1_1__leaf_osc_ck.n17 por_dig_0.clknet_1_1__leaf_osc_ck.n11 16.3913
R26180 por_dig_0.clknet_1_1__leaf_osc_ck.n28 por_dig_0.clknet_1_1__leaf_osc_ck.n22 15.4901
R26181 por_dig_0.clknet_1_1__leaf_osc_ck.n38 por_dig_0.clknet_1_1__leaf_osc_ck.n37 15.262
R26182 por_dig_0.clknet_1_1__leaf_osc_ck.n20 por_dig_0.clknet_1_1__leaf_osc_ck.n19 14.916
R26183 por_dig_0.clknet_1_1__leaf_osc_ck.n36 por_dig_0.clknet_1_1__leaf_osc_ck.n35 14.1296
R26184 por_dig_0.clknet_1_1__leaf_osc_ck.n32 por_dig_0.clknet_1_1__leaf_osc_ck.n31 13.8005
R26185 por_dig_0.clknet_1_1__leaf_osc_ck.n27 por_dig_0.clknet_1_1__leaf_osc_ck.n26 13.8005
R26186 por_dig_0.clknet_1_1__leaf_osc_ck.n56 por_dig_0.clknet_1_1__leaf_osc_ck.n40 13.177
R26187 por_dig_0.clknet_1_1__leaf_osc_ck.n16 por_dig_0.clknet_1_1__leaf_osc_ck 12.7032
R26188 por_dig_0.clknet_1_1__leaf_osc_ck.n16 por_dig_0.clknet_1_1__leaf_osc_ck 12.4091
R26189 por_dig_0.clknet_1_1__leaf_osc_ck.n55 por_dig_0.clknet_1_1__leaf_osc_ck.n54 10.4484
R26190 por_dig_0.clknet_1_1__leaf_osc_ck por_dig_0.clknet_1_1__leaf_osc_ck.n15 10.4234
R26191 por_dig_0.clknet_1_1__leaf_osc_ck por_dig_0.clknet_1_1__leaf_osc_ck.n13 10.4234
R26192 por_dig_0.clknet_1_1__leaf_osc_ck por_dig_0.clknet_1_1__leaf_osc_ck.n24 10.4234
R26193 por_dig_0.clknet_1_1__leaf_osc_ck.n35 por_dig_0.clknet_1_1__leaf_osc_ck.n32 9.99634
R26194 por_dig_0.clknet_1_1__leaf_osc_ck.n31 por_dig_0.clknet_1_1__leaf_osc_ck 9.32621
R26195 por_dig_0.clknet_1_1__leaf_osc_ck.n22 por_dig_0.clknet_1_1__leaf_osc_ck 9.32621
R26196 por_dig_0.clknet_1_1__leaf_osc_ck.n35 por_dig_0.clknet_1_1__leaf_osc_ck.n34 9.3005
R26197 por_dig_0.clknet_1_1__leaf_osc_ck.n37 por_dig_0.clknet_1_1__leaf_osc_ck.n36 9.3005
R26198 por_dig_0.clknet_1_1__leaf_osc_ck.n36 por_dig_0.clknet_1_1__leaf_osc_ck.n20 5.88649
R26199 por_dig_0.clknet_1_1__leaf_osc_ck.n17 por_dig_0.clknet_1_1__leaf_osc_ck.n16 4.5005
R26200 por_dig_0.clknet_1_1__leaf_osc_ck.n56 por_dig_0.clknet_1_1__leaf_osc_ck 3.13183
R26201 por_dig_0.clknet_1_1__leaf_osc_ck.n19 por_dig_0.clknet_1_1__leaf_osc_ck 3.10907
R26202 por_dig_0.clknet_1_1__leaf_osc_ck.n11 por_dig_0.clknet_1_1__leaf_osc_ck 3.10907
R26203 por_dig_0.clknet_1_1__leaf_osc_ck.n34 por_dig_0.clknet_1_1__leaf_osc_ck 3.10907
R26204 por_dig_0.clknet_1_1__leaf_osc_ck.n22 por_dig_0.clknet_1_1__leaf_osc_ck 3.10907
R26205 por_dig_0.clknet_1_1__leaf_osc_ck.n26 por_dig_0.clknet_1_1__leaf_osc_ck 3.10907
R26206 por_dig_0.clknet_1_1__leaf_osc_ck.n20 por_dig_0.clknet_1_1__leaf_osc_ck.n17 2.2972
R26207 por_dig_0.clknet_1_1__leaf_osc_ck por_dig_0.clknet_1_1__leaf_osc_ck.n27 2.21135
R26208 por_dig_0.clknet_1_1__leaf_osc_ck.n15 por_dig_0.clknet_1_1__leaf_osc_ck 2.01193
R26209 por_dig_0.clknet_1_1__leaf_osc_ck.n13 por_dig_0.clknet_1_1__leaf_osc_ck 2.01193
R26210 por_dig_0.clknet_1_1__leaf_osc_ck.n30 por_dig_0.clknet_1_1__leaf_osc_ck 2.01193
R26211 por_dig_0.clknet_1_1__leaf_osc_ck.n24 por_dig_0.clknet_1_1__leaf_osc_ck 2.01193
R26212 por_dig_0.clknet_1_1__leaf_osc_ck por_dig_0.clknet_1_1__leaf_osc_ck.n55 1.75844
R26213 por_dig_0.clknet_1_1__leaf_osc_ck.n31 por_dig_0.clknet_1_1__leaf_osc_ck.n30 1.09764
R26214 por_dig_0.clknet_1_1__leaf_osc_ck por_dig_0.clknet_1_1__leaf_osc_ck.n56 0.604792
R26215 por_dig_0.clknet_1_1__leaf_osc_ck.n28 por_dig_0.clknet_1_1__leaf_osc_ck 0.389923
R26216 por_dig_0.net22 por_dig_0.net22.n29 617.727
R26217 por_dig_0.net22.t11 por_dig_0.net22.t6 395.01
R26218 por_dig_0.net22 por_dig_0.net22.t11 320.745
R26219 por_dig_0.net22.n8 por_dig_0.net22.t5 261.887
R26220 por_dig_0.net22.n15 por_dig_0.net22.t23 254.256
R26221 por_dig_0.net22.n3 por_dig_0.net22.t4 241.536
R26222 por_dig_0.net22.n5 por_dig_0.net22.t18 241.536
R26223 por_dig_0.net22.n19 por_dig_0.net22.t16 241.536
R26224 por_dig_0.net22.n10 por_dig_0.net22.t20 241.536
R26225 por_dig_0.net22.n13 por_dig_0.net22.t9 239.505
R26226 por_dig_0.net22.n22 por_dig_0.net22.t19 230.155
R26227 por_dig_0.net22.n1 por_dig_0.net22.t21 229.369
R26228 por_dig_0.net22 por_dig_0.net22.n0 222.863
R26229 por_dig_0.net22.n15 por_dig_0.net22.t15 181.956
R26230 por_dig_0.net22.n3 por_dig_0.net22.t14 169.237
R26231 por_dig_0.net22.n5 por_dig_0.net22.t7 169.237
R26232 por_dig_0.net22.n19 por_dig_0.net22.t10 169.237
R26233 por_dig_0.net22.n10 por_dig_0.net22.t13 169.237
R26234 por_dig_0.net22.n13 por_dig_0.net22.t17 167.204
R26235 por_dig_0.net22.n6 por_dig_0.net22.n5 159.952
R26236 por_dig_0.net22.n20 por_dig_0.net22.n19 159.758
R26237 por_dig_0.net22.n22 por_dig_0.net22.t8 157.856
R26238 por_dig_0.net22.n1 por_dig_0.net22.t12 157.07
R26239 por_dig_0.net22.n8 por_dig_0.net22.t22 155.847
R26240 por_dig_0.net22.n2 por_dig_0.net22.n1 153.66
R26241 por_dig_0.net22.n14 por_dig_0.net22.n13 153.601
R26242 por_dig_0.net22.n23 por_dig_0.net22.n22 153.147
R26243 por_dig_0.net22.n9 por_dig_0.net22.n8 153.13
R26244 por_dig_0.net22.n16 por_dig_0.net22.n15 152.357
R26245 por_dig_0.net22.n4 por_dig_0.net22.n3 152
R26246 por_dig_0.net22.n11 por_dig_0.net22.n10 152
R26247 por_dig_0.net22.n0 por_dig_0.net22.t0 38.5719
R26248 por_dig_0.net22.n0 por_dig_0.net22.t1 38.5719
R26249 por_dig_0.net22.n29 por_dig_0.net22.t2 26.5955
R26250 por_dig_0.net22.n29 por_dig_0.net22.t3 26.5955
R26251 por_dig_0.net22.n27 por_dig_0.net22 25.7976
R26252 por_dig_0.net22.n17 por_dig_0.net22.n14 19.1121
R26253 por_dig_0.net22.n21 por_dig_0.net22.n20 14.5053
R26254 por_dig_0.net22.n17 por_dig_0.net22.n16 14.2892
R26255 por_dig_0.net22.n7 por_dig_0.net22 14.1918
R26256 por_dig_0.net22 por_dig_0.net22.n4 14.0693
R26257 por_dig_0.net22.n27 por_dig_0.net22 12.5005
R26258 por_dig_0.net22.n18 por_dig_0.net22.n12 11.9527
R26259 por_dig_0.net22.n12 por_dig_0.net22 11.4531
R26260 por_dig_0.net22.n28 por_dig_0.net22 11.3034
R26261 por_dig_0.net22.n26 por_dig_0.net22.n7 10.2027
R26262 por_dig_0.net22.n28 por_dig_0.net22 9.6005
R26263 por_dig_0.net22 por_dig_0.net22.n2 9.55096
R26264 por_dig_0.net22.n21 por_dig_0.net22.n18 9.40156
R26265 por_dig_0.net22.n24 por_dig_0.net22.n23 9.3005
R26266 por_dig_0.net22.n25 por_dig_0.net22.n9 9.3005
R26267 por_dig_0.net22.n18 por_dig_0.net22.n17 8.76698
R26268 por_dig_0.net22.n24 por_dig_0.net22.n21 7.10077
R26269 por_dig_0.net22 por_dig_0.net22.n27 5.29514
R26270 por_dig_0.net22.n7 por_dig_0.net22 4.73093
R26271 por_dig_0.net22.n2 por_dig_0.net22 4.26717
R26272 por_dig_0.net22.n14 por_dig_0.net22 3.8405
R26273 por_dig_0.net22 por_dig_0.net22.n6 3.33963
R26274 por_dig_0.net22.n6 por_dig_0.net22 3.29747
R26275 por_dig_0.net22.n23 por_dig_0.net22 3.24826
R26276 por_dig_0.net22.n9 por_dig_0.net22 3.2005
R26277 por_dig_0.net22.n20 por_dig_0.net22 3.10353
R26278 por_dig_0.net22.n16 por_dig_0.net22 3.02272
R26279 por_dig_0.net22.n27 por_dig_0.net22.n26 2.88099
R26280 por_dig_0.net22 por_dig_0.net22.n28 2.82403
R26281 por_dig_0.net22.n11 por_dig_0.net22 2.47068
R26282 por_dig_0.net22.n4 por_dig_0.net22 2.3087
R26283 por_dig_0.net22.n26 por_dig_0.net22.n25 2.19246
R26284 por_dig_0.net22.n12 por_dig_0.net22.n11 1.34787
R26285 por_dig_0.net22.n25 por_dig_0.net22.n24 1.11605
R26286 avss.n158 avss.n134 2.18688e+07
R26287 avss.n71 avss.n70 188352
R26288 avss.n896 avss.n860 160432
R26289 avss.n859 avss.n858 110146
R26290 avss.n133 avss.n50 100279
R26291 avss.n1019 avss.n50 100279
R26292 avss.n133 avss.n51 100279
R26293 avss.n1019 avss.n51 100279
R26294 avss.n70 avss.n69 92956.3
R26295 avss.n399 avss.n159 68021.9
R26296 avss.n1003 avss.n64 64733.3
R26297 avss.n70 avss.t298 48414.6
R26298 avss.n885 avss.n61 45524.4
R26299 avss.n885 avss.n62 45524.4
R26300 avss.n1005 avss.n61 45524.4
R26301 avss.n1005 avss.n62 45524.4
R26302 avss.n591 avss.n587 45524.4
R26303 avss.n791 avss.n587 45524.4
R26304 avss.n790 avss.n591 45524.4
R26305 avss.n791 avss.n790 45524.4
R26306 avss.n399 avss.n398 45183
R26307 avss.n1102 avss.n8 37415.6
R26308 avss.n1003 avss.n1002 29160.7
R26309 avss.n860 avss.t145 29031.2
R26310 avss.n1022 avss.n47 21059.4
R26311 avss.n1022 avss.n48 21059.4
R26312 avss.n1024 avss.n47 21059.4
R26313 avss.n1024 avss.n48 21059.4
R26314 avss.n988 avss.n73 18174.6
R26315 avss.n995 avss.n73 18174.6
R26316 avss.n995 avss.n72 18174.6
R26317 avss.n988 avss.n72 18174.6
R26318 avss.n842 avss.n567 18174.6
R26319 avss.n814 avss.n567 18174.6
R26320 avss.n842 avss.n841 18174.6
R26321 avss.n841 avss.n814 18174.6
R26322 avss.n857 avss.n578 17601.7
R26323 avss.n156 avss.n118 16300.9
R26324 avss.n403 avss.n118 16300.9
R26325 avss.n156 avss.n120 16300.9
R26326 avss.n403 avss.n120 16300.9
R26327 avss.n897 avss.n896 13864
R26328 avss.n208 avss.n159 12588.9
R26329 avss.n894 avss.n862 12517.1
R26330 avss.n888 avss.n862 12517.1
R26331 avss.n888 avss.n861 12517.1
R26332 avss.n894 avss.n861 12517.1
R26333 avss.n455 avss.n451 7742.83
R26334 avss.n457 avss.n451 7742.83
R26335 avss.n456 avss.n455 7742.83
R26336 avss.n457 avss.n456 7742.83
R26337 avss.n875 avss.n19 7610.36
R26338 avss.n875 avss.n20 7610.36
R26339 avss.n1079 avss.n20 7610.36
R26340 avss.n1079 avss.n19 7610.36
R26341 avss.n860 avss.n859 7383.98
R26342 avss.n54 avss.n52 6515.58
R26343 avss.n1018 avss.n52 6515.58
R26344 avss.n1017 avss.n54 6515.58
R26345 avss.n1018 avss.n1017 6515.58
R26346 avss.n1082 avss.n12 5644.38
R26347 avss.n1082 avss.n13 5644.38
R26348 avss.n1093 avss.n13 5644.38
R26349 avss.n1093 avss.n12 5644.38
R26350 avss.n159 avss.n158 4523.98
R26351 avss.n454 avss.n449 4175.68
R26352 avss.n458 avss.n449 4175.68
R26353 avss.n454 avss.n450 4175.68
R26354 avss.n458 avss.n450 4175.68
R26355 avss.n982 avss.n80 4139.43
R26356 avss.n978 avss.n80 4139.43
R26357 avss.n982 avss.n81 4139.43
R26358 avss.n978 avss.n81 4139.43
R26359 avss.n846 avss.n807 4139.43
R26360 avss.n812 avss.n807 4139.43
R26361 avss.n812 avss.n808 4139.43
R26362 avss.n846 avss.n808 4139.43
R26363 avss.n575 avss.n571 3978.07
R26364 avss.n575 avss.n572 3978.07
R26365 avss.n900 avss.n572 3978.07
R26366 avss.n900 avss.n571 3978.07
R26367 avss.n1001 avss.n66 3978.07
R26368 avss.n997 avss.n66 3978.07
R26369 avss.n997 avss.n65 3978.07
R26370 avss.n1001 avss.n65 3978.07
R26371 avss.t292 avss.t68 3966.94
R26372 avss.t294 avss.t292 3966.94
R26373 avss.t290 avss.t288 3966.94
R26374 avss.t288 avss.t64 3966.94
R26375 avss.n859 avss.n857 3945.98
R26376 avss.n1096 avss.n9 3902.33
R26377 avss.n1096 avss.n10 3902.33
R26378 avss.n1100 avss.n10 3902.33
R26379 avss.n1100 avss.n9 3902.33
R26380 avss.n896 avss.n895 3318.88
R26381 avss.n401 avss.n400 2998.14
R26382 avss.n1006 avss.n60 2957.93
R26383 avss.n792 avss.n585 2957.93
R26384 avss.n590 avss.n586 2957.93
R26385 avss.n792 avss.n586 2957.93
R26386 avss.n590 avss.n588 2940.24
R26387 avss.n884 avss.n60 2935.34
R26388 avss.n220 avss.n219 2905.02
R26389 avss.n232 avss.n231 2905.02
R26390 avss.n244 avss.n243 2905.02
R26391 avss.n256 avss.n255 2905.02
R26392 avss.n268 avss.n267 2905.02
R26393 avss.n280 avss.n279 2905.02
R26394 avss.n292 avss.n291 2905.02
R26395 avss.n304 avss.n303 2905.02
R26396 avss.n316 avss.n315 2905.02
R26397 avss.n328 avss.n327 2905.02
R26398 avss.n340 avss.n339 2905.02
R26399 avss.n352 avss.n351 2905.02
R26400 avss.n364 avss.n363 2905.02
R26401 avss.n376 avss.n375 2905.02
R26402 avss.n388 avss.n387 2905.02
R26403 avss.n1104 avss.n1103 2538.7
R26404 avss.t14 avss.n807 2436.62
R26405 avss.n808 avss.t145 2436.62
R26406 avss.n80 avss.t278 2436.62
R26407 avss.n1025 avss.n45 2366.87
R26408 avss.n1025 avss.n44 2366.87
R26409 avss.n1021 avss.n44 2344.28
R26410 avss.n1021 avss.n45 2344.28
R26411 avss.n843 avss.t68 2304.08
R26412 avss.t64 avss.n576 2304.08
R26413 avss.n501 avss.n485 2087.09
R26414 avss.n526 avss.n475 2084.98
R26415 avss.n839 avss.n566 2054.02
R26416 avss.n904 avss.n566 2054.02
R26417 avss.n994 avss.n74 2054.02
R26418 avss.n989 avss.n74 2054.02
R26419 avss.n519 avss.n517 2039.85
R26420 avss.n543 avss.n542 2039.84
R26421 avss.n840 avss.t294 1983.47
R26422 avss.n840 avss.t290 1983.47
R26423 avss.n904 avss.n903 1894.78
R26424 avss.n839 avss.n815 1894.78
R26425 avss.n991 avss.n989 1894.78
R26426 avss.n994 avss.n993 1894.78
R26427 avss.n404 avss.n117 1813.84
R26428 avss.n1106 avss.n6 1735.47
R26429 avss.n1107 avss.n6 1735.47
R26430 avss.n1107 avss.n5 1735.47
R26431 avss.n1106 avss.n5 1735.47
R26432 avss.t274 avss.n49 1637.21
R26433 avss.n154 avss.n153 1602.64
R26434 avss.n878 avss.n877 1487.81
R26435 avss.n877 avss.n58 1487.81
R26436 avss.n884 avss.n878 1439.24
R26437 avss.n1006 avss.n58 1439.24
R26438 avss.n889 avss.n874 1435.48
R26439 avss.n889 avss.n873 1435.48
R26440 avss.n400 avss.n132 1414.29
R26441 avss.t42 avss.t104 1389.88
R26442 avss.n893 avss.n864 1385.79
R26443 avss.n893 avss.n863 1385.79
R26444 avss.n845 avss.t18 1301
R26445 avss.n845 avss.t24 1301
R26446 avss.n983 avss.t276 1301
R26447 avss.t270 avss.n983 1301
R26448 avss.n1002 avss.t104 1143.92
R26449 avss.t24 avss.t16 1081.77
R26450 avss.t278 avss.t272 1081.77
R26451 avss.t20 avss.t14 1081.77
R26452 avss.t10 avss.t20 1081.77
R26453 avss.t12 avss.t10 1081.77
R26454 avss.t18 avss.t12 1081.77
R26455 avss.t16 avss.t22 1081.77
R26456 avss.t22 avss.t147 1081.77
R26457 avss.t272 avss.t268 1081.77
R26458 avss.t268 avss.t280 1081.77
R26459 avss.n453 avss.n446 976.942
R26460 avss.n453 avss.n452 976.942
R26461 avss.n460 avss.n459 976.188
R26462 avss.n459 avss.n448 974.683
R26463 avss.t296 avss.n49 964.784
R26464 avss.n400 avss.n399 939.895
R26465 avss.n813 avss.t18 925.769
R26466 avss.t24 avss.n813 925.769
R26467 avss.n844 avss.t145 887.293
R26468 avss.n1078 avss.n21 874.542
R26469 avss.n22 avss.n21 874.542
R26470 avss.n219 avss.n205 815.444
R26471 avss.n231 avss.n202 815.444
R26472 avss.n243 avss.n199 815.444
R26473 avss.n255 avss.n196 815.444
R26474 avss.n267 avss.n193 815.444
R26475 avss.n279 avss.n190 815.444
R26476 avss.n291 avss.n187 815.444
R26477 avss.n303 avss.n184 815.444
R26478 avss.n315 avss.n181 815.444
R26479 avss.n327 avss.n178 815.444
R26480 avss.n339 avss.n175 815.444
R26481 avss.n351 avss.n172 815.444
R26482 avss.n363 avss.n169 815.444
R26483 avss.n375 avss.n166 815.444
R26484 avss.n387 avss.n163 815.444
R26485 avss.n398 avss.n160 815.444
R26486 avss.n115 avss.n114 796.612
R26487 avss.n119 avss.n115 782.683
R26488 avss.n124 avss.n121 769.572
R26489 avss.n1076 avss.n1075 765.741
R26490 avss.n1077 avss.n1076 765.741
R26491 avss.n406 avss.n405 759.718
R26492 avss.n208 avss.t394 755.986
R26493 avss.n220 avss.t212 755.986
R26494 avss.n232 avss.t300 755.986
R26495 avss.n244 avss.t329 755.986
R26496 avss.n256 avss.t8 755.986
R26497 avss.n268 avss.t263 755.986
R26498 avss.n280 avss.t317 755.986
R26499 avss.n292 avss.t219 755.986
R26500 avss.n304 avss.t227 755.986
R26501 avss.n316 avss.t371 755.986
R26502 avss.n328 avss.t261 755.986
R26503 avss.n340 avss.t376 755.986
R26504 avss.n352 avss.t239 755.986
R26505 avss.n364 avss.t3 755.986
R26506 avss.n376 avss.t32 755.986
R26507 avss.n388 avss.t307 755.986
R26508 avss.t387 avss.t380 731.963
R26509 avss.t254 avss.t252 731.963
R26510 avss.t252 avss.n898 684.673
R26511 avss.n899 avss.t380 668.225
R26512 avss.n1092 avss.n14 649.788
R26513 avss.n1083 avss.n14 649.788
R26514 avss.n1004 avss.n1003 627.813
R26515 avss.n518 avss.t119 625.516
R26516 avss.n525 avss.t119 625.516
R26517 avss.t119 avss.n469 614.321
R26518 avss.n536 avss.t119 614.321
R26519 avss.n858 avss.t387 602.431
R26520 avss.n406 avss.n116 598.966
R26521 avss.t119 avss.n508 598.606
R26522 avss.n509 avss.t119 598.606
R26523 avss.n494 avss.t119 588.343
R26524 avss.n492 avss.t119 588.343
R26525 avss.n515 avss.n514 585
R26526 avss.n513 avss.n482 585
R26527 avss.n482 avss.n481 585
R26528 avss.n512 avss.n511 585
R26529 avss.n511 avss.n510 585
R26530 avss.n484 avss.n483 585
R26531 avss.n509 avss.n484 585
R26532 avss.n507 avss.n506 585
R26533 avss.n508 avss.n507 585
R26534 avss.n505 avss.n486 585
R26535 avss.n486 avss.n485 585
R26536 avss.n504 avss.n503 585
R26537 avss.n488 avss.n487 585
R26538 avss.n530 avss.n529 585
R26539 avss.n527 avss.n477 585
R26540 avss.n527 avss.n526 585
R26541 avss.n524 avss.n523 585
R26542 avss.n525 avss.n524 585
R26543 avss.n522 avss.n478 585
R26544 avss.n518 avss.n478 585
R26545 avss.n521 avss.n520 585
R26546 avss.n520 avss.n519 585
R26547 avss.n480 avss.n479 585
R26548 avss.n531 avss.n476 585
R26549 avss.n533 avss.n532 585
R26550 avss.n534 avss.n533 585
R26551 avss.n474 avss.n473 585
R26552 avss.n535 avss.n474 585
R26553 avss.n538 avss.n537 585
R26554 avss.n537 avss.n536 585
R26555 avss.n539 avss.n471 585
R26556 avss.n471 avss.n469 585
R26557 avss.n541 avss.n540 585
R26558 avss.n542 avss.n541 585
R26559 avss.n472 avss.n470 585
R26560 avss.n466 avss.n464 585
R26561 avss.n499 avss.n498 585
R26562 avss.n500 avss.n499 585
R26563 avss.n497 avss.n490 585
R26564 avss.n490 avss.n489 585
R26565 avss.n496 avss.n495 585
R26566 avss.n495 avss.n494 585
R26567 avss.n493 avss.n491 585
R26568 avss.n493 avss.n492 585
R26569 avss.n465 avss.n463 585
R26570 avss.n467 avss.n465 585
R26571 avss.n546 avss.n545 585
R26572 avss.n545 avss.n544 585
R26573 avss.n649 avss.n648 585
R26574 avss.n648 avss.n647 585
R26575 avss.n655 avss.n654 585
R26576 avss.n656 avss.n655 585
R26577 avss.n646 avss.n645 585
R26578 avss.n657 avss.n646 585
R26579 avss.n661 avss.n660 585
R26580 avss.n660 avss.n659 585
R26581 avss.n641 avss.n640 585
R26582 avss.n658 avss.n640 585
R26583 avss.n669 avss.n668 585
R26584 avss.n670 avss.n669 585
R26585 avss.n638 avss.n636 585
R26586 avss.n671 avss.n638 585
R26587 avss.n676 avss.n675 585
R26588 avss.n675 avss.n674 585
R26589 avss.n639 avss.n637 585
R26590 avss.n673 avss.n639 585
R26591 avss.n632 avss.n631 585
R26592 avss.n672 avss.n631 585
R26593 avss.n689 avss.n688 585
R26594 avss.n690 avss.n689 585
R26595 avss.n630 avss.n629 585
R26596 avss.n691 avss.n630 585
R26597 avss.n695 avss.n694 585
R26598 avss.n694 avss.n693 585
R26599 avss.n625 avss.n624 585
R26600 avss.n692 avss.n624 585
R26601 avss.n710 avss.n709 585
R26602 avss.n711 avss.n710 585
R26603 avss.n708 avss.n622 585
R26604 avss.n712 avss.n622 585
R26605 avss.n714 avss.n623 585
R26606 avss.n714 avss.n713 585
R26607 avss.n715 avss.n621 585
R26608 avss.n716 avss.n715 585
R26609 avss.n720 avss.n719 585
R26610 avss.n719 avss.n718 585
R26611 avss.n619 avss.n618 585
R26612 avss.n717 avss.n618 585
R26613 avss.n730 avss.n729 585
R26614 avss.n731 avss.n730 585
R26615 avss.n617 avss.n616 585
R26616 avss.n732 avss.n617 585
R26617 avss.n736 avss.n735 585
R26618 avss.n735 avss.n734 585
R26619 avss.n612 avss.n611 585
R26620 avss.n733 avss.n611 585
R26621 avss.n744 avss.n743 585
R26622 avss.n745 avss.n744 585
R26623 avss.n610 avss.n609 585
R26624 avss.n746 avss.n610 585
R26625 avss.n750 avss.n749 585
R26626 avss.n749 avss.n748 585
R26627 avss.n606 avss.n605 585
R26628 avss.n747 avss.n605 585
R26629 avss.n758 avss.n757 585
R26630 avss.n759 avss.n758 585
R26631 avss.n604 avss.n603 585
R26632 avss.n760 avss.n604 585
R26633 avss.n764 avss.n763 585
R26634 avss.n763 avss.n762 585
R26635 avss.n600 avss.n599 585
R26636 avss.n761 avss.n599 585
R26637 avss.n774 avss.n773 585
R26638 avss.n775 avss.n774 585
R26639 avss.n598 avss.n597 585
R26640 avss.n776 avss.n598 585
R26641 avss.n779 avss.n778 585
R26642 avss.n778 avss.n777 585
R26643 avss.n594 avss.n593 585
R26644 avss.n593 avss.n592 585
R26645 avss.n787 avss.n786 585
R26646 avss.n788 avss.n787 585
R26647 avss.n581 avss.n580 585
R26648 avss.n580 avss.n579 585
R26649 avss.n855 avss.n854 585
R26650 avss.n856 avss.n855 585
R26651 avss.n131 avss.n130 585
R26652 avss.n132 avss.n131 585
R26653 avss.n123 avss.n122 585
R26654 avss.n210 avss.n209 585
R26655 avss.n209 avss.n208 585
R26656 avss.n207 avss.n206 585
R26657 avss.n206 avss.n205 585
R26658 avss.n218 avss.n217 585
R26659 avss.n219 avss.n218 585
R26660 avss.n222 avss.n221 585
R26661 avss.n221 avss.n220 585
R26662 avss.n204 avss.n203 585
R26663 avss.n203 avss.n202 585
R26664 avss.n230 avss.n229 585
R26665 avss.n231 avss.n230 585
R26666 avss.n234 avss.n233 585
R26667 avss.n233 avss.n232 585
R26668 avss.n201 avss.n200 585
R26669 avss.n200 avss.n199 585
R26670 avss.n242 avss.n241 585
R26671 avss.n243 avss.n242 585
R26672 avss.n246 avss.n245 585
R26673 avss.n245 avss.n244 585
R26674 avss.n198 avss.n197 585
R26675 avss.n197 avss.n196 585
R26676 avss.n254 avss.n253 585
R26677 avss.n255 avss.n254 585
R26678 avss.n258 avss.n257 585
R26679 avss.n257 avss.n256 585
R26680 avss.n195 avss.n194 585
R26681 avss.n194 avss.n193 585
R26682 avss.n266 avss.n265 585
R26683 avss.n267 avss.n266 585
R26684 avss.n270 avss.n269 585
R26685 avss.n269 avss.n268 585
R26686 avss.n192 avss.n191 585
R26687 avss.n191 avss.n190 585
R26688 avss.n278 avss.n277 585
R26689 avss.n279 avss.n278 585
R26690 avss.n282 avss.n281 585
R26691 avss.n281 avss.n280 585
R26692 avss.n189 avss.n188 585
R26693 avss.n188 avss.n187 585
R26694 avss.n290 avss.n289 585
R26695 avss.n291 avss.n290 585
R26696 avss.n294 avss.n293 585
R26697 avss.n293 avss.n292 585
R26698 avss.n186 avss.n185 585
R26699 avss.n185 avss.n184 585
R26700 avss.n302 avss.n301 585
R26701 avss.n303 avss.n302 585
R26702 avss.n306 avss.n305 585
R26703 avss.n305 avss.n304 585
R26704 avss.n183 avss.n182 585
R26705 avss.n182 avss.n181 585
R26706 avss.n314 avss.n313 585
R26707 avss.n315 avss.n314 585
R26708 avss.n318 avss.n317 585
R26709 avss.n317 avss.n316 585
R26710 avss.n180 avss.n179 585
R26711 avss.n179 avss.n178 585
R26712 avss.n326 avss.n325 585
R26713 avss.n327 avss.n326 585
R26714 avss.n330 avss.n329 585
R26715 avss.n329 avss.n328 585
R26716 avss.n177 avss.n176 585
R26717 avss.n176 avss.n175 585
R26718 avss.n338 avss.n337 585
R26719 avss.n339 avss.n338 585
R26720 avss.n342 avss.n341 585
R26721 avss.n341 avss.n340 585
R26722 avss.n174 avss.n173 585
R26723 avss.n173 avss.n172 585
R26724 avss.n350 avss.n349 585
R26725 avss.n351 avss.n350 585
R26726 avss.n354 avss.n353 585
R26727 avss.n353 avss.n352 585
R26728 avss.n171 avss.n170 585
R26729 avss.n170 avss.n169 585
R26730 avss.n362 avss.n361 585
R26731 avss.n363 avss.n362 585
R26732 avss.n366 avss.n365 585
R26733 avss.n365 avss.n364 585
R26734 avss.n168 avss.n167 585
R26735 avss.n167 avss.n166 585
R26736 avss.n374 avss.n373 585
R26737 avss.n375 avss.n374 585
R26738 avss.n378 avss.n377 585
R26739 avss.n377 avss.n376 585
R26740 avss.n165 avss.n164 585
R26741 avss.n164 avss.n163 585
R26742 avss.n386 avss.n385 585
R26743 avss.n387 avss.n386 585
R26744 avss.n390 avss.n389 585
R26745 avss.n389 avss.n388 585
R26746 avss.n162 avss.n161 585
R26747 avss.n161 avss.n160 585
R26748 avss.n397 avss.n396 585
R26749 avss.n398 avss.n397 585
R26750 avss.n1084 avss.n15 540.989
R26751 avss.n1091 avss.n15 540.989
R26752 avss.n389 avss.n161 539.294
R26753 avss.n397 avss.n161 539.294
R26754 avss.n377 avss.n164 539.294
R26755 avss.n386 avss.n164 539.294
R26756 avss.n365 avss.n167 539.294
R26757 avss.n374 avss.n167 539.294
R26758 avss.n353 avss.n170 539.294
R26759 avss.n362 avss.n170 539.294
R26760 avss.n341 avss.n173 539.294
R26761 avss.n350 avss.n173 539.294
R26762 avss.n329 avss.n176 539.294
R26763 avss.n338 avss.n176 539.294
R26764 avss.n317 avss.n179 539.294
R26765 avss.n326 avss.n179 539.294
R26766 avss.n305 avss.n182 539.294
R26767 avss.n314 avss.n182 539.294
R26768 avss.n293 avss.n185 539.294
R26769 avss.n302 avss.n185 539.294
R26770 avss.n281 avss.n188 539.294
R26771 avss.n290 avss.n188 539.294
R26772 avss.n269 avss.n191 539.294
R26773 avss.n278 avss.n191 539.294
R26774 avss.n257 avss.n194 539.294
R26775 avss.n266 avss.n194 539.294
R26776 avss.n245 avss.n197 539.294
R26777 avss.n254 avss.n197 539.294
R26778 avss.n233 avss.n200 539.294
R26779 avss.n242 avss.n200 539.294
R26780 avss.n221 avss.n203 539.294
R26781 avss.n230 avss.n203 539.294
R26782 avss.n209 avss.n206 539.294
R26783 avss.n218 avss.n206 539.294
R26784 avss.n655 avss.n648 539.294
R26785 avss.n655 avss.n646 539.294
R26786 avss.n660 avss.n646 539.294
R26787 avss.n660 avss.n640 539.294
R26788 avss.n669 avss.n640 539.294
R26789 avss.n669 avss.n638 539.294
R26790 avss.n675 avss.n638 539.294
R26791 avss.n675 avss.n639 539.294
R26792 avss.n639 avss.n631 539.294
R26793 avss.n689 avss.n631 539.294
R26794 avss.n689 avss.n630 539.294
R26795 avss.n694 avss.n630 539.294
R26796 avss.n694 avss.n624 539.294
R26797 avss.n710 avss.n624 539.294
R26798 avss.n710 avss.n622 539.294
R26799 avss.n714 avss.n622 539.294
R26800 avss.n715 avss.n714 539.294
R26801 avss.n719 avss.n715 539.294
R26802 avss.n719 avss.n618 539.294
R26803 avss.n730 avss.n618 539.294
R26804 avss.n730 avss.n617 539.294
R26805 avss.n735 avss.n617 539.294
R26806 avss.n735 avss.n611 539.294
R26807 avss.n744 avss.n611 539.294
R26808 avss.n744 avss.n610 539.294
R26809 avss.n749 avss.n610 539.294
R26810 avss.n749 avss.n605 539.294
R26811 avss.n758 avss.n605 539.294
R26812 avss.n758 avss.n604 539.294
R26813 avss.n763 avss.n604 539.294
R26814 avss.n763 avss.n599 539.294
R26815 avss.n774 avss.n599 539.294
R26816 avss.n774 avss.n598 539.294
R26817 avss.n778 avss.n598 539.294
R26818 avss.n778 avss.n593 539.294
R26819 avss.n787 avss.n593 539.294
R26820 avss.n787 avss.n580 539.294
R26821 avss.n855 avss.n580 539.294
R26822 avss.n131 avss.n122 539.294
R26823 avss.n400 avss.t385 492.382
R26824 avss.n79 avss.t42 488.039
R26825 avss.n811 avss.n806 477.741
R26826 avss.n847 avss.n806 477.741
R26827 avss.n980 avss.n979 477.741
R26828 avss.n981 avss.n980 477.741
R26829 avss.t256 avss.n897 474.954
R26830 avss.n901 avss.n570 459.295
R26831 avss.n574 avss.n570 459.295
R26832 avss.n574 avss.n573 459.295
R26833 avss.n1000 avss.n67 459.295
R26834 avss.n1000 avss.n999 459.295
R26835 avss.n999 avss.n998 459.295
R26836 avss.n495 avss.n493 456.416
R26837 avss.n537 avss.n471 456.416
R26838 avss.n524 avss.n478 456.416
R26839 avss.n507 avss.n484 456.416
R26840 avss.n1099 avss.n11 425.264
R26841 avss.n1097 avss.n11 420.43
R26842 avss.n1098 avss.n1097 420.43
R26843 avss.n1099 avss.n1098 420.43
R26844 avss.n848 avss.n805 401.812
R26845 avss.n810 avss.n805 401.812
R26846 avss.n83 avss.n82 401.812
R26847 avss.n977 avss.n83 401.812
R26848 avss.n25 avss.t39 392.769
R26849 avss.n24 avss.t70 392.692
R26850 avss.n23 avss.t97 392.664
R26851 avss.n136 avss.t72 384.515
R26852 avss.n137 avss.t86 384.515
R26853 avss.n138 avss.t50 384.515
R26854 avss.n139 avss.t108 384.515
R26855 avss.n140 avss.t122 384.515
R26856 avss.n142 avss.t113 384.515
R26857 avss.n144 avss.t59 384.515
R26858 avss.n145 avss.t93 384.515
R26859 avss.n146 avss.t120 384.515
R26860 avss.n147 avss.t124 384.515
R26861 avss.n148 avss.t84 384.515
R26862 avss.n150 avss.t61 384.515
R26863 avss.n151 avss.t134 384.515
R26864 avss.n141 avss.t78 384.454
R26865 avss.n149 avss.t48 384.454
R26866 avss.n886 avss.t150 382.757
R26867 avss.n519 avss.n518 363.548
R26868 avss.n526 avss.n525 363.548
R26869 avss.n542 avss.n469 357.041
R26870 avss.n536 avss.n535 357.041
R26871 avss.n535 avss.n534 357.041
R26872 avss.n534 avss.n475 357.041
R26873 avss.n508 avss.n485 347.908
R26874 avss.n510 avss.n509 347.908
R26875 avss.n510 avss.n481 347.908
R26876 avss.n517 avss.n481 347.908
R26877 avss.n501 avss.n500 341.943
R26878 avss.n500 avss.n489 341.943
R26879 avss.n494 avss.n489 341.943
R26880 avss.n492 avss.n467 341.943
R26881 avss.n544 avss.n467 341.943
R26882 avss.n544 avss.n543 341.943
R26883 avss.n844 avss.n843 340.805
R26884 avss.n64 avss.t27 338.375
R26885 avss.n431 avss.n418 333.334
R26886 avss.n426 avss.n425 333.334
R26887 avss.n441 avss.n416 333.334
R26888 avss.t28 avss.n7 323.332
R26889 avss.t28 avss.n1104 323.332
R26890 avss.n902 avss.n569 318.495
R26891 avss.n990 avss.n68 318.495
R26892 avss.n400 avss.n7 301.202
R26893 avss.n528 avss.n475 283.521
R26894 avss.n517 avss.n516 283.521
R26895 avss.n405 avss.n404 274.072
R26896 avss.n155 avss.n114 270.683
R26897 avss.n895 avss.t55 262.885
R26898 avss.n887 avss.t55 262.885
R26899 avss.n502 avss.n501 262.719
R26900 avss.n543 avss.n468 262.719
R26901 avss.n1004 avss.t81 239.365
R26902 avss.n155 avss.n154 238.306
R26903 avss.n898 avss.n576 227.298
R26904 avss.t34 avss.n11 209.756
R26905 avss.n1098 avss.t34 209.756
R26906 avss.n119 avss.n116 208.189
R26907 avss.n1105 avss.n4 202.918
R26908 avss.n1108 avss.n4 202.918
R26909 avss.n132 avss.n121 200.215
R26910 avss.t147 avss.n844 194.476
R26911 avss.n1105 avss.n3 193.918
R26912 avss.n876 avss.t81 188.975
R26913 avss.n1109 avss.n1108 186.73
R26914 avss.t362 avss.t232 185.605
R26915 avss.t232 avss.t223 185.605
R26916 avss.t223 avss.t369 185.605
R26917 avss.t369 avss.t216 185.605
R26918 avss.t216 avss.t162 185.605
R26919 avss.t162 avss.t306 185.605
R26920 avss.t306 avss.t363 185.605
R26921 avss.t363 avss.t156 185.605
R26922 avss.n436 avss.n435 185
R26923 avss.n437 avss.n423 185
R26924 avss.n429 avss.n428 185
R26925 avss.n430 avss.n418 185
R26926 avss.t118 avss.n418 185
R26927 avss.n432 avss.n431 185
R26928 avss.n434 avss.n433 185
R26929 avss.n425 avss.n424 185
R26930 avss.n427 avss.n426 185
R26931 avss.n417 avss.n415 185
R26932 avss.n442 avss.n441 185
R26933 avss.n441 avss.t118 185
R26934 avss.n416 avss.n414 185
R26935 avss.n439 avss.n438 185
R26936 avss.n769 avss.n768 185
R26937 avss.n122 avss.n121 184.572
R26938 avss.n755 avss.t144 163.472
R26939 avss.t408 avss.t158 160.929
R26940 avss.t235 avss.t408 160.929
R26941 avss.t356 avss.t235 160.929
R26942 avss.t365 avss.t356 160.929
R26943 avss.t159 avss.t365 160.929
R26944 avss.t375 avss.t321 160.929
R26945 avss.t321 avss.t164 160.929
R26946 avss.t164 avss.t354 160.929
R26947 avss.t409 avss.t166 160.339
R26948 avss.t245 avss.t409 160.339
R26949 avss.t353 avss.t245 160.339
R26950 avss.t177 avss.t353 160.339
R26951 avss.t250 avss.t225 160.339
R26952 avss.t225 avss.t169 160.339
R26953 avss.t169 avss.t249 160.339
R26954 avss.t249 avss.t26 160.339
R26955 avss.t26 avss.t357 160.339
R26956 avss.t357 avss.t154 160.339
R26957 avss.t154 avss.t236 160.339
R26958 avss.t236 avss.t355 160.339
R26959 avss.t355 avss.t246 160.339
R26960 avss.t246 avss.t285 160.339
R26961 avss.n903 avss.n568 159.248
R26962 avss.n815 avss.n568 159.248
R26963 avss.n992 avss.n991 159.248
R26964 avss.n993 avss.n992 159.248
R26965 avss.n860 avss.n577 157.524
R26966 avss.n158 avss.t177 157.37
R26967 avss.n393 avss.t308 149.067
R26968 avss.n382 avss.t33 149.067
R26969 avss.n370 avss.t4 149.067
R26970 avss.n358 avss.t240 149.067
R26971 avss.n346 avss.t377 149.067
R26972 avss.n334 avss.t262 149.067
R26973 avss.n322 avss.t372 149.067
R26974 avss.n310 avss.t228 149.067
R26975 avss.n298 avss.t220 149.067
R26976 avss.n286 avss.t318 149.067
R26977 avss.n274 avss.t264 149.067
R26978 avss.n262 avss.t9 149.067
R26979 avss.n250 avss.t330 149.067
R26980 avss.n238 avss.t301 149.067
R26981 avss.n226 avss.t213 149.067
R26982 avss.n214 avss.t395 149.067
R26983 avss.n851 avss.t231 149.067
R26984 avss.n782 avss.t138 149.067
R26985 avss.n128 avss.t386 149.067
R26986 avss.n402 avss.t224 142.101
R26987 avss.n401 avss.t362 132.919
R26988 avss.n499 avss.n490 132.635
R26989 avss.n495 avss.n490 132.635
R26990 avss.n493 avss.n465 132.635
R26991 avss.n545 avss.n465 132.635
R26992 avss.n541 avss.n470 132.635
R26993 avss.n541 avss.n471 132.635
R26994 avss.n537 avss.n474 132.635
R26995 avss.n533 avss.n474 132.635
R26996 avss.n533 avss.n476 132.635
R26997 avss.n520 avss.n480 132.635
R26998 avss.n520 avss.n478 132.635
R26999 avss.n527 avss.n524 132.635
R27000 avss.n529 avss.n527 132.635
R27001 avss.n503 avss.n486 132.635
R27002 avss.n507 avss.n486 132.635
R27003 avss.n511 avss.n484 132.635
R27004 avss.n511 avss.n482 132.635
R27005 avss.n515 avss.n482 132.635
R27006 avss.n753 avss.t207 126.32
R27007 avss.n930 avss.t429 125.388
R27008 avss.n651 avss.t183 124.695
R27009 avss.n931 avss.t431 124.674
R27010 avss.n930 avss.t432 124.674
R27011 avss.n932 avss.t103 123.24
R27012 avss.n932 avss.t41 122.623
R27013 avss.t398 avss.n49 118.332
R27014 avss.t175 avss.t322 118.26
R27015 avss.t322 avss.t136 118.26
R27016 avss.t136 avss.t215 118.26
R27017 avss.t215 avss.t161 118.26
R27018 avss.t161 avss.t304 118.26
R27019 avss.n807 avss.n805 117.001
R27020 avss.n808 avss.n806 117.001
R27021 avss.n571 avss.n570 117.001
R27022 avss.n858 avss.n571 117.001
R27023 avss.n573 avss.n572 117.001
R27024 avss.n897 avss.n572 117.001
R27025 avss.n1001 avss.n1000 117.001
R27026 avss.n1002 avss.n1001 117.001
R27027 avss.n980 avss.n81 117.001
R27028 avss.n81 avss.n71 117.001
R27029 avss.n998 avss.n997 117.001
R27030 avss.n997 avss.n996 117.001
R27031 avss.n83 avss.n80 117.001
R27032 avss.n1106 avss.n1105 117.001
R27033 avss.t28 avss.n1106 117.001
R27034 avss.n1108 avss.n1107 117.001
R27035 avss.n1107 avss.t28 117.001
R27036 avss.n428 avss.n418 113.334
R27037 avss.n441 avss.n417 113.334
R27038 avss.n887 avss.n886 111.906
R27039 avss.t304 avss.t243 110.1
R27040 avss.t352 avss.n578 108.138
R27041 avss.t354 avss.n577 108.138
R27042 avss.t166 avss.n134 107.742
R27043 avss.n857 avss.t375 102.603
R27044 avss.n740 avss.n614 100.05
R27045 avss.n726 avss.n725 100.05
R27046 avss.n704 avss.n703 100.05
R27047 avss.n700 avss.n627 100.05
R27048 avss.n685 avss.n684 100.05
R27049 avss.n679 avss.n634 100.05
R27050 avss.n664 avss.n643 100.05
R27051 avss.n573 avss.n569 99.0123
R27052 avss.n998 avss.n68 99.0123
R27053 avss.n6 avss.n4 97.5005
R27054 avss.n1104 avss.n6 97.5005
R27055 avss.n5 avss.n3 97.5005
R27056 avss.n7 avss.n5 97.5005
R27057 avss.t157 avss.t174 96.6926
R27058 avss.n157 avss.t392 94.5922
R27059 avss.t323 avss.t244 91.065
R27060 avss.n796 avss.t15 88.2028
R27061 avss.n800 avss.t146 88.2028
R27062 avss.n936 avss.t334 88.2028
R27063 avss.n85 avss.t279 88.2028
R27064 avss.n89 avss.t299 88.2028
R27065 avss.n908 avss.t257 88.2028
R27066 avss.n938 avss.t43 87.8727
R27067 avss.n910 avss.t381 87.8727
R27068 avss.n423 avss.n421 87.6787
R27069 avss.n435 avss.n421 87.6787
R27070 avss.n937 avss.t332 87.5075
R27071 avss.n936 avss.t333 87.5075
R27072 avss.n909 avss.t255 87.5075
R27073 avss.n908 avss.t253 87.5075
R27074 avss.n1078 avss.n1077 86.2123
R27075 avss.n1075 avss.n22 86.2123
R27076 avss.n1092 avss.n1091 86.2123
R27077 avss.n1084 avss.n1083 86.2123
R27078 avss.n1110 avss.t29 85.1191
R27079 avss.t243 avss.n1102 84.4142
R27080 avss.n913 avss.t66 82.9912
R27081 avss.n554 avss.t128 82.9912
R27082 avss.n821 avss.t69 82.9912
R27083 avss.t133 avss.n832 82.9912
R27084 avss.t112 avss.n969 82.9912
R27085 avss.t96 avss.n966 82.9912
R27086 avss.n941 avss.t102 82.9912
R27087 avss.n104 avss.t47 82.9912
R27088 avss.n903 avss.n902 82.824
R27089 avss.n815 avss.n569 82.824
R27090 avss.n991 avss.n990 82.824
R27091 avss.n993 avss.n68 82.824
R27092 avss.t248 avss.t325 81.8562
R27093 avss.t118 avss.n419 77.7851
R27094 avss.t118 avss.n420 77.7851
R27095 avss.t309 avss.t320 76.3526
R27096 avss.t393 avss.t135 75.5042
R27097 avss.t210 avss.t211 75.5042
R27098 avss.t62 avss.t303 75.5042
R27099 avss.t302 avss.t49 75.5042
R27100 avss.t327 avss.t328 75.5042
R27101 avss.t85 avss.t7 75.5042
R27102 avss.t7 avss.t6 75.5042
R27103 avss.t125 avss.t266 75.5042
R27104 avss.t265 avss.t121 75.5042
R27105 avss.t316 avss.t315 75.5042
R27106 avss.t94 avss.t222 75.5042
R27107 avss.t221 avss.t60 75.5042
R27108 avss.t226 avss.t229 75.5042
R27109 avss.t114 avss.t374 75.5042
R27110 avss.t373 avss.t79 75.5042
R27111 avss.t79 avss.t260 75.5042
R27112 avss.t259 avss.t123 75.5042
R27113 avss.t379 avss.t378 75.5042
R27114 avss.t109 avss.t237 75.5042
R27115 avss.t238 avss.t51 75.5042
R27116 avss.t87 avss.t31 75.5042
R27117 avss.t30 avss.t73 75.5042
R27118 avss.t310 avss.t309 75.5042
R27119 avss.t160 avss.t259 73.8075
R27120 avss.n1103 avss.t156 73.162
R27121 avss.t170 avss.t125 72.9591
R27122 avss.n1103 avss.t175 71.6444
R27123 avss.n798 avss.n797 70.9775
R27124 avss.n796 avss.n795 70.9775
R27125 avss.n802 avss.n801 70.9775
R27126 avss.n800 avss.n799 70.9775
R27127 avss.n87 avss.n86 70.9775
R27128 avss.n85 avss.n84 70.9775
R27129 avss.n91 avss.n90 70.9775
R27130 avss.n89 avss.n88 70.9775
R27131 avss.n560 avss.n559 70.9612
R27132 avss.n558 avss.n557 70.9612
R27133 avss.n564 avss.n563 70.9612
R27134 avss.n837 avss.n836 70.9612
R27135 avss.n820 avss.n817 70.9612
R27136 avss.n834 avss.n833 70.9612
R27137 avss.n110 avss.n109 70.9612
R27138 avss.n108 avss.n107 70.9612
R27139 avss.n97 avss.n96 70.9612
R27140 avss.n95 avss.n94 70.9612
R27141 avss.n971 avss.n970 70.9612
R27142 avss.n968 avss.n967 70.9612
R27143 avss.t118 avss.n422 70.8113
R27144 avss.t118 avss.n440 70.8113
R27145 avss.t341 avss.t234 70.601
R27146 avss.n435 avss.n434 70.0005
R27147 avss.n439 avss.n423 70.0005
R27148 avss.t328 avss.t1 68.7174
R27149 avss.t151 avss.t152 67.9453
R27150 avss.t153 avss.t151 67.9453
R27151 avss.t150 avss.t153 67.9453
R27152 avss.t374 avss.t0 67.869
R27153 avss.t73 avss.t173 67.0206
R27154 avss.t367 avss.t379 64.4756
R27155 avss.t270 avss.t282 63.8987
R27156 avss.n899 avss.t254 63.7388
R27157 avss.t267 avss.t265 63.6272
R27158 avss.n79 avss.t276 63.1818
R27159 avss.n64 avss.n63 61.8334
R27160 avss.t305 avss.t335 61.3923
R27161 avss.n1095 avss.t37 61.1365
R27162 avss.n1101 avss.t364 60.3691
R27163 avss.n470 avss.n468 59.5655
R27164 avss.n503 avss.n502 59.5655
R27165 avss.n502 avss.n488 59.5655
R27166 avss.n468 avss.n466 59.5655
R27167 avss.t394 avss.n205 59.46
R27168 avss.t212 avss.n202 59.46
R27169 avss.t300 avss.n199 59.46
R27170 avss.t329 avss.n196 59.46
R27171 avss.t8 avss.n193 59.46
R27172 avss.t263 avss.n190 59.46
R27173 avss.t317 avss.n187 59.46
R27174 avss.t219 avss.n184 59.46
R27175 avss.t227 avss.n181 59.46
R27176 avss.t371 avss.n178 59.46
R27177 avss.t261 avss.n175 59.46
R27178 avss.t376 avss.n172 59.46
R27179 avss.t239 avss.n169 59.46
R27180 avss.t3 avss.n166 59.46
R27181 avss.t32 avss.n163 59.46
R27182 avss.t307 avss.n160 59.46
R27183 avss.t49 avss.t366 59.3854
R27184 avss.t229 avss.t360 58.5371
R27185 avss.n857 avss.t159 58.3266
R27186 avss.t31 avss.t155 57.6887
R27187 avss.n869 avss.t110 57.0602
R27188 avss.n985 avss.t296 56.675
R27189 avss.t149 avss.t109 55.1437
R27190 avss.t382 avss.t165 54.4857
R27191 avss.t241 avss.t316 54.2953
R27192 avss.t311 avss.t393 53.4469
R27193 avss.n814 avss.n568 53.1823
R27194 avss.n814 avss.n576 53.1823
R27195 avss.n842 avss.n566 53.1823
R27196 avss.n843 avss.n842 53.1823
R27197 avss.n74 avss.n72 53.1823
R27198 avss.n985 avss.n72 53.1823
R27199 avss.n992 avss.n73 53.1823
R27200 avss.n985 avss.n73 53.1823
R27201 avss.n18 avss.t163 52.9509
R27202 avss.n46 avss.t35 51.9277
R27203 avss.t303 avss.t171 50.0535
R27204 avss.n848 avss.n847 49.8123
R27205 avss.n811 avss.n810 49.8123
R27206 avss.n979 avss.n977 49.8123
R27207 avss.n981 avss.n82 49.8123
R27208 avss.t60 avss.t312 49.2052
R27209 avss.t118 avss.n421 48.6621
R27210 avss.t5 avss.t242 48.3568
R27211 avss.n898 avss.t256 47.2902
R27212 avss.t287 avss.t238 45.8117
R27213 avss.t384 avss.t340 45.5327
R27214 avss.t98 avss.t343 45.5327
R27215 avss.t40 avss.t337 45.5327
R27216 avss.n11 avss.n9 45.0005
R27217 avss.t35 avss.n9 45.0005
R27218 avss.n1098 avss.n10 45.0005
R27219 avss.t35 avss.n10 45.0005
R27220 avss.t361 avss.t94 44.9634
R27221 avss.n986 avss.t274 44.1554
R27222 avss.n984 avss.t298 44.1554
R27223 avss.t172 avss.t210 44.115
R27224 avss.t218 avss.n18 43.7421
R27225 avss.t285 avss.n157 43.6909
R27226 avss.t2 avss.n135 43.6909
R27227 avss.n431 avss.n422 43.3803
R27228 avss.n440 avss.n416 43.3803
R27229 avss.n434 avss.n422 43.3803
R27230 avss.n440 avss.n439 43.3803
R27231 avss.t152 avss.n49 42.7523
R27232 avss.n1081 avss.n1080 42.7189
R27233 avss.n996 avss.n71 42.3223
R27234 avss.t319 avss.t382 42.2073
R27235 avss.n656 avss.n647 40.8713
R27236 avss.n659 avss.n657 40.8713
R27237 avss.n671 avss.n670 40.8713
R27238 avss.n691 avss.n690 40.8713
R27239 avss.n693 avss.n692 40.8713
R27240 avss.n718 avss.n717 40.8713
R27241 avss.n732 avss.n731 40.8713
R27242 avss.n748 avss.n746 40.8713
R27243 avss.n762 avss.n760 40.8713
R27244 avss.n788 avss.n592 40.8713
R27245 avss.n856 avss.n579 40.8713
R27246 avss.t211 avss.t284 40.7216
R27247 avss.t222 avss.t286 39.8732
R27248 avss.n996 avss.t298 39.7462
R27249 avss.n658 avss.t184 39.5941
R27250 avss.t188 avss.n716 39.5941
R27251 avss.n775 avss.t370 39.5941
R27252 avss.n777 avss.t233 39.5941
R27253 avss.t51 avss.t214 39.0249
R27254 avss.n1016 avss.n1015 38.6099
R27255 avss.n1016 avss.n53 38.6076
R27256 avss.n1015 avss.n1014 38.5956
R27257 avss.t143 avss.n759 37.8912
R27258 avss.t230 avss.n788 37.8912
R27259 avss.n711 avss.t200 37.0397
R27260 avss.t206 avss.n747 37.0397
R27261 avss.n759 avss.t359 37.0397
R27262 avss.t158 avss.n856 37.0397
R27263 avss.t214 avss.t2 36.4798
R27264 avss.t174 avss.n1101 36.324
R27265 avss.n390 avss.n162 36.1417
R27266 avss.n396 avss.n162 36.1417
R27267 avss.n378 avss.n165 36.1417
R27268 avss.n385 avss.n165 36.1417
R27269 avss.n366 avss.n168 36.1417
R27270 avss.n373 avss.n168 36.1417
R27271 avss.n354 avss.n171 36.1417
R27272 avss.n361 avss.n171 36.1417
R27273 avss.n342 avss.n174 36.1417
R27274 avss.n349 avss.n174 36.1417
R27275 avss.n330 avss.n177 36.1417
R27276 avss.n337 avss.n177 36.1417
R27277 avss.n318 avss.n180 36.1417
R27278 avss.n325 avss.n180 36.1417
R27279 avss.n306 avss.n183 36.1417
R27280 avss.n313 avss.n183 36.1417
R27281 avss.n294 avss.n186 36.1417
R27282 avss.n301 avss.n186 36.1417
R27283 avss.n282 avss.n189 36.1417
R27284 avss.n289 avss.n189 36.1417
R27285 avss.n270 avss.n192 36.1417
R27286 avss.n277 avss.n192 36.1417
R27287 avss.n258 avss.n195 36.1417
R27288 avss.n265 avss.n195 36.1417
R27289 avss.n246 avss.n198 36.1417
R27290 avss.n253 avss.n198 36.1417
R27291 avss.n234 avss.n201 36.1417
R27292 avss.n241 avss.n201 36.1417
R27293 avss.n222 avss.n204 36.1417
R27294 avss.n229 avss.n204 36.1417
R27295 avss.n654 avss.n649 36.1417
R27296 avss.n654 avss.n645 36.1417
R27297 avss.n661 avss.n645 36.1417
R27298 avss.n661 avss.n641 36.1417
R27299 avss.n668 avss.n641 36.1417
R27300 avss.n668 avss.n636 36.1417
R27301 avss.n676 avss.n636 36.1417
R27302 avss.n676 avss.n637 36.1417
R27303 avss.n637 avss.n632 36.1417
R27304 avss.n688 avss.n632 36.1417
R27305 avss.n688 avss.n629 36.1417
R27306 avss.n695 avss.n629 36.1417
R27307 avss.n695 avss.n625 36.1417
R27308 avss.n709 avss.n625 36.1417
R27309 avss.n709 avss.n708 36.1417
R27310 avss.n708 avss.n623 36.1417
R27311 avss.n623 avss.n621 36.1417
R27312 avss.n720 avss.n621 36.1417
R27313 avss.n720 avss.n619 36.1417
R27314 avss.n729 avss.n619 36.1417
R27315 avss.n729 avss.n616 36.1417
R27316 avss.n736 avss.n616 36.1417
R27317 avss.n736 avss.n612 36.1417
R27318 avss.n743 avss.n612 36.1417
R27319 avss.n743 avss.n609 36.1417
R27320 avss.n750 avss.n609 36.1417
R27321 avss.n750 avss.n606 36.1417
R27322 avss.n757 avss.n606 36.1417
R27323 avss.n757 avss.n603 36.1417
R27324 avss.n764 avss.n603 36.1417
R27325 avss.n764 avss.n600 36.1417
R27326 avss.n773 avss.n600 36.1417
R27327 avss.n773 avss.n597 36.1417
R27328 avss.n779 avss.n597 36.1417
R27329 avss.n779 avss.n594 36.1417
R27330 avss.n786 avss.n594 36.1417
R27331 avss.n786 avss.n581 36.1417
R27332 avss.n854 avss.n581 36.1417
R27333 avss.n130 avss.n123 36.1417
R27334 avss.n124 avss.n123 36.1417
R27335 avss.n210 avss.n207 36.1417
R27336 avss.n217 avss.n207 36.1417
R27337 avss.n153 avss.n117 36.1417
R27338 avss.n1013 avss.n53 35.7393
R27339 avss.t286 avss.t221 35.6315
R27340 avss.n432 avss.n430 35.5561
R27341 avss.n427 avss.n424 35.5561
R27342 avss.n499 avss.n488 35.1094
R27343 avss.n545 avss.n466 35.1094
R27344 avss.t284 avss.t62 34.7831
R27345 avss.n672 avss.t192 34.4853
R27346 avss.n734 avss.t178 34.4853
R27347 avss.n745 avss.t313 34.4853
R27348 avss.n404 avss.n403 34.4123
R27349 avss.n403 avss.n402 34.4123
R27350 avss.n156 avss.n155 34.4123
R27351 avss.n157 avss.n156 34.4123
R27352 avss.n776 avss.t139 33.6338
R27353 avss.n1023 avss.t217 33.2544
R27354 avss.t137 avss.n776 32.7823
R27355 avss.n875 avss.n22 32.5005
R27356 avss.t150 avss.n875 32.5005
R27357 avss.n873 avss.n861 32.5005
R27358 avss.n861 avss.t55 32.5005
R27359 avss.n874 avss.n862 32.5005
R27360 avss.n862 avss.t55 32.5005
R27361 avss.n1100 avss.n1099 32.5005
R27362 avss.n1101 avss.n1100 32.5005
R27363 avss.n1097 avss.n1096 32.5005
R27364 avss.n1096 avss.n1095 32.5005
R27365 avss.n1093 avss.n1092 32.5005
R27366 avss.n1094 avss.n1093 32.5005
R27367 avss.n1083 avss.n1082 32.5005
R27368 avss.n1082 avss.n1081 32.5005
R27369 avss.n1079 avss.n1078 32.5005
R27370 avss.n1080 avss.n1079 32.5005
R27371 avss.t190 avss.n672 31.9308
R27372 avss.n734 avss.t196 31.9308
R27373 avss.n135 avss.t5 31.8139
R27374 avss.n1081 avss.t305 31.4638
R27375 avss.t135 avss.t172 31.3897
R27376 avss.t315 avss.t361 30.5413
R27377 avss.t237 avss.t287 29.693
R27378 avss.n506 avss.n483 29.6559
R27379 avss.n523 avss.n522 29.6559
R27380 avss.n539 avss.n538 29.6559
R27381 avss.n428 avss.n419 29.4328
R27382 avss.n425 avss.n420 29.4328
R27383 avss.n426 avss.n419 29.4328
R27384 avss.n420 avss.n417 29.4328
R27385 avss.t182 avss.n656 29.3764
R27386 avss.t202 avss.n711 29.3764
R27387 avss.n713 avss.t368 29.3764
R27388 avss.n902 avss.n901 28.9887
R27389 avss.n990 avss.n67 28.9887
R27390 avss.t247 avss.t98 28.9058
R27391 avss.t71 avss.t398 28.65
R27392 avss.t242 avss.t87 27.1479
R27393 avss.n874 avss.n864 27.1064
R27394 avss.n873 avss.n863 27.1064
R27395 avss.t27 avss.t81 26.5545
R27396 avss.n1041 avss.t129 26.4633
R27397 avss.n1036 avss.t88 26.4633
R27398 avss.n41 avss.t115 26.4633
R27399 avss.n1031 avss.t76 26.4633
R27400 avss.n1050 avss.t90 26.4633
R27401 avss.n1056 avss.t52 26.4633
R27402 avss.n1066 avss.t80 26.4633
R27403 avss.n1061 avss.t36 26.4633
R27404 avss.n28 avss.t105 26.4633
R27405 avss.n36 avss.t57 26.4633
R27406 avss.t312 avss.t226 26.2995
R27407 avss.t244 avss.t341 26.092
R27408 avss.t171 avss.t302 25.4512
R27409 avss.n870 avss.t74 25.2191
R27410 avss.n867 avss.t54 25.2191
R27411 avss.t186 avss.n671 24.2676
R27412 avss.t168 avss.n673 24.2676
R27413 avss.t35 avss.t319 23.7898
R27414 avss.n16 avss.t339 23.7186
R27415 avss.n1086 avss.t336 23.4728
R27416 avss.n1089 avss.t342 23.4728
R27417 avss.n16 avss.t383 23.4728
R27418 avss.t176 avss.t71 23.2782
R27419 avss.n762 avss.t141 22.5646
R27420 avss.n1080 avss.t217 22.5108
R27421 avss.n901 avss.n900 22.5005
R27422 avss.n900 avss.n899 22.5005
R27423 avss.n575 avss.n574 22.5005
R27424 avss.n899 avss.n575 22.5005
R27425 avss.n67 avss.n65 22.5005
R27426 avss.n78 avss.n65 22.5005
R27427 avss.n999 avss.n66 22.5005
R27428 avss.n78 avss.n66 22.5005
R27429 avss.n1094 avss.t234 22.255
R27430 avss.t343 avss.t176 22.255
R27431 avss.n987 avss.t270 22.0815
R27432 avss.t392 avss.t311 22.0578
R27433 avss.t251 avss.n658 21.7131
R27434 avss.n693 avss.t198 21.7131
R27435 avss.n746 avss.t204 21.7131
R27436 avss.n793 avss.n584 21.3347
R27437 avss.n768 avss.t142 21.2805
R27438 avss.n768 avss.t140 21.2805
R27439 avss.n614 avss.t179 21.2805
R27440 avss.n614 avss.t205 21.2805
R27441 avss.n725 avss.t195 21.2805
R27442 avss.n725 avss.t197 21.2805
R27443 avss.n703 avss.t209 21.2805
R27444 avss.n703 avss.t189 21.2805
R27445 avss.n627 avss.t201 21.2805
R27446 avss.n627 avss.t203 21.2805
R27447 avss.n684 avss.t193 21.2805
R27448 avss.n684 avss.t199 21.2805
R27449 avss.n634 avss.t187 21.2805
R27450 avss.n634 avss.t191 21.2805
R27451 avss.n643 avss.t181 21.2805
R27452 avss.n643 avss.t185 21.2805
R27453 avss.t121 avss.t241 21.2094
R27454 avss.n589 avss.n584 21.1018
R27455 avss.n589 avss.n583 20.9741
R27456 avss.n847 avss.n846 20.8934
R27457 avss.n846 avss.n845 20.8934
R27458 avss.n812 avss.n811 20.8934
R27459 avss.n813 avss.n812 20.8934
R27460 avss.n979 avss.n978 20.8934
R27461 avss.n978 avss.n77 20.8934
R27462 avss.n982 avss.n981 20.8934
R27463 avss.n983 avss.n982 20.8934
R27464 avss.t335 avss.t396 20.7202
R27465 avss.t208 avss.n8 20.4359
R27466 avss.n1040 avss.n1039 20.3733
R27467 avss.n1038 avss.n1037 20.3733
R27468 avss.n1028 avss.n1027 20.3733
R27469 avss.n1030 avss.n1029 20.3733
R27470 avss.n1053 avss.n1052 20.3733
R27471 avss.n1055 avss.n1054 20.3733
R27472 avss.n1065 avss.n1064 20.3733
R27473 avss.n1063 avss.n1062 20.3733
R27474 avss.n33 avss.n32 20.3733
R27475 avss.n35 avss.n34 20.3733
R27476 avss.t378 avss.t149 20.361
R27477 avss avss.n436 20.2672
R27478 avss.n14 avss.n12 20.1729
R27479 avss.n18 avss.n12 20.1729
R27480 avss.n15 avss.n13 20.1729
R27481 avss.n18 avss.n13 20.1729
R27482 avss.n1088 avss.n1087 20.1668
R27483 avss.t282 avss.n986 19.7448
R27484 avss.t296 avss.n984 19.7448
R27485 avss.n647 avss.t352 19.1587
R27486 avss.t204 avss.n745 19.1587
R27487 avss.t141 avss.n761 18.3072
R27488 avss.n402 avss.t320 18.2402
R27489 avss.n1041 avss.t131 18.0193
R27490 avss.t89 avss.n1036 18.0193
R27491 avss.n41 avss.t117 18.0193
R27492 avss.n1031 avss.t77 18.0193
R27493 avss.n1050 avss.t92 18.0193
R27494 avss.n1056 avss.t53 18.0193
R27495 avss.n1066 avss.t83 18.0193
R27496 avss.t38 avss.n1061 18.0193
R27497 avss.n28 avss.t107 18.0193
R27498 avss.n36 avss.t58 18.0193
R27499 avss.n529 avss.n528 17.9618
R27500 avss.n516 avss.n480 17.9618
R27501 avss.n516 avss.n515 17.9618
R27502 avss.n528 avss.n476 17.9618
R27503 avss.n443 avss.n442 17.9561
R27504 avss.t155 avss.t30 17.816
R27505 avss.n588 avss.n585 17.6946
R27506 avss.n443 avss.n414 17.6005
R27507 avss.n870 avss.t75 17.2863
R27508 avss.n867 avss.t56 17.2863
R27509 avss.t360 avss.t114 16.9676
R27510 avss.n496 avss 16.7292
R27511 avss.t340 avss.t247 16.6274
R27512 avss.n674 avss.t186 16.6043
R27513 avss.n674 avss.t168 16.6043
R27514 avss.n731 avss.t194 16.6043
R27515 avss.n797 avss.t13 16.5305
R27516 avss.n797 avss.t19 16.5305
R27517 avss.n795 avss.t21 16.5305
R27518 avss.n795 avss.t11 16.5305
R27519 avss.n801 avss.t25 16.5305
R27520 avss.n801 avss.t17 16.5305
R27521 avss.n799 avss.t23 16.5305
R27522 avss.n799 avss.t148 16.5305
R27523 avss.n559 avss.t344 16.5305
R27524 avss.n559 avss.t65 16.5305
R27525 avss.n557 avss.t289 16.5305
R27526 avss.n557 avss.t127 16.5305
R27527 avss.n563 avss.t347 16.5305
R27528 avss.n563 avss.t345 16.5305
R27529 avss.n836 avss.t295 16.5305
R27530 avss.n836 avss.t291 16.5305
R27531 avss.t69 avss.n820 16.5305
R27532 avss.n820 avss.t346 16.5305
R27533 avss.n833 avss.t133 16.5305
R27534 avss.n833 avss.t293 16.5305
R27535 avss.n86 avss.t281 16.5305
R27536 avss.n86 avss.t277 16.5305
R27537 avss.n84 avss.t273 16.5305
R27538 avss.n84 avss.t269 16.5305
R27539 avss.n90 avss.t271 16.5305
R27540 avss.n90 avss.t283 16.5305
R27541 avss.n88 avss.t275 16.5305
R27542 avss.n88 avss.t297 16.5305
R27543 avss.n109 avss.t349 16.5305
R27544 avss.n109 avss.t101 16.5305
R27545 avss.n107 avss.t389 16.5305
R27546 avss.n107 avss.t46 16.5305
R27547 avss.n96 avss.t351 16.5305
R27548 avss.n96 avss.t348 16.5305
R27549 avss.n94 avss.t391 16.5305
R27550 avss.n94 avss.t388 16.5305
R27551 avss.n970 avss.t112 16.5305
R27552 avss.n970 avss.t350 16.5305
R27553 avss.n967 avss.t96 16.5305
R27554 avss.n967 avss.t390 16.5305
R27555 avss.t366 avss.t327 16.1193
R27556 avss.n771 avss.n770 16.0275
R27557 avss.n794 avss.n583 15.8429
R27558 avss.t258 avss.t194 15.3271
R27559 avss.n437 avss 15.2894
R27560 avss.n769 avss.n767 15.2801
R27561 avss.n1077 avss.n17 14.9605
R27562 avss.n1091 avss.n1090 14.9605
R27563 avss.n1085 avss.n1084 14.9605
R27564 avss.n1075 avss.n1074 14.9605
R27565 avss.t325 avss.t218 14.8368
R27566 avss.t396 avss.t248 14.581
R27567 avss.n913 avss.t63 14.0925
R27568 avss.n554 avss.t126 14.0925
R27569 avss.n821 avss.t67 14.0925
R27570 avss.n832 avss.t132 14.0925
R27571 avss.n969 avss.t111 14.0925
R27572 avss.n966 avss.t95 14.0925
R27573 avss.n941 avss.t99 14.0925
R27574 avss.n104 avss.t44 14.0925
R27575 avss.n46 avss.t338 14.0694
R27576 avss.n659 avss.t180 14.0498
R27577 avss.t358 avss.n691 14.0498
R27578 avss.n713 avss.t208 14.0498
R27579 avss.t398 avss.n1020 13.0463
R27580 avss.n491 avss 12.9272
R27581 avss.n412 avss.t167 12.8791
R27582 avss.n1095 avss.t165 12.7905
R27583 avss.n21 avss.n19 12.7179
R27584 avss.t151 avss.n19 12.7179
R27585 avss.n1076 avss.n20 12.7179
R27586 avss.t151 avss.n20 12.7179
R27587 avss.t331 avss.n77 12.513
R27588 avss.n1102 avss.t157 12.2789
R27589 avss.n59 avss.n56 12.189
R27590 avss.n433 avss.n432 12.0894
R27591 avss.n430 avss.n429 12.0894
R27592 avss.n438 avss.n414 12.0894
R27593 avss.n442 avss.n415 12.0894
R27594 avss.n881 avss.t314 11.9874
R27595 avss.t266 avss.t267 11.8775
R27596 avss.n1110 avss.n1109 11.8447
R27597 avss.n63 avss.t81 11.7601
R27598 avss.n657 avss.t182 11.4954
R27599 avss.n712 avss.t202 11.4954
R27600 avss.t368 avss.n712 11.4954
R27601 avss.n78 avss.t331 11.409
R27602 avss.t123 avss.t367 11.0291
R27603 avss.n69 avss.n49 10.9999
R27604 avss.n987 avss.n77 10.673
R27605 avss.n93 avss.n82 10.3632
R27606 avss.n977 avss.n976 10.3105
R27607 avss.n849 avss.n848 10.3105
R27608 avss.n810 avss.n809 10.3105
R27609 avss.n550 avss.n549 10.2952
R27610 avss.n1044 avss.n1026 9.42076
R27611 avss.n1034 avss.n1026 9.42076
R27612 avss.n650 avss.n649 9.36464
R27613 avss.n408 avss.n116 9.35869
R27614 avss.n409 avss.n115 9.35222
R27615 avss.n410 avss.n114 9.34791
R27616 avss.n407 avss.n406 9.33929
R27617 avss.n405 avss.n55 9.33929
R27618 avss.n129 avss.n128 9.30641
R27619 avss.n652 avss.n651 9.3005
R27620 avss.n651 avss.n650 9.3005
R27621 avss.n664 avss.n663 9.3005
R27622 avss.n680 avss.n679 9.3005
R27623 avss.n679 avss.n678 9.3005
R27624 avss.n679 avss.n635 9.3005
R27625 avss.n685 avss.n628 9.3005
R27626 avss.n686 avss.n685 9.3005
R27627 avss.n685 avss.n682 9.3005
R27628 avss.n701 avss.n700 9.3005
R27629 avss.n700 avss.n699 9.3005
R27630 avss.n700 avss.n698 9.3005
R27631 avss.n705 avss.n704 9.3005
R27632 avss.n726 avss.n615 9.3005
R27633 avss.n727 avss.n726 9.3005
R27634 avss.n726 avss.n723 9.3005
R27635 avss.n741 avss.n740 9.3005
R27636 avss.n740 avss.n613 9.3005
R27637 avss.n740 avss.n739 9.3005
R27638 avss.n770 avss.n601 9.3005
R27639 avss.n783 avss.n782 9.3005
R27640 avss.n782 avss.n781 9.3005
R27641 avss.n852 avss.n851 9.3005
R27642 avss.n851 avss.n582 9.3005
R27643 avss.n754 avss.n753 9.3005
R27644 avss.n753 avss.n752 9.3005
R27645 avss.n654 avss.n653 9.3005
R27646 avss.n645 avss.n644 9.3005
R27647 avss.n662 avss.n661 9.3005
R27648 avss.n642 avss.n641 9.3005
R27649 avss.n668 avss.n667 9.3005
R27650 avss.n666 avss.n636 9.3005
R27651 avss.n677 avss.n676 9.3005
R27652 avss.n637 avss.n633 9.3005
R27653 avss.n681 avss.n632 9.3005
R27654 avss.n688 avss.n687 9.3005
R27655 avss.n683 avss.n629 9.3005
R27656 avss.n696 avss.n695 9.3005
R27657 avss.n697 avss.n625 9.3005
R27658 avss.n709 avss.n626 9.3005
R27659 avss.n708 avss.n707 9.3005
R27660 avss.n706 avss.n623 9.3005
R27661 avss.n702 avss.n621 9.3005
R27662 avss.n721 avss.n720 9.3005
R27663 avss.n722 avss.n619 9.3005
R27664 avss.n729 avss.n728 9.3005
R27665 avss.n724 avss.n616 9.3005
R27666 avss.n737 avss.n736 9.3005
R27667 avss.n738 avss.n612 9.3005
R27668 avss.n743 avss.n742 9.3005
R27669 avss.n609 avss.n608 9.3005
R27670 avss.n751 avss.n750 9.3005
R27671 avss.n607 avss.n606 9.3005
R27672 avss.n757 avss.n756 9.3005
R27673 avss.n603 avss.n602 9.3005
R27674 avss.n765 avss.n764 9.3005
R27675 avss.n766 avss.n600 9.3005
R27676 avss.n773 avss.n772 9.3005
R27677 avss.n597 avss.n596 9.3005
R27678 avss.n780 avss.n779 9.3005
R27679 avss.n595 avss.n594 9.3005
R27680 avss.n786 avss.n785 9.3005
R27681 avss.n784 avss.n581 9.3005
R27682 avss.n854 avss.n853 9.3005
R27683 avss.n891 avss.n864 9.3005
R27684 avss.n865 avss.n863 9.3005
R27685 avss.n879 avss.n878 9.3005
R27686 avss.n1008 avss.n58 9.3005
R27687 avss.n128 avss.n127 9.3005
R27688 avss.n130 avss.n129 9.3005
R27689 avss.n126 avss.n123 9.3005
R27690 avss.n125 avss.n124 9.3005
R27691 avss.n215 avss.n214 9.3005
R27692 avss.n214 avss.n213 9.3005
R27693 avss.n227 avss.n226 9.3005
R27694 avss.n226 avss.n225 9.3005
R27695 avss.n239 avss.n238 9.3005
R27696 avss.n238 avss.n237 9.3005
R27697 avss.n251 avss.n250 9.3005
R27698 avss.n250 avss.n249 9.3005
R27699 avss.n263 avss.n262 9.3005
R27700 avss.n262 avss.n261 9.3005
R27701 avss.n275 avss.n274 9.3005
R27702 avss.n274 avss.n273 9.3005
R27703 avss.n287 avss.n286 9.3005
R27704 avss.n286 avss.n285 9.3005
R27705 avss.n299 avss.n298 9.3005
R27706 avss.n298 avss.n297 9.3005
R27707 avss.n311 avss.n310 9.3005
R27708 avss.n310 avss.n309 9.3005
R27709 avss.n323 avss.n322 9.3005
R27710 avss.n322 avss.n321 9.3005
R27711 avss.n335 avss.n334 9.3005
R27712 avss.n334 avss.n333 9.3005
R27713 avss.n347 avss.n346 9.3005
R27714 avss.n346 avss.n345 9.3005
R27715 avss.n359 avss.n358 9.3005
R27716 avss.n358 avss.n357 9.3005
R27717 avss.n371 avss.n370 9.3005
R27718 avss.n370 avss.n369 9.3005
R27719 avss.n383 avss.n382 9.3005
R27720 avss.n382 avss.n381 9.3005
R27721 avss.n393 avss.n0 9.3005
R27722 avss.n394 avss.n393 9.3005
R27723 avss.n223 avss.n222 9.3005
R27724 avss.n224 avss.n204 9.3005
R27725 avss.n229 avss.n228 9.3005
R27726 avss.n235 avss.n234 9.3005
R27727 avss.n236 avss.n201 9.3005
R27728 avss.n241 avss.n240 9.3005
R27729 avss.n247 avss.n246 9.3005
R27730 avss.n248 avss.n198 9.3005
R27731 avss.n253 avss.n252 9.3005
R27732 avss.n259 avss.n258 9.3005
R27733 avss.n260 avss.n195 9.3005
R27734 avss.n265 avss.n264 9.3005
R27735 avss.n271 avss.n270 9.3005
R27736 avss.n272 avss.n192 9.3005
R27737 avss.n277 avss.n276 9.3005
R27738 avss.n283 avss.n282 9.3005
R27739 avss.n284 avss.n189 9.3005
R27740 avss.n289 avss.n288 9.3005
R27741 avss.n295 avss.n294 9.3005
R27742 avss.n296 avss.n186 9.3005
R27743 avss.n301 avss.n300 9.3005
R27744 avss.n307 avss.n306 9.3005
R27745 avss.n308 avss.n183 9.3005
R27746 avss.n313 avss.n312 9.3005
R27747 avss.n319 avss.n318 9.3005
R27748 avss.n320 avss.n180 9.3005
R27749 avss.n325 avss.n324 9.3005
R27750 avss.n331 avss.n330 9.3005
R27751 avss.n332 avss.n177 9.3005
R27752 avss.n337 avss.n336 9.3005
R27753 avss.n343 avss.n342 9.3005
R27754 avss.n344 avss.n174 9.3005
R27755 avss.n349 avss.n348 9.3005
R27756 avss.n355 avss.n354 9.3005
R27757 avss.n356 avss.n171 9.3005
R27758 avss.n361 avss.n360 9.3005
R27759 avss.n367 avss.n366 9.3005
R27760 avss.n368 avss.n168 9.3005
R27761 avss.n373 avss.n372 9.3005
R27762 avss.n379 avss.n378 9.3005
R27763 avss.n380 avss.n165 9.3005
R27764 avss.n385 avss.n384 9.3005
R27765 avss.n391 avss.n390 9.3005
R27766 avss.n392 avss.n162 9.3005
R27767 avss.n396 avss.n395 9.3005
R27768 avss.n211 avss.n210 9.3005
R27769 avss.n212 avss.n207 9.3005
R27770 avss.n217 avss.n216 9.3005
R27771 avss.n154 avss.n152 9.3005
R27772 avss.n1011 avss.n1010 9.20927
R27773 avss.n673 avss.t190 8.94099
R27774 avss.n717 avss.t258 8.94099
R27775 avss.t196 avss.n732 8.94099
R27776 avss.t276 avss.n78 8.83289
R27777 avss.t274 avss.n985 8.83289
R27778 avss.n882 avss.n880 8.81442
R27779 avss.n829 avss.t414 8.80038
R27780 avss.n828 avss.t433 8.80038
R27781 avss.n827 avss.t415 8.80038
R27782 avss.n826 avss.t424 8.80038
R27783 avss.n825 avss.t416 8.80038
R27784 avss.n824 avss.t437 8.80038
R27785 avss.n823 avss.t419 8.80038
R27786 avss.n553 avss.t438 8.80038
R27787 avss.n963 avss.t426 8.80038
R27788 avss.n962 avss.t410 8.80038
R27789 avss.n961 avss.t441 8.80038
R27790 avss.n960 avss.t427 8.80038
R27791 avss.n959 avss.t411 8.80038
R27792 avss.n958 avss.t428 8.80038
R27793 avss.n957 avss.t412 8.80038
R27794 avss.n956 avss.t442 8.80038
R27795 avss.n919 avss.t418 8.73382
R27796 avss.n920 avss.t436 8.73382
R27797 avss.n921 avss.t421 8.73382
R27798 avss.n922 avss.t425 8.73382
R27799 avss.n923 avss.t422 8.73382
R27800 avss.n924 avss.t439 8.73382
R27801 avss.n925 avss.t423 8.73382
R27802 avss.n926 avss.t440 8.73382
R27803 avss.n947 avss.t430 8.73382
R27804 avss.n948 avss.t413 8.73382
R27805 avss.n949 avss.t443 8.73382
R27806 avss.n950 avss.t434 8.73382
R27807 avss.n951 avss.t417 8.73382
R27808 avss.n952 avss.t435 8.73382
R27809 avss.n953 avss.t420 8.73382
R27810 avss.n954 avss.t444 8.73382
R27811 avss.n504 avss.n487 8.61832
R27812 avss.n505 avss.n504 8.61832
R27813 avss.n506 avss.n505 8.61832
R27814 avss.n512 avss.n483 8.61832
R27815 avss.n513 avss.n512 8.61832
R27816 avss.n514 avss.n513 8.61832
R27817 avss.n521 avss.n479 8.61832
R27818 avss.n522 avss.n521 8.61832
R27819 avss.n523 avss.n477 8.61832
R27820 avss.n530 avss.n477 8.61832
R27821 avss.n472 avss.n464 8.61832
R27822 avss.n540 avss.n472 8.61832
R27823 avss.n540 avss.n539 8.61832
R27824 avss.n538 avss.n473 8.61832
R27825 avss.n532 avss.n473 8.61832
R27826 avss.n532 avss.n531 8.61832
R27827 avss.n498 avss.n497 8.61832
R27828 avss.n497 avss.n496 8.61832
R27829 avss.n491 avss.n463 8.61832
R27830 avss.t173 avss.t310 8.48406
R27831 avss.n880 avss.n59 8.4666
R27832 avss.n891 avss.n890 8.37766
R27833 avss.n890 avss.n865 8.37766
R27834 avss.n38 avss.n30 8.11041
R27835 avss.n1070 avss.n30 8.11041
R27836 avss.n777 avss.t137 8.08952
R27837 avss.n1008 avss.n1007 8.02619
R27838 avss.n1007 avss.n59 8.00675
R27839 avss.n892 avss.n865 7.938
R27840 avss.n892 avss.n891 7.938
R27841 avss avss.n850 7.87749
R27842 avss.t0 avss.t373 7.63571
R27843 avss.n927 avss.n553 7.62598
R27844 avss.n956 avss.n955 7.62598
R27845 avss.n883 avss.n879 7.48375
R27846 avss.n436 avss.n433 7.46717
R27847 avss.n438 avss.n437 7.46717
R27848 avss.n429 avss.n427 7.46717
R27849 avss.n424 avss.n415 7.46717
R27850 avss.t139 avss.n775 7.23804
R27851 avss.n883 avss.n882 7.16066
R27852 avss.n934 avss.n933 7.079
R27853 avss.t338 avss.t364 6.90708
R27854 avss.n879 avss.n57 6.89147
R27855 avss.n1008 avss.n57 6.89083
R27856 avss.n48 avss.n45 6.88285
R27857 avss.n63 avss.n48 6.88285
R27858 avss.n47 avss.n44 6.88285
R27859 avss.n47 avss.n46 6.88285
R27860 avss.t1 avss.t85 6.78735
R27861 avss.n413 avss 6.6041
R27862 avss.n412 avss.n411 6.54285
R27863 avss.n894 avss.n893 6.5005
R27864 avss.n895 avss.n894 6.5005
R27865 avss.n889 avss.n888 6.5005
R27866 avss.n888 avss.n887 6.5005
R27867 avss.n905 avss.n565 6.47706
R27868 avss.n905 avss.n561 6.47706
R27869 avss.n838 avss.n835 6.47706
R27870 avss.n838 avss.n556 6.47706
R27871 avss.n972 avss.n76 6.47706
R27872 avss.n111 avss.n76 6.47706
R27873 avss.n102 avss.n75 6.47706
R27874 avss.n106 avss.n75 6.47706
R27875 avss.n547 avss.n463 6.46387
R27876 avss.n690 avss.t192 6.38657
R27877 avss.n716 avss.n8 6.38657
R27878 avss.t178 avss.n733 6.38657
R27879 avss.n733 avss.t313 6.38657
R27880 avss.n1112 avss.n1111 6.05765
R27881 avss.n1022 avss.n1021 5.90959
R27882 avss.n1023 avss.n1022 5.90959
R27883 avss.n1025 avss.n1024 5.90959
R27884 avss.n1024 avss.n1023 5.90959
R27885 avss.n69 avss.t40 5.88388
R27886 avss.n1111 avss.n2 5.78505
R27887 avss.n881 avss.n872 5.7846
R27888 avss.n871 avss.n870 5.76099
R27889 avss.n868 avss.n867 5.76099
R27890 avss.n850 avss.n794 5.71512
R27891 avss.n1035 avss.n1034 5.70305
R27892 avss.n1033 avss.n1032 5.70305
R27893 avss.n1058 avss.n1057 5.70305
R27894 avss.n1060 avss.n1059 5.70305
R27895 avss.n38 avss.n37 5.70305
R27896 avss.n866 avss.n865 5.6605
R27897 avss.n1042 avss.n1041 5.6605
R27898 avss.n1036 avss.n1035 5.6605
R27899 avss.n1044 avss.n1043 5.6605
R27900 avss.n42 avss.n41 5.6605
R27901 avss.n1032 avss.n1031 5.6605
R27902 avss.n1046 avss.n1045 5.6605
R27903 avss.n1051 avss.n1050 5.6605
R27904 avss.n1057 avss.n1056 5.6605
R27905 avss.n1049 avss.n31 5.6605
R27906 avss.n1067 avss.n1066 5.6605
R27907 avss.n1061 avss.n1060 5.6605
R27908 avss.n1069 avss.n1068 5.6605
R27909 avss.n29 avss.n28 5.6605
R27910 avss.n37 avss.n36 5.6605
R27911 avss.n1071 avss.n1070 5.6605
R27912 avss.n891 avss.n872 5.6605
R27913 avss.t163 avss.t323 5.62808
R27914 avss.n794 avss.n793 5.46789
R27915 avss.n551 avss.n112 5.276
R27916 avss.n790 avss.n586 5.27077
R27917 avss.n790 avss.n789 5.27077
R27918 avss.n587 avss.n585 5.27077
R27919 avss.n789 avss.n587 5.27077
R27920 avss.n1006 avss.n1005 5.27077
R27921 avss.n1005 avss.n1004 5.27077
R27922 avss.n885 avss.n884 5.27077
R27923 avss.n886 avss.n885 5.27077
R27924 avss.t180 avss.t251 5.10935
R27925 avss.t198 avss.t358 5.10935
R27926 avss.n558 avss.n556 5.07277
R27927 avss.n838 avss.n837 5.07277
R27928 avss.n835 avss.n834 5.07277
R27929 avss.n108 avss.n106 5.07277
R27930 avss.n95 avss.n75 5.07277
R27931 avss.n968 avss.n102 5.07277
R27932 avss.n792 avss.n791 5.0436
R27933 avss.n791 avss.n577 5.0436
R27934 avss.n591 avss.n590 5.0436
R27935 avss.n591 avss.n578 5.0436
R27936 avss.n62 avss.n60 5.0436
R27937 avss.t27 avss.n62 5.0436
R27938 avss.n877 avss.n61 5.0436
R27939 avss.t27 avss.n61 5.0436
R27940 avss.n1019 avss.n1018 5.0436
R27941 avss.n1020 avss.n1019 5.0436
R27942 avss.n133 avss.n54 5.0436
R27943 avss.n134 avss.n133 5.0436
R27944 avss.n459 avss.n458 5.0005
R27945 avss.n458 avss.n457 5.0005
R27946 avss.n450 avss.n446 5.0005
R27947 avss.n456 avss.n450 5.0005
R27948 avss.n454 avss.n453 5.0005
R27949 avss.n455 avss.n454 5.0005
R27950 avss.n452 avss.n449 5.0005
R27951 avss.n451 avss.n449 5.0005
R27952 avss.n561 avss.n560 4.95167
R27953 avss.n817 avss.n565 4.95167
R27954 avss.n111 avss.n110 4.95167
R27955 avss.n972 avss.n971 4.95167
R27956 avss.n550 avss.n413 4.93439
R27957 avss.n1013 avss.n1012 4.86769
R27958 avss.n153 avss.n118 4.6805
R27959 avss.t60 avss.n118 4.6805
R27960 avss.n120 avss.n119 4.6805
R27961 avss.t60 avss.n120 4.6805
R27962 avss.n665 avss.n664 4.63624
R27963 avss.n704 avss.n620 4.63624
R27964 avss.n955 avss.n954 4.60905
R27965 avss.n927 avss.n926 4.60905
R27966 avss.n555 avss.n554 4.5005
R27967 avss.n914 avss.n913 4.5005
R27968 avss.n906 avss.n905 4.5005
R27969 avss.n916 avss.n915 4.5005
R27970 avss.n918 avss.n917 4.5005
R27971 avss.n832 avss.n831 4.5005
R27972 avss.n822 avss.n821 4.5005
R27973 avss.n830 avss.n816 4.5005
R27974 avss.n819 avss.n818 4.5005
R27975 avss.n98 avss.n76 4.5005
R27976 avss.n105 avss.n104 4.5005
R27977 avss.n942 avss.n941 4.5005
R27978 avss.n946 avss.n945 4.5005
R27979 avss.n944 avss.n943 4.5005
R27980 avss.n966 avss.n965 4.5005
R27981 avss.n969 avss.n100 4.5005
R27982 avss.n964 avss.n101 4.5005
R27983 avss.n974 avss.n973 4.5005
R27984 avss.n447 avss.n444 4.3603
R27985 avss.n461 avss.n445 4.34678
R27986 avss.n447 avss.n445 4.34003
R27987 avss.n866 avss.n26 4.00655
R27988 avss.n841 avss.n839 3.9532
R27989 avss.n841 avss.n840 3.9532
R27990 avss.n904 avss.n567 3.9532
R27991 avss.n840 avss.n567 3.9532
R27992 avss.n989 avss.n988 3.9532
R27993 avss.n988 avss.n987 3.9532
R27994 avss.n995 avss.n994 3.9532
R27995 avss.n996 avss.n995 3.9532
R27996 avss.n1111 avss.n1110 3.94537
R27997 avss.n929 avss.n928 3.9105
R27998 avss.n1020 avss.t337 3.83749
R27999 avss.n692 avss.t200 3.83214
R28000 avss.n748 avss.t206 3.83214
R28001 avss.n747 avss.t359 3.83214
R28002 avss.n462 avss.n461 3.78259
R28003 avss.n819 avss.n562 3.77378
R28004 avss.n975 avss.n974 3.77378
R28005 avss.n907 avss.n906 3.77209
R28006 avss.n99 avss.n98 3.77209
R28007 avss.n915 avss.n912 3.77014
R28008 avss.n943 avss.n940 3.77014
R28009 avss.n1074 avss.n1073 3.68964
R28010 avss.n1043 avss.n40 3.57087
R28011 avss.n1047 avss.n1046 3.57087
R28012 avss.n1049 avss.n1048 3.57087
R28013 avss.n1068 avss.n27 3.57087
R28014 avss.n1072 avss.n1071 3.57087
R28015 avss.n93 avss.n92 3.4105
R28016 avss.n939 avss.n938 3.4105
R28017 avss.n911 avss.n910 3.4105
R28018 avss.n804 avss.n803 3.4105
R28019 avss.n1039 avss.t405 3.3065
R28020 avss.n1039 avss.t130 3.3065
R28021 avss.n1037 avss.t89 3.3065
R28022 avss.n1037 avss.t403 3.3065
R28023 avss.n1027 avss.t407 3.3065
R28024 avss.n1027 avss.t116 3.3065
R28025 avss.t77 avss.n1030 3.3065
R28026 avss.n1030 avss.t404 3.3065
R28027 avss.n1052 avss.t399 3.3065
R28028 avss.n1052 avss.t91 3.3065
R28029 avss.t53 avss.n1055 3.3065
R28030 avss.n1055 avss.t397 3.3065
R28031 avss.n1064 avss.t402 3.3065
R28032 avss.n1064 avss.t82 3.3065
R28033 avss.n1062 avss.t38 3.3065
R28034 avss.n1062 avss.t400 3.3065
R28035 avss.n32 avss.t401 3.3065
R28036 avss.n32 avss.t106 3.3065
R28037 avss.t58 avss.n35 3.3065
R28038 avss.n35 avss.t406 3.3065
R28039 avss.n1087 avss.t324 3.3065
R28040 avss.n1087 avss.t326 3.3065
R28041 avss.t150 avss.n876 3.2875
R28042 avss.n818 avss.n565 3.23878
R28043 avss.n916 avss.n561 3.23878
R28044 avss.n835 avss.n816 3.23878
R28045 avss.n917 avss.n556 3.23878
R28046 avss.n973 avss.n972 3.23878
R28047 avss.n944 avss.n111 3.23878
R28048 avss.n102 avss.n101 3.23878
R28049 avss.n945 avss.n106 3.23878
R28050 avss.n919 avss.n918 3.21858
R28051 avss.n947 avss.n946 3.21858
R28052 avss.n830 avss.n829 3.12292
R28053 avss.n964 avss.n963 3.12292
R28054 avss.n548 avss.n547 3.1005
R28055 avss.n760 avss.t143 2.98066
R28056 avss.n158 avss.t250 2.96975
R28057 avss.n1014 avss.n1013 2.83532
R28058 avss.n1109 avss.n3 2.6005
R28059 avss.n789 avss.n579 2.55493
R28060 avss.t6 avss.t170 2.54557
R28061 avss.n551 avss.n550 2.47021
R28062 avss.n1070 avss.n1069 2.42291
R28063 avss.n1069 avss.n31 2.42291
R28064 avss.n1045 avss.n1044 2.42291
R28065 avss.n1034 avss.n1033 2.42291
R28066 avss.n1059 avss.n1058 2.42291
R28067 avss.n1059 avss.n38 2.42291
R28068 avss.n514 avss.n479 2.40842
R28069 avss.n531 avss.n530 2.40842
R28070 avss.n549 avss.n443 2.32925
R28071 avss.n1009 avss.n1008 2.31886
R28072 avss.n879 avss.n26 2.31886
R28073 avss.n498 avss.n487 2.28169
R28074 avss.n546 avss.n464 2.28169
R28075 avss.n452 avss.n448 2.25932
R28076 avss.n882 avss.n881 2.2505
R28077 avss.n929 avss.n56 2.221
R28078 avss.n548 avss.n462 2.17339
R28079 avss.n547 avss.n546 2.15496
R28080 avss avss.n932 2.13136
R28081 avss.n928 avss.n927 2.12151
R28082 avss.n818 avss.n816 2.11769
R28083 avss.n917 avss.n916 2.11769
R28084 avss.n973 avss.n101 2.11769
R28085 avss.n945 avss.n944 2.11769
R28086 avss.n552 avss.n551 2.10921
R28087 avss.n1010 avss.n56 2.058
R28088 avss.n935 avss.n103 1.90581
R28089 avss.n928 avss.n552 1.90581
R28090 avss.n911 avss.n552 1.80585
R28091 avss.n1045 avss.n43 1.80222
R28092 avss.n1033 avss.n39 1.80222
R28093 avss.t260 avss.t160 1.69721
R28094 avss.n409 avss.n408 1.6605
R28095 avss.n934 avss.n929 1.65831
R28096 avss.n975 avss.n99 1.58008
R28097 avss.n940 avss.n99 1.58008
R28098 avss.n912 avss.n907 1.58008
R28099 avss.n907 avss.n562 1.58008
R28100 avss.n413 avss.n412 1.55609
R28101 avss.n1017 avss.n51 1.50436
R28102 avss.n135 avss.n51 1.50436
R28103 avss.n52 avss.n50 1.50436
R28104 avss.n135 avss.n50 1.50436
R28105 avss.n211 avss.n113 1.48467
R28106 avss.n933 avss 1.41066
R28107 avss.n136 avss.n1 1.34141
R28108 avss.n410 avss.n409 1.338
R28109 avss.n152 avss.n151 1.32209
R28110 avss.n955 avss.n103 1.31665
R28111 avss.n1023 avss.t384 1.2795
R28112 avss.n670 avss.t184 1.27771
R28113 avss.n718 avss.t188 1.27771
R28114 avss.n761 avss.t370 1.27771
R28115 avss.t233 avss.n592 1.27771
R28116 avss.n407 avss.n55 1.27675
R28117 avss.t224 avss.n401 1.27303
R28118 avss.n876 avss.n64 1.27293
R28119 avss.n141 avss.n140 1.14936
R28120 avss.n149 avss.n148 1.14936
R28121 avss.n142 avss.n141 1.14839
R28122 avss.n150 avss.n149 1.14811
R28123 avss.n137 avss.n136 1.08686
R28124 avss.n138 avss.n137 1.08686
R28125 avss.n139 avss.n138 1.08686
R28126 avss.n140 avss.n139 1.08686
R28127 avss.n145 avss.n144 1.08686
R28128 avss.n147 avss.n146 1.08686
R28129 avss.n148 avss.n147 1.08686
R28130 avss.n151 avss.n150 1.08686
R28131 avss.n146 avss.n145 1.08005
R28132 avss.n1040 avss.n1038 1.05355
R28133 avss.n1029 avss.n1028 1.05355
R28134 avss.n1054 avss.n1053 1.05355
R28135 avss.n1065 avss.n1063 1.05355
R28136 avss.n34 avss.n33 1.05355
R28137 avss.n408 avss.n407 1.00987
R28138 avss.n112 avss.n103 1.00659
R28139 avss.n143 avss.n142 1.00505
R28140 avss.n939 avss.n935 1.00226
R28141 avss.n871 avss.n869 0.955426
R28142 avss.n869 avss.n868 0.953203
R28143 avss.n1011 avss.n1 0.902375
R28144 avss avss.n1112 0.899013
R28145 avss.n411 avss.n113 0.839875
R28146 avss.n829 avss.n828 0.807835
R28147 avss.n828 avss.n827 0.807835
R28148 avss.n827 avss.n826 0.807835
R28149 avss.n826 avss.n825 0.807835
R28150 avss.n825 avss.n824 0.807835
R28151 avss.n824 avss.n823 0.807835
R28152 avss.n823 avss.n553 0.807835
R28153 avss.n963 avss.n962 0.807835
R28154 avss.n962 avss.n961 0.807835
R28155 avss.n961 avss.n960 0.807835
R28156 avss.n960 avss.n959 0.807835
R28157 avss.n959 avss.n958 0.807835
R28158 avss.n958 avss.n957 0.807835
R28159 avss.n957 avss.n956 0.807835
R28160 avss.n920 avss.n919 0.80776
R28161 avss.n921 avss.n920 0.80776
R28162 avss.n922 avss.n921 0.80776
R28163 avss.n923 avss.n922 0.80776
R28164 avss.n924 avss.n923 0.80776
R28165 avss.n925 avss.n924 0.80776
R28166 avss.n926 avss.n925 0.80776
R28167 avss.n948 avss.n947 0.80776
R28168 avss.n949 avss.n948 0.80776
R28169 avss.n950 avss.n949 0.80776
R28170 avss.n951 avss.n950 0.80776
R28171 avss.n952 avss.n951 0.80776
R28172 avss.n953 avss.n952 0.80776
R28173 avss.n954 avss.n953 0.80776
R28174 avss.n460 avss.n446 0.753441
R28175 avss.n770 avss.n769 0.747945
R28176 avss.n802 avss.n800 0.695812
R28177 avss.n914 avss.n555 0.695812
R28178 avss.n560 avss.n558 0.695812
R28179 avss.n834 avss.n817 0.695812
R28180 avss.n831 avss.n822 0.695812
R28181 avss.n937 avss.n936 0.695812
R28182 avss.n91 avss.n89 0.695812
R28183 avss.n110 avss.n108 0.695812
R28184 avss.n97 avss.n95 0.695812
R28185 avss.n971 avss.n968 0.695812
R28186 avss.n942 avss.n105 0.695812
R28187 avss.n965 avss.n100 0.695812
R28188 avss.n909 avss.n908 0.695812
R28189 avss.t280 avss.n79 0.69443
R28190 avss.n931 avss.n930 0.693859
R28191 avss.n798 avss.n796 0.679185
R28192 avss.n87 avss.n85 0.679185
R28193 avss.n837 avss.n564 0.676856
R28194 avss.n803 avss.n802 0.654797
R28195 avss.n92 avss.n91 0.654797
R28196 avss.n1074 avss.n25 0.635318
R28197 avss.n935 avss.n934 0.622375
R28198 avss.n43 avss.n31 0.62119
R28199 avss.n1058 avss.n39 0.62119
R28200 avss.n918 avss.n555 0.572766
R28201 avss.n831 avss.n830 0.572766
R28202 avss.n946 avss.n105 0.572766
R28203 avss.n965 avss.n964 0.572766
R28204 avss.n462 avss.n444 0.571446
R28205 avss.n1038 avss.n1035 0.527027
R28206 avss.n1042 avss.n1040 0.527027
R28207 avss.n1032 avss.n1029 0.527027
R28208 avss.n1028 avss.n42 0.527027
R28209 avss.n1057 avss.n1054 0.527027
R28210 avss.n1053 avss.n1051 0.527027
R28211 avss.n1063 avss.n1060 0.527027
R28212 avss.n1067 avss.n1065 0.527027
R28213 avss.n37 avss.n34 0.527027
R28214 avss.n33 avss.n29 0.527027
R28215 avss.t37 avss.n1094 0.512098
R28216 avss.n1073 avss.n26 0.505881
R28217 avss.n1073 avss.n1072 0.497189
R28218 avss.n1072 avss.n27 0.478977
R28219 avss.n1048 avss.n27 0.478977
R28220 avss.n1048 avss.n1047 0.478977
R28221 avss.n1047 avss.n40 0.478977
R28222 avss.n915 avss.n914 0.451672
R28223 avss.n906 avss.n564 0.451672
R28224 avss.n822 avss.n819 0.451672
R28225 avss.n98 avss.n97 0.451672
R28226 avss.n943 avss.n942 0.451672
R28227 avss.n974 avss.n100 0.451672
R28228 avss.n789 avss.t230 0.426238
R28229 avss.n933 avss.n931 0.416516
R28230 avss.n1010 avss.n1009 0.387296
R28231 avss.n1009 avss.n40 0.380881
R28232 avss.n1112 avss.n1 0.364875
R28233 avss.n986 avss.t100 0.344476
R28234 avss.n938 avss.n937 0.311047
R28235 avss.n910 avss.n909 0.311047
R28236 avss.n1089 avss.n1088 0.291392
R28237 avss.n1088 avss.n1086 0.291392
R28238 avss.n448 avss.n447 0.274029
R28239 avss.n459 avss.n445 0.266214
R28240 avss.n461 avss.n460 0.266214
R28241 avss.n453 avss.n444 0.266214
R28242 avss.n223 avss 0.248811
R28243 avss.n235 avss 0.248811
R28244 avss.n247 avss 0.248811
R28245 avss.n259 avss 0.248811
R28246 avss.n271 avss 0.248811
R28247 avss.n283 avss 0.248811
R28248 avss.n295 avss 0.248811
R28249 avss.n307 avss 0.248811
R28250 avss.n319 avss 0.248811
R28251 avss.n331 avss 0.248811
R28252 avss.n343 avss 0.248811
R28253 avss.n355 avss 0.248811
R28254 avss.n367 avss 0.248811
R28255 avss.n379 avss 0.248811
R28256 avss.n391 avss 0.248811
R28257 avss.n940 avss.n939 0.237405
R28258 avss.n912 avss.n911 0.237405
R28259 avss.n23 avss.n17 0.182466
R28260 avss.n984 avss.t45 0.176117
R28261 avss.n411 avss.n410 0.153
R28262 avss.n152 avss.n113 0.128909
R28263 avss.n1090 avss.n16 0.119588
R28264 avss.n976 avss.n975 0.118318
R28265 avss.n809 avss.n562 0.118318
R28266 avss.n45 avss.n43 0.11675
R28267 avss.n44 avss.n39 0.11675
R28268 avss.n24 avss.n23 0.11673
R28269 avss avss.n112 0.116631
R28270 avss.n976 avss.n93 0.114189
R28271 avss.n809 avss.n804 0.114189
R28272 avss.n25 avss.n24 0.113554
R28273 avss.n893 avss.n892 0.109912
R28274 avss.n890 avss.n889 0.109912
R28275 avss.n1012 avss.n1011 0.10175
R28276 avss.n1021 avss.n30 0.0994362
R28277 avss.n1026 avss.n1025 0.0994362
R28278 avss.n588 avss.n583 0.0907913
R28279 avss.n884 avss.n883 0.0890714
R28280 avss.n1007 avss.n1006 0.0890714
R28281 avss.n586 avss.n584 0.0890714
R28282 avss.n877 avss.n57 0.0866111
R28283 avss.n1015 avss.n54 0.0850455
R28284 avss.n1018 avss.n53 0.0850455
R28285 avss.n880 avss.n60 0.0850455
R28286 avss.n590 avss.n589 0.0850455
R28287 avss.n793 avss.n792 0.0850455
R28288 avss.n144 avss.n143 0.0823182
R28289 avss.n126 avss.n125 0.0815811
R28290 avss.n212 avss.n211 0.0815811
R28291 avss.n224 avss.n223 0.0815811
R28292 avss.n236 avss.n235 0.0815811
R28293 avss.n248 avss.n247 0.0815811
R28294 avss.n260 avss.n259 0.0815811
R28295 avss.n272 avss.n271 0.0815811
R28296 avss.n284 avss.n283 0.0815811
R28297 avss.n296 avss.n295 0.0815811
R28298 avss.n308 avss.n307 0.0815811
R28299 avss.n320 avss.n319 0.0815811
R28300 avss.n332 avss.n331 0.0815811
R28301 avss.n344 avss.n343 0.0815811
R28302 avss.n356 avss.n355 0.0815811
R28303 avss.n368 avss.n367 0.0815811
R28304 avss.n380 avss.n379 0.0815811
R28305 avss.n392 avss.n391 0.0815811
R28306 avss.n850 avss.n849 0.0798919
R28307 avss.n662 avss.n644 0.0794474
R28308 avss.n667 avss.n666 0.0794474
R28309 avss.n697 avss.n696 0.0794474
R28310 avss.n707 avss.n706 0.0794474
R28311 avss.n722 avss.n721 0.0794474
R28312 avss.n751 avss.n608 0.0794474
R28313 avss.n765 avss.n602 0.0794474
R28314 avss.n780 avss.n596 0.0794474
R28315 avss.n785 avss.n784 0.0794474
R28316 avss.n143 avss.n117 0.0793136
R28317 avss.n549 avss.n548 0.0784703
R28318 avss.n682 avss.n681 0.072046
R28319 avss.n739 avss.n737 0.072046
R28320 avss.n905 avss.n904 0.0674065
R28321 avss.n839 avss.n838 0.0674065
R28322 avss.n994 avss.n75 0.0674065
R28323 avss.n989 avss.n76 0.0674065
R28324 avss.n681 avss.n680 0.0671118
R28325 avss.n737 avss.n615 0.0671118
R28326 avss.n771 avss.n596 0.0638224
R28327 avss.n755 avss.n602 0.0621776
R28328 avss.n767 avss.n765 0.0555987
R28329 avss.n216 avss.n213 0.0553986
R28330 avss.n228 avss.n225 0.0553986
R28331 avss.n240 avss.n237 0.0553986
R28332 avss.n252 avss.n249 0.0553986
R28333 avss.n264 avss.n261 0.0553986
R28334 avss.n276 avss.n273 0.0553986
R28335 avss.n288 avss.n285 0.0553986
R28336 avss.n300 avss.n297 0.0553986
R28337 avss.n312 avss.n309 0.0553986
R28338 avss.n324 avss.n321 0.0553986
R28339 avss.n336 avss.n333 0.0553986
R28340 avss.n348 avss.n345 0.0553986
R28341 avss.n360 avss.n357 0.0553986
R28342 avss.n372 avss.n369 0.0553986
R28343 avss.n384 avss.n381 0.0553986
R28344 avss.n395 avss.n394 0.0553986
R28345 avss.n781 avss.n595 0.0539539
R28346 avss.n853 avss.n582 0.0539539
R28347 avss.n1085 avss.n17 0.0538514
R28348 avss.n849 avss.n804 0.0532162
R28349 avss.n666 avss.n635 0.0523092
R28350 avss.n687 avss.n686 0.0523092
R28351 avss.n701 avss.n626 0.0523092
R28352 avss.n723 avss.n722 0.0523092
R28353 avss.n738 avss.n613 0.0523092
R28354 avss.n752 avss.n607 0.0498421
R28355 avss.n663 avss.n642 0.047375
R28356 avss.n678 avss.n633 0.047375
R28357 avss.n696 avss.n628 0.047375
R28358 avss.n705 avss.n702 0.047375
R28359 avss.n727 avss.n724 0.047375
R28360 avss.n741 avss.n608 0.047375
R28361 avss.n653 avss.n652 0.0449079
R28362 avss.n772 avss.n601 0.0440855
R28363 avss.n872 avss.n871 0.0436892
R28364 avss.n1043 avss.n1042 0.0430541
R28365 avss.n1046 avss.n42 0.0430541
R28366 avss.n1051 avss.n1049 0.0430541
R28367 avss.n1068 avss.n1067 0.0430541
R28368 avss.n1071 avss.n29 0.0430541
R28369 avss.n1090 avss.n1089 0.0430541
R28370 avss.n868 avss.n866 0.0430541
R28371 avss.n665 avss.n642 0.0428468
R28372 avss.n702 avss.n620 0.0428468
R28373 avss.n1086 avss.n1085 0.0427365
R28374 avss.n125 avss 0.0410405
R28375 avss.n756 avss 0.0399737
R28376 avss.n785 avss 0.0399737
R28377 avss.n667 avss.n665 0.0379126
R28378 avss.n721 avss.n620 0.0379126
R28379 avss.n766 avss.n601 0.0358618
R28380 avss.n215 avss 0.0351284
R28381 avss.n227 avss 0.0351284
R28382 avss.n239 avss 0.0351284
R28383 avss.n251 avss 0.0351284
R28384 avss.n263 avss 0.0351284
R28385 avss.n275 avss 0.0351284
R28386 avss.n287 avss 0.0351284
R28387 avss.n299 avss 0.0351284
R28388 avss.n311 avss 0.0351284
R28389 avss.n323 avss 0.0351284
R28390 avss.n335 avss 0.0351284
R28391 avss.n347 avss 0.0351284
R28392 avss.n359 avss 0.0351284
R28393 avss.n371 avss 0.0351284
R28394 avss.n383 avss 0.0351284
R28395 avss avss.n0 0.0351284
R28396 avss.n652 avss.n644 0.0350395
R28397 avss avss.n783 0.0342171
R28398 avss.n852 avss 0.0342171
R28399 avss.n127 avss.n2 0.0334392
R28400 avss.n663 avss.n662 0.0325724
R28401 avss.n678 avss.n677 0.0325724
R28402 avss.n683 avss.n628 0.0325724
R28403 avss.n699 avss 0.0325724
R28404 avss.n706 avss.n705 0.0325724
R28405 avss.n728 avss.n727 0.0325724
R28406 avss.n742 avss.n741 0.0325724
R28407 avss.n752 avss.n751 0.0301053
R28408 avss avss.n754 0.0301053
R28409 avss.n677 avss.n635 0.0276382
R28410 avss.n686 avss.n683 0.0276382
R28411 avss avss.n698 0.0276382
R28412 avss.n707 avss.n701 0.0276382
R28413 avss.n728 avss.n723 0.0276382
R28414 avss.n742 avss.n613 0.0276382
R28415 avss.n127 avss.n126 0.0266824
R28416 avss.n213 avss.n212 0.0266824
R28417 avss.n225 avss.n224 0.0266824
R28418 avss.n237 avss.n236 0.0266824
R28419 avss.n249 avss.n248 0.0266824
R28420 avss.n261 avss.n260 0.0266824
R28421 avss.n273 avss.n272 0.0266824
R28422 avss.n285 avss.n284 0.0266824
R28423 avss.n297 avss.n296 0.0266824
R28424 avss.n309 avss.n308 0.0266824
R28425 avss.n321 avss.n320 0.0266824
R28426 avss.n333 avss.n332 0.0266824
R28427 avss.n345 avss.n344 0.0266824
R28428 avss.n357 avss.n356 0.0266824
R28429 avss.n369 avss.n368 0.0266824
R28430 avss.n381 avss.n380 0.0266824
R28431 avss.n394 avss.n392 0.0266824
R28432 avss.n781 avss.n780 0.0259934
R28433 avss.n784 avss.n582 0.0259934
R28434 avss.n1014 avss.n52 0.0258406
R28435 avss.n1017 avss.n1016 0.0258406
R28436 avss.n767 avss.n766 0.0243487
R28437 avss.n129 avss.n2 0.0224595
R28438 avss.n803 avss.n798 0.0190811
R28439 avss.n92 avss.n87 0.0190811
R28440 avss.n756 avss.n755 0.0177697
R28441 avss.n772 avss.n771 0.016125
R28442 avss.n653 avss.n650 0.0153026
R28443 avss.n680 avss.n633 0.0128355
R28444 avss.n698 avss.n697 0.0128355
R28445 avss.n724 avss.n615 0.0128355
R28446 avss.n754 avss.n607 0.0103684
R28447 avss.n687 avss.n682 0.00790132
R28448 avss.n699 avss.n626 0.00790132
R28449 avss.n739 avss.n738 0.00790132
R28450 avss.n216 avss.n215 0.00641216
R28451 avss.n228 avss.n227 0.00641216
R28452 avss.n240 avss.n239 0.00641216
R28453 avss.n252 avss.n251 0.00641216
R28454 avss.n264 avss.n263 0.00641216
R28455 avss.n276 avss.n275 0.00641216
R28456 avss.n288 avss.n287 0.00641216
R28457 avss.n300 avss.n299 0.00641216
R28458 avss.n312 avss.n311 0.00641216
R28459 avss.n324 avss.n323 0.00641216
R28460 avss.n336 avss.n335 0.00641216
R28461 avss.n348 avss.n347 0.00641216
R28462 avss.n360 avss.n359 0.00641216
R28463 avss.n372 avss.n371 0.00641216
R28464 avss.n384 avss.n383 0.00641216
R28465 avss.n395 avss.n0 0.00641216
R28466 avss.n783 avss.n595 0.00625658
R28467 avss.n853 avss.n852 0.00625658
R28468 avss.n1012 avss.n55 0.004875
R28469 por.n2 por.n0 243.458
R28470 por.n2 por.n1 205.059
R28471 por.n4 por.n3 205.059
R28472 por.n6 por.n5 205.059
R28473 por.n8 por.n7 205.059
R28474 por.n10 por.n9 205.059
R28475 por.n12 por.n11 205.059
R28476 por.n14 por.n13 205.059
R28477 por.n17 por.n15 133.534
R28478 por.n17 por.n16 99.1759
R28479 por.n19 por.n18 99.1759
R28480 por.n21 por.n20 99.1759
R28481 por.n23 por.n22 99.1759
R28482 por.n25 por.n24 99.1759
R28483 por.n27 por.n26 99.1759
R28484 por por.n28 97.4305
R28485 por.n4 por.n2 38.4005
R28486 por.n6 por.n4 38.4005
R28487 por.n8 por.n6 38.4005
R28488 por.n10 por.n8 38.4005
R28489 por.n12 por.n10 38.4005
R28490 por.n14 por.n12 38.4005
R28491 por.n19 por.n17 34.3584
R28492 por.n21 por.n19 34.3584
R28493 por.n23 por.n21 34.3584
R28494 por.n25 por.n23 34.3584
R28495 por.n27 por.n25 34.3584
R28496 por.n29 por.n27 34.3584
R28497 por.n13 por.t31 26.5955
R28498 por.n13 por.t18 26.5955
R28499 por.n0 por.t26 26.5955
R28500 por.n0 por.t30 26.5955
R28501 por.n1 por.t21 26.5955
R28502 por.n1 por.t29 26.5955
R28503 por.n3 por.t28 26.5955
R28504 por.n3 por.t24 26.5955
R28505 por.n5 por.t27 26.5955
R28506 por.n5 por.t25 26.5955
R28507 por.n7 por.t23 26.5955
R28508 por.n7 por.t20 26.5955
R28509 por.n9 por.t19 26.5955
R28510 por.n9 por.t17 26.5955
R28511 por.n11 por.t16 26.5955
R28512 por.n11 por.t22 26.5955
R28513 por.n28 por.t1 24.9236
R28514 por.n28 por.t4 24.9236
R28515 por.n15 por.t12 24.9236
R28516 por.n15 por.t0 24.9236
R28517 por.n16 por.t7 24.9236
R28518 por.n16 por.t15 24.9236
R28519 por.n18 por.t14 24.9236
R28520 por.n18 por.t10 24.9236
R28521 por.n20 por.t13 24.9236
R28522 por.n20 por.t11 24.9236
R28523 por.n22 por.t9 24.9236
R28524 por.n22 por.t6 24.9236
R28525 por.n24 por.t5 24.9236
R28526 por.n24 por.t3 24.9236
R28527 por.n26 por.t2 24.9236
R28528 por.n26 por.t8 24.9236
R28529 por.n30 por 24.0418
R28530 por por.n14 18.4247
R28531 por.n30 por.n29 10.0853
R28532 por.n29 por 1.74595
R28533 por por.n30 1.35808
R28534 osc_ck.n11 osc_ck.t6 236.258
R28535 osc_ck.n8 osc_ck.n6 214.567
R28536 osc_ck.n10 osc_ck.n5 207.792
R28537 osc_ck.n0 osc_ck.t13 184.768
R28538 osc_ck.n1 osc_ck.t9 184.768
R28539 osc_ck.n2 osc_ck.t14 184.768
R28540 osc_ck.n3 osc_ck.t10 184.768
R28541 osc_ck.n4 osc_ck.n3 171.375
R28542 osc_ck.n0 osc_ck.t11 146.208
R28543 osc_ck.n1 osc_ck.t15 146.208
R28544 osc_ck.n2 osc_ck.t12 146.208
R28545 osc_ck.n3 osc_ck.t8 146.208
R28546 osc_ck.n9 osc_ck.t5 88.3503
R28547 osc_ck.n12 osc_ck.n11 80.8585
R28548 osc_ck.n8 osc_ck.n7 70.9231
R28549 osc_ck.n1 osc_ck.n0 40.6397
R28550 osc_ck.n2 osc_ck.n1 40.6397
R28551 osc_ck.n3 osc_ck.n2 40.6397
R28552 osc_ck.n6 osc_ck.t2 29.5505
R28553 osc_ck.n6 osc_ck.t0 29.5505
R28554 osc_ck.n5 osc_ck.t4 28.5655
R28555 osc_ck.n5 osc_ck.t3 28.5655
R28556 osc_ck.n7 osc_ck.t1 18.0005
R28557 osc_ck.n7 osc_ck.t7 18.0005
R28558 osc_ck.n12 osc_ck 15.2808
R28559 osc_ck.n10 osc_ck.n9 13.4303
R28560 osc_ck osc_ck.n4 9.14336
R28561 osc_ck.n9 osc_ck.n8 7.92796
R28562 osc_ck.n4 osc_ck 4.67352
R28563 osc_ck osc_ck.n12 0.835533
R28564 osc_ck.n11 osc_ck.n10 0.0968612
R28565 por_dig_0.net23.n30 por_dig_0.net23.n1 589.152
R28566 por_dig_0.net23.n16 por_dig_0.net23.t19 471.289
R28567 por_dig_0.net23.n10 por_dig_0.net23.t4 241.536
R28568 por_dig_0.net23.n2 por_dig_0.net23.t17 238.194
R28569 por_dig_0.net23.n21 por_dig_0.net23.t8 236.18
R28570 por_dig_0.net23.n19 por_dig_0.net23.t22 231.017
R28571 por_dig_0.net23.n12 por_dig_0.net23.t11 231.017
R28572 por_dig_0.net23.n8 por_dig_0.net23.t12 231.017
R28573 por_dig_0.net23.n25 por_dig_0.net23.t23 224.984
R28574 por_dig_0.net23 por_dig_0.net23.n31 216.464
R28575 por_dig_0.net23.n25 por_dig_0.net23.t14 187.714
R28576 por_dig_0.net23.n14 por_dig_0.net23.t7 173.34
R28577 por_dig_0.net23.n4 por_dig_0.net23.t18 173.34
R28578 por_dig_0.net23.n10 por_dig_0.net23.t16 169.237
R28579 por_dig_0.net23.n2 por_dig_0.net23.t10 165.893
R28580 por_dig_0.net23.n21 por_dig_0.net23.t13 163.881
R28581 por_dig_0.net23.n14 por_dig_0.net23.t21 162.81
R28582 por_dig_0.net23.n4 por_dig_0.net23.t5 162.81
R28583 por_dig_0.net23.n17 por_dig_0.net23.n16 161.775
R28584 por_dig_0.net23 por_dig_0.net23.n14 159.565
R28585 por_dig_0.net23.n19 por_dig_0.net23.t9 158.716
R28586 por_dig_0.net23.n12 por_dig_0.net23.t15 158.716
R28587 por_dig_0.net23.n8 por_dig_0.net23.t6 158.716
R28588 por_dig_0.net23.n6 por_dig_0.net23.n4 156.268
R28589 por_dig_0.net23.n3 por_dig_0.net23.n2 153.477
R28590 por_dig_0.net23.n13 por_dig_0.net23.n12 153.358
R28591 por_dig_0.net23.n9 por_dig_0.net23.n8 153.303
R28592 por_dig_0.net23.n11 por_dig_0.net23.n10 153.26
R28593 por_dig_0.net23.n26 por_dig_0.net23.n25 152
R28594 por_dig_0.net23.n22 por_dig_0.net23.n21 152
R28595 por_dig_0.net23.n20 por_dig_0.net23.n19 152
R28596 por_dig_0.net23.n16 por_dig_0.net23.t20 148.35
R28597 por_dig_0.net23.n31 por_dig_0.net23.t0 38.5719
R28598 por_dig_0.net23.n31 por_dig_0.net23.t1 38.5719
R28599 por_dig_0.net23 por_dig_0.net23.n30 34.7569
R28600 por_dig_0.net23.n1 por_dig_0.net23.t3 26.5955
R28601 por_dig_0.net23.n1 por_dig_0.net23.t2 26.5955
R28602 por_dig_0.net23.n0 por_dig_0.net23.n15 25.5914
R28603 por_dig_0.net23.n7 por_dig_0.net23.n3 22.6426
R28604 por_dig_0.net23.n27 por_dig_0.net23 19.8943
R28605 por_dig_0.net23.n0 por_dig_0.net23.n13 19.6865
R28606 por_dig_0.net23.n22 por_dig_0.net23 16.5338
R28607 por_dig_0.net23.n23 por_dig_0.net23.n20 15.1342
R28608 por_dig_0.net23.n18 por_dig_0.net23.n17 14.5053
R28609 por_dig_0.net23.n23 por_dig_0.net23.n22 14.4719
R28610 por_dig_0.net23.n29 por_dig_0.net23.n7 12.9649
R28611 por_dig_0.net23 por_dig_0.net23.n11 12.0867
R28612 por_dig_0.net23.n29 por_dig_0.net23.n28 11.2972
R28613 por_dig_0.net23.n28 por_dig_0.net23.n27 10.9511
R28614 por_dig_0.net23.n18 por_dig_0.net23.n0 10.4613
R28615 por_dig_0.net23.n28 por_dig_0.net23.n9 10.1368
R28616 por_dig_0.net23.n30 por_dig_0.net23.n29 9.59462
R28617 por_dig_0.net23.n7 por_dig_0.net23.n6 9.3005
R28618 por_dig_0.net23.n6 por_dig_0.net23.n5 8.92171
R28619 por_dig_0.net23.n15 por_dig_0.net23 8.43686
R28620 por_dig_0.net23 por_dig_0.net23.n26 8.0005
R28621 por_dig_0.net23.n24 por_dig_0.net23.n23 6.89885
R28622 por_dig_0.net23.n15 por_dig_0.net23 5.62474
R28623 por_dig_0.net23.n3 por_dig_0.net23 4.18512
R28624 por_dig_0.net23.n26 por_dig_0.net23 4.08939
R28625 por_dig_0.net23.n17 por_dig_0.net23 3.95686
R28626 por_dig_0.net23.n9 por_dig_0.net23 3.68864
R28627 por_dig_0.net23.n11 por_dig_0.net23 3.56771
R28628 por_dig_0.net23.n13 por_dig_0.net23 3.29747
R28629 por_dig_0.net23.n24 por_dig_0.net23.n18 2.60077
R28630 por_dig_0.net23.n5 por_dig_0.net23 2.37576
R28631 por_dig_0.net23.n20 por_dig_0.net23 2.32777
R28632 por_dig_0.net23.n0 por_dig_0.net23 2.19624
R28633 por_dig_0.net23.n27 por_dig_0.net23.n24 1.99363
R28634 por_dig_0.net23.n5 por_dig_0.net23 0.970197
R28635 por_ana_0.comparator_1.vpp.t16 por_ana_0.comparator_1.vpp.n2 241.742
R28636 por_ana_0.comparator_1.vpp.n2 por_ana_0.comparator_1.vpp.n9 204.284
R28637 por_ana_0.comparator_1.vpp.n2 por_ana_0.comparator_1.vpp.n23 204.284
R28638 por_ana_0.comparator_1.vpp.n2 por_ana_0.comparator_1.vpp.n22 204.284
R28639 por_ana_0.comparator_1.vpp.n2 por_ana_0.comparator_1.vpp.n21 204.284
R28640 por_ana_0.comparator_1.vpp.n2 por_ana_0.comparator_1.vpp.n20 204.284
R28641 por_ana_0.comparator_1.vpp.n2 por_ana_0.comparator_1.vpp.n19 204.284
R28642 por_ana_0.comparator_1.vpp.n2 por_ana_0.comparator_1.vpp.n18 204.284
R28643 por_ana_0.comparator_1.vpp.n2 por_ana_0.comparator_1.vpp.n6 199.786
R28644 por_ana_0.comparator_1.vpp.n2 por_ana_0.comparator_1.vpp.n5 199.65
R28645 por_ana_0.comparator_1.vpp.n2 por_ana_0.comparator_1.vpp.n7 199.65
R28646 por_ana_0.comparator_1.vpp.n2 por_ana_0.comparator_1.vpp.n8 199.65
R28647 por_ana_0.comparator_1.vpp.n1 por_ana_0.comparator_1.vpp.n10 71.9371
R28648 por_ana_0.comparator_1.vpp.n1 por_ana_0.comparator_1.vpp.n17 70.9612
R28649 por_ana_0.comparator_1.vpp.n1 por_ana_0.comparator_1.vpp.n16 70.9612
R28650 por_ana_0.comparator_1.vpp.n1 por_ana_0.comparator_1.vpp.n15 70.9612
R28651 por_ana_0.comparator_1.vpp.n1 por_ana_0.comparator_1.vpp.n14 70.9612
R28652 por_ana_0.comparator_1.vpp.n1 por_ana_0.comparator_1.vpp.n13 70.9612
R28653 por_ana_0.comparator_1.vpp.n1 por_ana_0.comparator_1.vpp.n12 70.9612
R28654 por_ana_0.comparator_1.vpp.n1 por_ana_0.comparator_1.vpp.n11 70.9612
R28655 por_ana_0.comparator_1.vpp.n6 por_ana_0.comparator_1.vpp.t13 27.6955
R28656 por_ana_0.comparator_1.vpp.n6 por_ana_0.comparator_1.vpp.t9 27.6955
R28657 por_ana_0.comparator_1.vpp.n5 por_ana_0.comparator_1.vpp.t5 27.6955
R28658 por_ana_0.comparator_1.vpp.n5 por_ana_0.comparator_1.vpp.t1 27.6955
R28659 por_ana_0.comparator_1.vpp.n7 por_ana_0.comparator_1.vpp.t11 27.6955
R28660 por_ana_0.comparator_1.vpp.n7 por_ana_0.comparator_1.vpp.t7 27.6955
R28661 por_ana_0.comparator_1.vpp.n8 por_ana_0.comparator_1.vpp.t3 27.6955
R28662 por_ana_0.comparator_1.vpp.n8 por_ana_0.comparator_1.vpp.t15 27.6955
R28663 por_ana_0.comparator_1.vpp.n9 por_ana_0.comparator_1.vpp.t24 27.6955
R28664 por_ana_0.comparator_1.vpp.n9 por_ana_0.comparator_1.vpp.t25 27.6955
R28665 por_ana_0.comparator_1.vpp.n23 por_ana_0.comparator_1.vpp.t26 27.6955
R28666 por_ana_0.comparator_1.vpp.n23 por_ana_0.comparator_1.vpp.t17 27.6955
R28667 por_ana_0.comparator_1.vpp.n22 por_ana_0.comparator_1.vpp.t27 27.6955
R28668 por_ana_0.comparator_1.vpp.n22 por_ana_0.comparator_1.vpp.t18 27.6955
R28669 por_ana_0.comparator_1.vpp.n21 por_ana_0.comparator_1.vpp.t28 27.6955
R28670 por_ana_0.comparator_1.vpp.n21 por_ana_0.comparator_1.vpp.t19 27.6955
R28671 por_ana_0.comparator_1.vpp.n20 por_ana_0.comparator_1.vpp.t29 27.6955
R28672 por_ana_0.comparator_1.vpp.n20 por_ana_0.comparator_1.vpp.t20 27.6955
R28673 por_ana_0.comparator_1.vpp.n19 por_ana_0.comparator_1.vpp.t22 27.6955
R28674 por_ana_0.comparator_1.vpp.n19 por_ana_0.comparator_1.vpp.t23 27.6955
R28675 por_ana_0.comparator_1.vpp.n18 por_ana_0.comparator_1.vpp.t30 27.6955
R28676 por_ana_0.comparator_1.vpp.n18 por_ana_0.comparator_1.vpp.t21 27.6955
R28677 por_ana_0.comparator_1.vpp.n1 por_ana_0.comparator_1.vpp.t59 23.5879
R28678 por_ana_0.comparator_1.vpp.n2 por_ana_0.comparator_1.vpp.n1 18.1658
R28679 por_ana_0.comparator_1.vpp.n1 por_ana_0.comparator_1.vpp.n0 18.106
R28680 por_ana_0.comparator_1.vpp.n1 por_ana_0.comparator_1.vpp.n3 16.9748
R28681 por_ana_0.comparator_1.vpp.n17 por_ana_0.comparator_1.vpp.t34 16.5305
R28682 por_ana_0.comparator_1.vpp.n17 por_ana_0.comparator_1.vpp.t39 16.5305
R28683 por_ana_0.comparator_1.vpp.n16 por_ana_0.comparator_1.vpp.t43 16.5305
R28684 por_ana_0.comparator_1.vpp.n16 por_ana_0.comparator_1.vpp.t31 16.5305
R28685 por_ana_0.comparator_1.vpp.n15 por_ana_0.comparator_1.vpp.t35 16.5305
R28686 por_ana_0.comparator_1.vpp.n15 por_ana_0.comparator_1.vpp.t40 16.5305
R28687 por_ana_0.comparator_1.vpp.n14 por_ana_0.comparator_1.vpp.t38 16.5305
R28688 por_ana_0.comparator_1.vpp.n14 por_ana_0.comparator_1.vpp.t46 16.5305
R28689 por_ana_0.comparator_1.vpp.n13 por_ana_0.comparator_1.vpp.t36 16.5305
R28690 por_ana_0.comparator_1.vpp.n13 por_ana_0.comparator_1.vpp.t41 16.5305
R28691 por_ana_0.comparator_1.vpp.n12 por_ana_0.comparator_1.vpp.t44 16.5305
R28692 por_ana_0.comparator_1.vpp.n12 por_ana_0.comparator_1.vpp.t32 16.5305
R28693 por_ana_0.comparator_1.vpp.n11 por_ana_0.comparator_1.vpp.t37 16.5305
R28694 por_ana_0.comparator_1.vpp.n11 por_ana_0.comparator_1.vpp.t42 16.5305
R28695 por_ana_0.comparator_1.vpp.n10 por_ana_0.comparator_1.vpp.t45 16.5305
R28696 por_ana_0.comparator_1.vpp.n10 por_ana_0.comparator_1.vpp.t33 16.5305
R28697 por_ana_0.comparator_1.vpp.n0 por_ana_0.comparator_1.vpp.t62 16.3148
R28698 por_ana_0.comparator_1.vpp.n0 por_ana_0.comparator_1.vpp.t50 16.3148
R28699 por_ana_0.comparator_1.vpp.n4 por_ana_0.comparator_1.vpp.t51 16.3148
R28700 por_ana_0.comparator_1.vpp.n0 por_ana_0.comparator_1.vpp.t52 16.3148
R28701 por_ana_0.comparator_1.vpp.n0 por_ana_0.comparator_1.vpp.t53 16.3148
R28702 por_ana_0.comparator_1.vpp.n1 por_ana_0.comparator_1.vpp.t60 16.3148
R28703 por_ana_0.comparator_1.vpp.n1 por_ana_0.comparator_1.vpp.t54 16.3148
R28704 por_ana_0.comparator_1.vpp.n3 por_ana_0.comparator_1.vpp.t47 16.3148
R28705 por_ana_0.comparator_1.vpp.n2 por_ana_0.comparator_1.vpp.t14 14.2251
R28706 por_ana_0.comparator_1.vpp.n2 por_ana_0.comparator_1.vpp.t2 14.2251
R28707 por_ana_0.comparator_1.vpp.n2 por_ana_0.comparator_1.vpp.t6 14.2251
R28708 por_ana_0.comparator_1.vpp.n2 por_ana_0.comparator_1.vpp.t10 14.2251
R28709 por_ana_0.comparator_1.vpp.n2 por_ana_0.comparator_1.vpp.t0 14.2251
R28710 por_ana_0.comparator_1.vpp.n2 por_ana_0.comparator_1.vpp.t4 14.2251
R28711 por_ana_0.comparator_1.vpp.n2 por_ana_0.comparator_1.vpp.t12 14.2251
R28712 por_ana_0.comparator_1.vpp.n2 por_ana_0.comparator_1.vpp.t8 14.2251
R28713 por_ana_0.comparator_1.vpp.n0 por_ana_0.comparator_1.vpp.n4 14.2134
R28714 por_ana_0.comparator_1.vpp.n0 por_ana_0.comparator_1.vpp.t48 12.0866
R28715 por_ana_0.comparator_1.vpp.n0 por_ana_0.comparator_1.vpp.t55 12.0866
R28716 por_ana_0.comparator_1.vpp.n4 por_ana_0.comparator_1.vpp.t56 12.0866
R28717 por_ana_0.comparator_1.vpp.n0 por_ana_0.comparator_1.vpp.t57 12.0866
R28718 por_ana_0.comparator_1.vpp.n0 por_ana_0.comparator_1.vpp.t58 12.0866
R28719 por_ana_0.comparator_1.vpp.n1 por_ana_0.comparator_1.vpp.t61 12.0866
R28720 por_ana_0.comparator_1.vpp.n3 por_ana_0.comparator_1.vpp.t49 12.0866
R28721 dcomp.n2 dcomp.n0 243.458
R28722 dcomp.n2 dcomp.n1 205.059
R28723 dcomp.n4 dcomp.n3 205.059
R28724 dcomp.n6 dcomp.n5 205.059
R28725 dcomp.n8 dcomp.n7 205.059
R28726 dcomp.n10 dcomp.n9 205.059
R28727 dcomp.n12 dcomp.n11 205.059
R28728 dcomp.n14 dcomp.n13 205.059
R28729 dcomp.n17 dcomp.n15 133.534
R28730 dcomp.n17 dcomp.n16 99.1759
R28731 dcomp.n19 dcomp.n18 99.1759
R28732 dcomp.n21 dcomp.n20 99.1759
R28733 dcomp.n23 dcomp.n22 99.1759
R28734 dcomp.n25 dcomp.n24 99.1759
R28735 dcomp.n27 dcomp.n26 99.1759
R28736 dcomp dcomp.n28 97.4305
R28737 dcomp.n4 dcomp.n2 38.4005
R28738 dcomp.n6 dcomp.n4 38.4005
R28739 dcomp.n8 dcomp.n6 38.4005
R28740 dcomp.n10 dcomp.n8 38.4005
R28741 dcomp.n12 dcomp.n10 38.4005
R28742 dcomp.n14 dcomp.n12 38.4005
R28743 dcomp.n19 dcomp.n17 34.3584
R28744 dcomp.n21 dcomp.n19 34.3584
R28745 dcomp.n23 dcomp.n21 34.3584
R28746 dcomp.n25 dcomp.n23 34.3584
R28747 dcomp.n27 dcomp.n25 34.3584
R28748 dcomp.n29 dcomp.n27 34.3584
R28749 dcomp.n30 dcomp 32.7152
R28750 dcomp.n13 dcomp.t17 26.5955
R28751 dcomp.n13 dcomp.t20 26.5955
R28752 dcomp.n0 dcomp.t28 26.5955
R28753 dcomp.n0 dcomp.t16 26.5955
R28754 dcomp.n1 dcomp.t23 26.5955
R28755 dcomp.n1 dcomp.t31 26.5955
R28756 dcomp.n3 dcomp.t30 26.5955
R28757 dcomp.n3 dcomp.t26 26.5955
R28758 dcomp.n5 dcomp.t29 26.5955
R28759 dcomp.n5 dcomp.t27 26.5955
R28760 dcomp.n7 dcomp.t25 26.5955
R28761 dcomp.n7 dcomp.t22 26.5955
R28762 dcomp.n9 dcomp.t21 26.5955
R28763 dcomp.n9 dcomp.t19 26.5955
R28764 dcomp.n11 dcomp.t18 26.5955
R28765 dcomp.n11 dcomp.t24 26.5955
R28766 dcomp.n28 dcomp.t7 24.9236
R28767 dcomp.n28 dcomp.t10 24.9236
R28768 dcomp.n15 dcomp.t2 24.9236
R28769 dcomp.n15 dcomp.t6 24.9236
R28770 dcomp.n16 dcomp.t13 24.9236
R28771 dcomp.n16 dcomp.t5 24.9236
R28772 dcomp.n18 dcomp.t4 24.9236
R28773 dcomp.n18 dcomp.t0 24.9236
R28774 dcomp.n20 dcomp.t3 24.9236
R28775 dcomp.n20 dcomp.t1 24.9236
R28776 dcomp.n22 dcomp.t15 24.9236
R28777 dcomp.n22 dcomp.t12 24.9236
R28778 dcomp.n24 dcomp.t11 24.9236
R28779 dcomp.n24 dcomp.t9 24.9236
R28780 dcomp.n26 dcomp.t8 24.9236
R28781 dcomp.n26 dcomp.t14 24.9236
R28782 dcomp dcomp.n14 18.4247
R28783 dcomp.n30 dcomp.n29 10.0853
R28784 dcomp.n29 dcomp 1.74595
R28785 dcomp dcomp.n30 1.35808
R28786 por_ana_0.rstring_mux_0.vtrip3.n5 por_ana_0.rstring_mux_0.vtrip3.n3 50.7022
R28787 por_ana_0.rstring_mux_0.vtrip3.n2 por_ana_0.rstring_mux_0.vtrip3.n0 50.7022
R28788 por_ana_0.rstring_mux_0.vtrip3.n6 por_ana_0.rstring_mux_0.vtrip3.n5 14.2209
R28789 por_ana_0.rstring_mux_0.vtrip3.n5 por_ana_0.rstring_mux_0.vtrip3.n4 13.8791
R28790 por_ana_0.rstring_mux_0.vtrip3.n2 por_ana_0.rstring_mux_0.vtrip3.n1 13.8791
R28791 por_ana_0.rstring_mux_0.vtrip3.t4 por_ana_0.rstring_mux_0.vtrip3.n7 10.5857
R28792 por_ana_0.rstring_mux_0.vtrip3.n7 por_ana_0.rstring_mux_0.vtrip3.t9 10.5847
R28793 por_ana_0.rstring_mux_0.vtrip3.n6 por_ana_0.rstring_mux_0.vtrip3.n2 5.7125
R28794 por_ana_0.rstring_mux_0.vtrip3.n3 por_ana_0.rstring_mux_0.vtrip3.t3 5.5395
R28795 por_ana_0.rstring_mux_0.vtrip3.n3 por_ana_0.rstring_mux_0.vtrip3.t2 5.5395
R28796 por_ana_0.rstring_mux_0.vtrip3.n0 por_ana_0.rstring_mux_0.vtrip3.t7 5.5395
R28797 por_ana_0.rstring_mux_0.vtrip3.n0 por_ana_0.rstring_mux_0.vtrip3.t8 5.5395
R28798 por_ana_0.rstring_mux_0.vtrip3.n4 por_ana_0.rstring_mux_0.vtrip3.t1 3.3065
R28799 por_ana_0.rstring_mux_0.vtrip3.n4 por_ana_0.rstring_mux_0.vtrip3.t0 3.3065
R28800 por_ana_0.rstring_mux_0.vtrip3.n1 por_ana_0.rstring_mux_0.vtrip3.t5 3.3065
R28801 por_ana_0.rstring_mux_0.vtrip3.n1 por_ana_0.rstring_mux_0.vtrip3.t6 3.3065
R28802 por_ana_0.rstring_mux_0.vtrip3.n7 por_ana_0.rstring_mux_0.vtrip3.n6 3.16869
R28803 por_ana_0.rstring_mux_0.vtrip2.n5 por_ana_0.rstring_mux_0.vtrip2.n3 50.7022
R28804 por_ana_0.rstring_mux_0.vtrip2.n2 por_ana_0.rstring_mux_0.vtrip2.n0 50.7022
R28805 por_ana_0.rstring_mux_0.vtrip2.n7 por_ana_0.rstring_mux_0.vtrip2.n6 23.8383
R28806 por_ana_0.rstring_mux_0.vtrip2.n6 por_ana_0.rstring_mux_0.vtrip2.n5 14.3726
R28807 por_ana_0.rstring_mux_0.vtrip2.n5 por_ana_0.rstring_mux_0.vtrip2.n4 13.8791
R28808 por_ana_0.rstring_mux_0.vtrip2.n2 por_ana_0.rstring_mux_0.vtrip2.n1 13.8791
R28809 por_ana_0.rstring_mux_0.vtrip2.n7 por_ana_0.rstring_mux_0.vtrip2.t5 10.6303
R28810 por_ana_0.rstring_mux_0.vtrip2.n3 por_ana_0.rstring_mux_0.vtrip2.t9 5.5395
R28811 por_ana_0.rstring_mux_0.vtrip2.n3 por_ana_0.rstring_mux_0.vtrip2.t8 5.5395
R28812 por_ana_0.rstring_mux_0.vtrip2.n0 por_ana_0.rstring_mux_0.vtrip2.t6 5.5395
R28813 por_ana_0.rstring_mux_0.vtrip2.n0 por_ana_0.rstring_mux_0.vtrip2.t7 5.5395
R28814 por_ana_0.rstring_mux_0.vtrip2.n6 por_ana_0.rstring_mux_0.vtrip2.n2 4.21994
R28815 por_ana_0.rstring_mux_0.vtrip2.n4 por_ana_0.rstring_mux_0.vtrip2.t4 3.3065
R28816 por_ana_0.rstring_mux_0.vtrip2.n4 por_ana_0.rstring_mux_0.vtrip2.t3 3.3065
R28817 por_ana_0.rstring_mux_0.vtrip2.n1 por_ana_0.rstring_mux_0.vtrip2.t0 3.3065
R28818 por_ana_0.rstring_mux_0.vtrip2.n1 por_ana_0.rstring_mux_0.vtrip2.t1 3.3065
R28819 por_ana_0.rstring_mux_0.vtrip2 por_ana_0.rstring_mux_0.vtrip2.t2 0.769662
R28820 por_ana_0.rstring_mux_0.vtrip2 por_ana_0.rstring_mux_0.vtrip2.n7 0.0563195
R28821 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[6].n1 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[6].n0 873.303
R28822 por_ana_0.sky130_fd_sc_hvl__lsbuflv2hv_1_0[0|7].X por_ana_0.rstring_mux_0.vtrip_decoded_avdd[6].n1 585
R28823 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[6].t0 por_ana_0.sky130_fd_sc_hvl__lsbuflv2hv_1_0[0|7].X 511.971
R28824 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[6].n2 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[6].t3 384.704
R28825 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[6].n2 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[6].t4 384.226
R28826 por_ana_0.sky130_fd_sc_hvl__lsbuflv2hv_1_0[0|7].X por_ana_0.rstring_mux_0.vtrip_decoded_avdd[6].t1 155.607
R28827 por_ana_0.rstring_mux_0.sky130_fd_sc_hvl__inv_1_0[14].A por_ana_0.rstring_mux_0.vtrip_decoded_avdd[6].n3 153.165
R28828 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[6].n1 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[6].t0 147.756
R28829 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[6].n3 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[6].t2 114.031
R28830 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[6].n3 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[6].t5 81.5883
R28831 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[6].n6 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[6].n5 37.3303
R28832 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[6].n5 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[6].n4 13.8005
R28833 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[6].n5 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[6].n2 9.66769
R28834 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[6].n0 por_ana_0.sky130_fd_sc_hvl__lsbuflv2hv_1_0[0|7].X 8.85549
R28835 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[6].n4 por_ana_0.rstring_mux_0.sky130_fd_sc_hvl__inv_1_0[14].A 7.97972
R28836 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[6].n4 por_ana_0.rstring_mux_0.sky130_fd_sc_hvl__inv_1_0[14].A 7.97972
R28837 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[6].n6 por_ana_0.sky130_fd_sc_hvl__lsbuflv2hv_1_0[0|7].X 7.49318
R28838 por_ana_0.sky130_fd_sc_hvl__lsbuflv2hv_1_0[0|7].X por_ana_0.rstring_mux_0.vtrip_decoded_avdd[6].n0 4.05904
R28839 por_ana_0.sky130_fd_sc_hvl__lsbuflv2hv_1_0[0|7].X por_ana_0.rstring_mux_0.vtrip_decoded_avdd[6].n6 4.05904
R28840 por_dig_0._034_.n6 por_dig_0._034_.t13 241.536
R28841 por_dig_0._034_.n14 por_dig_0._034_.n12 235.923
R28842 por_dig_0._034_.n4 por_dig_0._034_.t15 231.835
R28843 por_dig_0._034_.n9 por_dig_0._034_.t10 229.001
R28844 por_dig_0._034_.n14 por_dig_0._034_.n13 206.25
R28845 por_dig_0._034_.n2 por_dig_0._034_.n0 204.565
R28846 por_dig_0._034_ por_dig_0._034_.n1 199.148
R28847 por_dig_0._034_.n11 por_dig_0._034_.n3 190.911
R28848 por_dig_0._034_.n6 por_dig_0._034_.t11 169.237
R28849 por_dig_0._034_.n4 por_dig_0._034_.t12 157.07
R28850 por_dig_0._034_.n9 por_dig_0._034_.t14 156.702
R28851 por_dig_0._034_.n7 por_dig_0._034_.n6 153.745
R28852 por_dig_0._034_.n10 por_dig_0._034_.n9 152
R28853 por_dig_0._034_.n5 por_dig_0._034_.n4 152
R28854 por_dig_0._034_.n11 por_dig_0._034_ 50.2687
R28855 por_dig_0._034_.n15 por_dig_0._034_.n14 38.9823
R28856 por_dig_0._034_ por_dig_0._034_.n2 26.7641
R28857 por_dig_0._034_.n0 por_dig_0._034_.t7 26.5955
R28858 por_dig_0._034_.n0 por_dig_0._034_.t6 26.5955
R28859 por_dig_0._034_.n3 por_dig_0._034_.t2 26.5955
R28860 por_dig_0._034_.n3 por_dig_0._034_.t3 26.5955
R28861 por_dig_0._034_.n12 por_dig_0._034_.t8 26.5955
R28862 por_dig_0._034_.n12 por_dig_0._034_.t9 26.5955
R28863 por_dig_0._034_.n13 por_dig_0._034_.t1 26.5955
R28864 por_dig_0._034_.n13 por_dig_0._034_.t0 26.5955
R28865 por_dig_0._034_.n8 por_dig_0._034_.n5 25.2315
R28866 por_dig_0._034_.n1 por_dig_0._034_.t5 24.9236
R28867 por_dig_0._034_.n1 por_dig_0._034_.t4 24.9236
R28868 por_dig_0._034_.n15 por_dig_0._034_.n11 15.34
R28869 por_dig_0._034_.n15 por_dig_0._034_ 13.0914
R28870 por_dig_0._034_ por_dig_0._034_.n10 10.8774
R28871 por_dig_0._034_.n10 por_dig_0._034_ 10.6672
R28872 por_dig_0._034_.n8 por_dig_0._034_.n7 9.3005
R28873 por_dig_0._034_ por_dig_0._034_.n15 4.26717
R28874 por_dig_0._034_.n7 por_dig_0._034_ 3.49141
R28875 por_dig_0._034_.n2 por_dig_0._034_ 2.53744
R28876 por_dig_0._034_.n5 por_dig_0._034_ 2.3045
R28877 por_dig_0._034_ por_dig_0._034_.n8 1.65091
R28878 por_ana_0.ibias_gen_0.vp.n10 por_ana_0.ibias_gen_0.vp.t6 56.5501
R28879 por_ana_0.ibias_gen_0.vp.n4 por_ana_0.ibias_gen_0.vp.t8 50.9767
R28880 por_ana_0.ibias_gen_0.vp.n5 por_ana_0.ibias_gen_0.vp.t8 50.9767
R28881 por_ana_0.ibias_gen_0.vp.t11 por_ana_0.ibias_gen_0.vp.n6 50.9767
R28882 por_ana_0.ibias_gen_0.vp.t7 por_ana_0.ibias_gen_0.vp.n4 48.6451
R28883 por_ana_0.ibias_gen_0.vp.n7 por_ana_0.ibias_gen_0.vp.t11 48.6451
R28884 por_ana_0.ibias_gen_0.vp.n6 por_ana_0.ibias_gen_0.vp.t10 48.6451
R28885 por_ana_0.ibias_gen_0.vp.n5 por_ana_0.ibias_gen_0.vp.t7 48.6451
R28886 por_ana_0.ibias_gen_0.vp.t10 por_ana_0.ibias_gen_0.vp.n3 48.6451
R28887 por_ana_0.ibias_gen_0.vp.n0 por_ana_0.ibias_gen_0.vp.n11 42.5266
R28888 por_ana_0.ibias_gen_0.vp.n0 por_ana_0.ibias_gen_0.vp.n2 42.4505
R28889 por_ana_0.ibias_gen_0.vp.n9 por_ana_0.ibias_gen_0.vp.n8 26.1532
R28890 por_ana_0.ibias_gen_0.vp.n8 por_ana_0.ibias_gen_0.vp.t9 25.4891
R28891 por_ana_0.ibias_gen_0.vp.n8 por_ana_0.ibias_gen_0.vp.t12 24.3233
R28892 por_ana_0.ibias_gen_0.vp.n13 por_ana_0.ibias_gen_0.vp.n12 15.1165
R28893 por_ana_0.ibias_gen_0.vp.n12 por_ana_0.ibias_gen_0.vp.n1 14.8365
R28894 por_ana_0.ibias_gen_0.vp.n10 por_ana_0.ibias_gen_0.vp.n9 8.08875
R28895 por_ana_0.ibias_gen_0.vp.n12 por_ana_0.ibias_gen_0.vp.n0 7.57893
R28896 por_ana_0.ibias_gen_0.vp.n0 por_ana_0.ibias_gen_0.vp.n10 6.28836
R28897 por_ana_0.ibias_gen_0.vp.n2 por_ana_0.ibias_gen_0.vp.t2 5.5395
R28898 por_ana_0.ibias_gen_0.vp.t0 por_ana_0.ibias_gen_0.vp.n2 5.5395
R28899 por_ana_0.ibias_gen_0.vp.n11 por_ana_0.ibias_gen_0.vp.t0 5.5395
R28900 por_ana_0.ibias_gen_0.vp.n11 por_ana_0.ibias_gen_0.vp.t4 5.5395
R28901 por_ana_0.ibias_gen_0.vp.n1 por_ana_0.ibias_gen_0.vp.t5 3.3065
R28902 por_ana_0.ibias_gen_0.vp.t1 por_ana_0.ibias_gen_0.vp.n1 3.3065
R28903 por_ana_0.ibias_gen_0.vp.t1 por_ana_0.ibias_gen_0.vp.n13 3.3065
R28904 por_ana_0.ibias_gen_0.vp.n13 por_ana_0.ibias_gen_0.vp.t3 3.3065
R28905 por_ana_0.ibias_gen_0.vp.n9 por_ana_0.ibias_gen_0.vp.n7 2.37524
R28906 por_ana_0.ibias_gen_0.vp.n6 por_ana_0.ibias_gen_0.vp.n5 2.33202
R28907 por_ana_0.ibias_gen_0.vp.n4 por_ana_0.ibias_gen_0.vp.n3 2.33202
R28908 por_ana_0.ibias_gen_0.vp.n7 por_ana_0.ibias_gen_0.vp.n3 2.33126
R28909 por_ana_0.ibias_gen_0.ibias0.n0 por_ana_0.ibias_gen_0.ibias0.t2 233.487
R28910 por_ana_0.ibias_gen_0.ibias0.n0 por_ana_0.ibias_gen_0.ibias0.t3 88.1251
R28911 por_ana_0.ibias_gen_0.ibias0.n1 por_ana_0.ibias_gen_0.ibias0.n0 71.4893
R28912 por_ana_0.ibias_gen_0.ibias0.t1 por_ana_0.ibias_gen_0.ibias0.n1 5.5395
R28913 por_ana_0.ibias_gen_0.ibias0.n1 por_ana_0.ibias_gen_0.ibias0.t0 5.5395
R28914 force_short_oneshot.n0 force_short_oneshot.t2 276.464
R28915 force_short_oneshot.n0 force_short_oneshot.t3 196.131
R28916 force_short_oneshot.n1 force_short_oneshot.n0 153.083
R28917 force_short_oneshot.n3 force_short_oneshot.n2 92.6423
R28918 force_short_oneshot.n2 force_short_oneshot.t0 16.5305
R28919 force_short_oneshot.n2 force_short_oneshot.t1 16.5305
R28920 force_short_oneshot force_short_oneshot.n1 9.39918
R28921 force_short_oneshot.n1 force_short_oneshot 3.06529
R28922 force_short_oneshot.n3 force_short_oneshot 0.904467
R28923 force_short_oneshot force_short_oneshot.n3 0.6585
R28924 por_dig_0.net7.n2 por_dig_0.net7.t15 323.55
R28925 por_dig_0.net7.n1 por_dig_0.net7.t1 319.171
R28926 por_dig_0.net7.n18 por_dig_0.net7.t13 241.536
R28927 por_dig_0.net7.n16 por_dig_0.net7.t2 241.536
R28928 por_dig_0.net7.n6 por_dig_0.net7.t11 229.001
R28929 por_dig_0.net7 por_dig_0.net7.t0 209.923
R28930 por_dig_0.net7.n12 por_dig_0.net7.t18 204.656
R28931 por_dig_0.net7.n8 por_dig_0.net7.t8 201.369
R28932 por_dig_0.net7.n15 por_dig_0.net7.t7 196.549
R28933 por_dig_0.net7.n5 por_dig_0.net7.t5 196.549
R28934 por_dig_0.net7.n2 por_dig_0.net7.t12 195.017
R28935 por_dig_0.net7.n21 por_dig_0.net7.t3 183.505
R28936 por_dig_0.net7.n18 por_dig_0.net7.t19 169.237
R28937 por_dig_0.net7.n16 por_dig_0.net7.t16 169.237
R28938 por_dig_0.net7 por_dig_0.net7.n15 159.024
R28939 por_dig_0.net7 por_dig_0.net7.n5 159.024
R28940 por_dig_0.net7.n6 por_dig_0.net7.t17 156.702
R28941 por_dig_0.net7 por_dig_0.net7.n16 156.329
R28942 por_dig_0.net7.n22 por_dig_0.net7.n21 153.863
R28943 por_dig_0.net7 por_dig_0.net7.n2 153.409
R28944 por_dig_0.net7.n14 por_dig_0.net7.n11 153.13
R28945 por_dig_0.net7.n9 por_dig_0.net7.n8 152.827
R28946 por_dig_0.net7.n19 por_dig_0.net7.n18 152
R28947 por_dig_0.net7.n13 por_dig_0.net7.n12 152
R28948 por_dig_0.net7.n7 por_dig_0.net7.n6 152
R28949 por_dig_0.net7.n15 por_dig_0.net7.t4 148.35
R28950 por_dig_0.net7.n5 por_dig_0.net7.t14 148.35
R28951 por_dig_0.net7.n8 por_dig_0.net7.t9 132.282
R28952 por_dig_0.net7.n11 por_dig_0.net7.t6 121.109
R28953 por_dig_0.net7.n21 por_dig_0.net7.t10 114.532
R28954 por_dig_0.net7.n12 por_dig_0.net7.n11 40.9982
R28955 por_dig_0.net7.n20 por_dig_0.net7.n19 23.2299
R28956 por_dig_0.net7.n17 por_dig_0.net7 18.9005
R28957 por_dig_0.net7.n7 por_dig_0.net7 18.7264
R28958 por_dig_0.net7.n0 por_dig_0.net7 16.4928
R28959 por_dig_0.net7.n4 por_dig_0.net7 16.0005
R28960 por_dig_0.net7 por_dig_0.net7.n22 13.8485
R28961 por_dig_0.net7.n0 por_dig_0.net7 11.9542
R28962 por_dig_0.net7.n10 por_dig_0.net7.n9 11.2528
R28963 por_dig_0.net7.n20 por_dig_0.net7.n17 11.1609
R28964 por_dig_0.net7.n0 por_dig_0.net7.n10 10.8257
R28965 por_dig_0.net7.n10 por_dig_0.net7.n7 10.7227
R28966 por_dig_0.net7.n0 por_dig_0.net7.n14 10.6051
R28967 por_dig_0.net7 por_dig_0.net7.n13 9.6005
R28968 por_dig_0.net7.n17 por_dig_0.net7.n0 9.47709
R28969 por_dig_0.net7.n23 por_dig_0.net7 9.3005
R28970 por_dig_0.net7.n23 por_dig_0.net7.n4 8.88939
R28971 por_dig_0.net7 por_dig_0.net7.n23 7.82272
R28972 por_dig_0.net7 por_dig_0.net7.n1 7.73474
R28973 por_dig_0.net7 por_dig_0.net7.n20 6.93567
R28974 por_dig_0.net7 por_dig_0.net7.n3 6.34564
R28975 por_dig_0.net7.n4 por_dig_0.net7 6.0165
R28976 por_dig_0.net7.n4 por_dig_0.net7 5.7605
R28977 por_dig_0.net7.n14 por_dig_0.net7 3.2005
R28978 por_dig_0.net7.n13 por_dig_0.net7 3.2005
R28979 por_dig_0.net7.n1 por_dig_0.net7 2.48634
R28980 por_dig_0.net7.n3 por_dig_0.net7 2.19479
R28981 por_dig_0.net7.n19 por_dig_0.net7 2.07109
R28982 por_dig_0.net7.n22 por_dig_0.net7 1.97868
R28983 por_dig_0.net7.n3 por_dig_0.net7 1.80756
R28984 por_dig_0.net7.n9 por_dig_0.net7 1.75534
R28985 por_ana_0.rstring_mux_0.vtrip5.n5 por_ana_0.rstring_mux_0.vtrip5.n3 50.7022
R28986 por_ana_0.rstring_mux_0.vtrip5.n2 por_ana_0.rstring_mux_0.vtrip5.n0 50.7022
R28987 por_ana_0.rstring_mux_0.vtrip5.n6 por_ana_0.rstring_mux_0.vtrip5.n2 14.7069
R28988 por_ana_0.rstring_mux_0.vtrip5.n5 por_ana_0.rstring_mux_0.vtrip5.n4 13.8791
R28989 por_ana_0.rstring_mux_0.vtrip5.n2 por_ana_0.rstring_mux_0.vtrip5.n1 13.8791
R28990 por_ana_0.rstring_mux_0.vtrip5.t0 por_ana_0.rstring_mux_0.vtrip5.n7 10.5857
R28991 por_ana_0.rstring_mux_0.vtrip5.n7 por_ana_0.rstring_mux_0.vtrip5.t1 10.5847
R28992 por_ana_0.rstring_mux_0.vtrip5.n3 por_ana_0.rstring_mux_0.vtrip5.t7 5.5395
R28993 por_ana_0.rstring_mux_0.vtrip5.n3 por_ana_0.rstring_mux_0.vtrip5.t6 5.5395
R28994 por_ana_0.rstring_mux_0.vtrip5.n0 por_ana_0.rstring_mux_0.vtrip5.t2 5.5395
R28995 por_ana_0.rstring_mux_0.vtrip5.n0 por_ana_0.rstring_mux_0.vtrip5.t3 5.5395
R28996 por_ana_0.rstring_mux_0.vtrip5.n7 por_ana_0.rstring_mux_0.vtrip5.n6 5.07153
R28997 por_ana_0.rstring_mux_0.vtrip5.n6 por_ana_0.rstring_mux_0.vtrip5.n5 3.33746
R28998 por_ana_0.rstring_mux_0.vtrip5.n4 por_ana_0.rstring_mux_0.vtrip5.t5 3.3065
R28999 por_ana_0.rstring_mux_0.vtrip5.n4 por_ana_0.rstring_mux_0.vtrip5.t4 3.3065
R29000 por_ana_0.rstring_mux_0.vtrip5.n1 por_ana_0.rstring_mux_0.vtrip5.t9 3.3065
R29001 por_ana_0.rstring_mux_0.vtrip5.n1 por_ana_0.rstring_mux_0.vtrip5.t8 3.3065
R29002 por_ana_0.rstring_mux_0.vtrip6.n5 por_ana_0.rstring_mux_0.vtrip6.n3 50.7022
R29003 por_ana_0.rstring_mux_0.vtrip6.n2 por_ana_0.rstring_mux_0.vtrip6.n0 50.7022
R29004 por_ana_0.rstring_mux_0.vtrip6.n7 por_ana_0.rstring_mux_0.vtrip6.n6 21.6754
R29005 por_ana_0.rstring_mux_0.vtrip6.n6 por_ana_0.rstring_mux_0.vtrip6.n5 14.944
R29006 por_ana_0.rstring_mux_0.vtrip6.n5 por_ana_0.rstring_mux_0.vtrip6.n4 13.8791
R29007 por_ana_0.rstring_mux_0.vtrip6.n2 por_ana_0.rstring_mux_0.vtrip6.n1 13.8791
R29008 por_ana_0.rstring_mux_0.vtrip6 por_ana_0.rstring_mux_0.vtrip6.t5 10.5739
R29009 por_ana_0.rstring_mux_0.vtrip6.n3 por_ana_0.rstring_mux_0.vtrip6.t4 5.5395
R29010 por_ana_0.rstring_mux_0.vtrip6.n3 por_ana_0.rstring_mux_0.vtrip6.t3 5.5395
R29011 por_ana_0.rstring_mux_0.vtrip6.n0 por_ana_0.rstring_mux_0.vtrip6.t9 5.5395
R29012 por_ana_0.rstring_mux_0.vtrip6.n0 por_ana_0.rstring_mux_0.vtrip6.t8 5.5395
R29013 por_ana_0.rstring_mux_0.vtrip6.n6 por_ana_0.rstring_mux_0.vtrip6.n2 5.01904
R29014 por_ana_0.rstring_mux_0.vtrip6.n4 por_ana_0.rstring_mux_0.vtrip6.t2 3.3065
R29015 por_ana_0.rstring_mux_0.vtrip6.n4 por_ana_0.rstring_mux_0.vtrip6.t1 3.3065
R29016 por_ana_0.rstring_mux_0.vtrip6.n1 por_ana_0.rstring_mux_0.vtrip6.t7 3.3065
R29017 por_ana_0.rstring_mux_0.vtrip6.n1 por_ana_0.rstring_mux_0.vtrip6.t6 3.3065
R29018 por_ana_0.rstring_mux_0.vtrip6.n7 por_ana_0.rstring_mux_0.vtrip6.t0 0.826075
R29019 por_ana_0.rstring_mux_0.vtrip6 por_ana_0.rstring_mux_0.vtrip6.n7 0.0563195
R29020 por_ana_0.schmitt_trigger_0.in.n3 por_ana_0.schmitt_trigger_0.in.t4 240.778
R29021 por_ana_0.schmitt_trigger_0.in.n0 por_ana_0.schmitt_trigger_0.in.t12 240.778
R29022 por_ana_0.schmitt_trigger_0.in.n3 por_ana_0.schmitt_trigger_0.in.t9 240.349
R29023 por_ana_0.schmitt_trigger_0.in.n2 por_ana_0.schmitt_trigger_0.in.t1 240.349
R29024 por_ana_0.schmitt_trigger_0.in.n1 por_ana_0.schmitt_trigger_0.in.t5 240.349
R29025 por_ana_0.schmitt_trigger_0.in.n0 por_ana_0.schmitt_trigger_0.in.t11 240.349
R29026 por_ana_0.schmitt_trigger_0.in.n12 por_ana_0.schmitt_trigger_0.in.t2 236.423
R29027 por_ana_0.schmitt_trigger_0.in.n12 por_ana_0.schmitt_trigger_0.in.t3 236.011
R29028 por_ana_0.schmitt_trigger_0.in.n10 por_ana_0.schmitt_trigger_0.in.n9 28.545
R29029 por_ana_0.schmitt_trigger_0.in.n11 por_ana_0.schmitt_trigger_0.in.n10 19.9248
R29030 por_ana_0.schmitt_trigger_0.in.n10 por_ana_0.schmitt_trigger_0.in.t0 5.93425
R29031 por_ana_0.schmitt_trigger_0.in por_ana_0.schmitt_trigger_0.in.n12 4.93075
R29032 por_ana_0.schmitt_trigger_0.in.n11 por_ana_0.schmitt_trigger_0.in.n4 4.72087
R29033 por_ana_0.schmitt_trigger_0.in.n1 por_ana_0.schmitt_trigger_0.in.n0 0.429848
R29034 por_ana_0.schmitt_trigger_0.in.n2 por_ana_0.schmitt_trigger_0.in.n1 0.429848
R29035 por_ana_0.schmitt_trigger_0.in.n4 por_ana_0.schmitt_trigger_0.in.n2 0.285826
R29036 por_ana_0.schmitt_trigger_0.in por_ana_0.schmitt_trigger_0.in.n11 0.216402
R29037 por_ana_0.schmitt_trigger_0.in.n4 por_ana_0.schmitt_trigger_0.in.n3 0.0956087
R29038 por_ana_0.schmitt_trigger_0.in.n5 por_ana_0.schmitt_trigger_0.in.t6 0.0791747
R29039 por_ana_0.schmitt_trigger_0.in.n6 por_ana_0.schmitt_trigger_0.in.n5 0.06865
R29040 por_ana_0.schmitt_trigger_0.in.n7 por_ana_0.schmitt_trigger_0.in.n6 0.06865
R29041 por_ana_0.schmitt_trigger_0.in.n8 por_ana_0.schmitt_trigger_0.in.n7 0.06865
R29042 por_ana_0.schmitt_trigger_0.in.n9 por_ana_0.schmitt_trigger_0.in.n8 0.06865
R29043 por_ana_0.schmitt_trigger_0.in.n5 por_ana_0.schmitt_trigger_0.in.t14 0.0110247
R29044 por_ana_0.schmitt_trigger_0.in.n6 por_ana_0.schmitt_trigger_0.in.t8 0.0110247
R29045 por_ana_0.schmitt_trigger_0.in.n7 por_ana_0.schmitt_trigger_0.in.t7 0.0110247
R29046 por_ana_0.schmitt_trigger_0.in.n8 por_ana_0.schmitt_trigger_0.in.t13 0.0110247
R29047 por_ana_0.schmitt_trigger_0.in.n9 por_ana_0.schmitt_trigger_0.in.t10 0.0110247
R29048 por_ana_0.schmitt_trigger_0.m.n5 por_ana_0.schmitt_trigger_0.m.t17 240.764
R29049 por_ana_0.schmitt_trigger_0.m.n6 por_ana_0.schmitt_trigger_0.m.t14 240.713
R29050 por_ana_0.schmitt_trigger_0.m.n7 por_ana_0.schmitt_trigger_0.m.t15 240.529
R29051 por_ana_0.schmitt_trigger_0.m.n5 por_ana_0.schmitt_trigger_0.m.t16 240.349
R29052 por_ana_0.schmitt_trigger_0.m.n10 por_ana_0.schmitt_trigger_0.m.n8 211.214
R29053 por_ana_0.schmitt_trigger_0.m.n2 por_ana_0.schmitt_trigger_0.m.n0 207.804
R29054 por_ana_0.schmitt_trigger_0.m.n2 por_ana_0.schmitt_trigger_0.m.n1 207.585
R29055 por_ana_0.schmitt_trigger_0.m.n4 por_ana_0.schmitt_trigger_0.m.n3 204.175
R29056 por_ana_0.schmitt_trigger_0.m.n10 por_ana_0.schmitt_trigger_0.m.n9 204.175
R29057 por_ana_0.schmitt_trigger_0.m.n13 por_ana_0.schmitt_trigger_0.m.n12 70.9014
R29058 por_ana_0.schmitt_trigger_0.m.n15 por_ana_0.schmitt_trigger_0.m.n14 70.9014
R29059 por_ana_0.schmitt_trigger_0.m.n8 por_ana_0.schmitt_trigger_0.m.t13 28.5655
R29060 por_ana_0.schmitt_trigger_0.m.n8 por_ana_0.schmitt_trigger_0.m.t11 28.5655
R29061 por_ana_0.schmitt_trigger_0.m.n3 por_ana_0.schmitt_trigger_0.m.t4 28.5655
R29062 por_ana_0.schmitt_trigger_0.m.n3 por_ana_0.schmitt_trigger_0.m.t6 28.5655
R29063 por_ana_0.schmitt_trigger_0.m.n1 por_ana_0.schmitt_trigger_0.m.t5 28.5655
R29064 por_ana_0.schmitt_trigger_0.m.n1 por_ana_0.schmitt_trigger_0.m.t7 28.5655
R29065 por_ana_0.schmitt_trigger_0.m.n0 por_ana_0.schmitt_trigger_0.m.t2 28.5655
R29066 por_ana_0.schmitt_trigger_0.m.n0 por_ana_0.schmitt_trigger_0.m.t3 28.5655
R29067 por_ana_0.schmitt_trigger_0.m.n9 por_ana_0.schmitt_trigger_0.m.t9 28.5655
R29068 por_ana_0.schmitt_trigger_0.m.n9 por_ana_0.schmitt_trigger_0.m.t8 28.5655
R29069 por_ana_0.schmitt_trigger_0.m.n12 por_ana_0.schmitt_trigger_0.m.t12 17.4005
R29070 por_ana_0.schmitt_trigger_0.m.n12 por_ana_0.schmitt_trigger_0.m.t10 17.4005
R29071 por_ana_0.schmitt_trigger_0.m.n14 por_ana_0.schmitt_trigger_0.m.t0 17.4005
R29072 por_ana_0.schmitt_trigger_0.m.n14 por_ana_0.schmitt_trigger_0.m.t1 17.4005
R29073 por_ana_0.schmitt_trigger_0.m.n7 por_ana_0.schmitt_trigger_0.m.n6 12.9318
R29074 por_ana_0.schmitt_trigger_0.m.n11 por_ana_0.schmitt_trigger_0.m.n10 8.3606
R29075 por_ana_0.schmitt_trigger_0.m.n4 por_ana_0.schmitt_trigger_0.m.n2 3.62811
R29076 por_ana_0.schmitt_trigger_0.m por_ana_0.schmitt_trigger_0.m.n4 0.819515
R29077 por_ana_0.schmitt_trigger_0.m por_ana_0.schmitt_trigger_0.m.n15 0.73133
R29078 por_ana_0.schmitt_trigger_0.m.n15 por_ana_0.schmitt_trigger_0.m.n13 0.688
R29079 por_ana_0.schmitt_trigger_0.m.n11 por_ana_0.schmitt_trigger_0.m.n7 0.358635
R29080 por_ana_0.schmitt_trigger_0.m.n13 por_ana_0.schmitt_trigger_0.m.n11 0.251558
R29081 por_ana_0.schmitt_trigger_0.m.n6 por_ana_0.schmitt_trigger_0.m.n5 0.0297969
R29082 por_ana_0.comparator_0.vnn.n7 por_ana_0.comparator_0.vnn.t14 244.34
R29083 por_ana_0.comparator_0.vnn.n7 por_ana_0.comparator_0.vnn.n20 204.284
R29084 por_ana_0.comparator_0.vnn.n7 por_ana_0.comparator_0.vnn.n21 204.284
R29085 por_ana_0.comparator_0.vnn.n7 por_ana_0.comparator_0.vnn.n22 204.284
R29086 por_ana_0.comparator_0.vnn.n7 por_ana_0.comparator_0.vnn.n23 204.284
R29087 por_ana_0.comparator_0.vnn.n7 por_ana_0.comparator_0.vnn.n25 204.284
R29088 por_ana_0.comparator_0.vnn.n7 por_ana_0.comparator_0.vnn.n26 204.284
R29089 por_ana_0.comparator_0.vnn.n7 por_ana_0.comparator_0.vnn.n24 204.284
R29090 por_ana_0.comparator_0.vnn.n6 por_ana_0.comparator_0.vnn.n17 199.784
R29091 por_ana_0.comparator_0.vnn.n6 por_ana_0.comparator_0.vnn.n16 199.65
R29092 por_ana_0.comparator_0.vnn.n6 por_ana_0.comparator_0.vnn.n18 199.65
R29093 por_ana_0.comparator_0.vnn.n6 por_ana_0.comparator_0.vnn.n19 199.65
R29094 por_ana_0.comparator_0.vnn.n0 por_ana_0.comparator_0.vnn.n8 71.9371
R29095 por_ana_0.comparator_0.vnn.n0 por_ana_0.comparator_0.vnn.n15 70.9612
R29096 por_ana_0.comparator_0.vnn.n0 por_ana_0.comparator_0.vnn.n14 70.9612
R29097 por_ana_0.comparator_0.vnn.n0 por_ana_0.comparator_0.vnn.n13 70.9612
R29098 por_ana_0.comparator_0.vnn.n0 por_ana_0.comparator_0.vnn.n12 70.9612
R29099 por_ana_0.comparator_0.vnn.n0 por_ana_0.comparator_0.vnn.n11 70.9612
R29100 por_ana_0.comparator_0.vnn.n0 por_ana_0.comparator_0.vnn.n10 70.9612
R29101 por_ana_0.comparator_0.vnn.n0 por_ana_0.comparator_0.vnn.n9 70.9612
R29102 por_ana_0.comparator_0.vnn.n20 por_ana_0.comparator_0.vnn.t2 27.6955
R29103 por_ana_0.comparator_0.vnn.n20 por_ana_0.comparator_0.vnn.t4 27.6955
R29104 por_ana_0.comparator_0.vnn.n21 por_ana_0.comparator_0.vnn.t12 27.6955
R29105 por_ana_0.comparator_0.vnn.n21 por_ana_0.comparator_0.vnn.t1 27.6955
R29106 por_ana_0.comparator_0.vnn.n22 por_ana_0.comparator_0.vnn.t0 27.6955
R29107 por_ana_0.comparator_0.vnn.n22 por_ana_0.comparator_0.vnn.t3 27.6955
R29108 por_ana_0.comparator_0.vnn.n23 por_ana_0.comparator_0.vnn.t9 27.6955
R29109 por_ana_0.comparator_0.vnn.n23 por_ana_0.comparator_0.vnn.t10 27.6955
R29110 por_ana_0.comparator_0.vnn.n25 por_ana_0.comparator_0.vnn.t8 27.6955
R29111 por_ana_0.comparator_0.vnn.n25 por_ana_0.comparator_0.vnn.t7 27.6955
R29112 por_ana_0.comparator_0.vnn.n26 por_ana_0.comparator_0.vnn.t6 27.6955
R29113 por_ana_0.comparator_0.vnn.n26 por_ana_0.comparator_0.vnn.t5 27.6955
R29114 por_ana_0.comparator_0.vnn.n17 por_ana_0.comparator_0.vnn.t44 27.6955
R29115 por_ana_0.comparator_0.vnn.n17 por_ana_0.comparator_0.vnn.t46 27.6955
R29116 por_ana_0.comparator_0.vnn.n16 por_ana_0.comparator_0.vnn.t38 27.6955
R29117 por_ana_0.comparator_0.vnn.n16 por_ana_0.comparator_0.vnn.t42 27.6955
R29118 por_ana_0.comparator_0.vnn.n18 por_ana_0.comparator_0.vnn.t36 27.6955
R29119 por_ana_0.comparator_0.vnn.n18 por_ana_0.comparator_0.vnn.t40 27.6955
R29120 por_ana_0.comparator_0.vnn.n19 por_ana_0.comparator_0.vnn.t32 27.6955
R29121 por_ana_0.comparator_0.vnn.n19 por_ana_0.comparator_0.vnn.t34 27.6955
R29122 por_ana_0.comparator_0.vnn.n24 por_ana_0.comparator_0.vnn.t11 27.6955
R29123 por_ana_0.comparator_0.vnn.n24 por_ana_0.comparator_0.vnn.t13 27.6955
R29124 por_ana_0.comparator_0.vnn.n15 por_ana_0.comparator_0.vnn.t19 16.5305
R29125 por_ana_0.comparator_0.vnn.n15 por_ana_0.comparator_0.vnn.t23 16.5305
R29126 por_ana_0.comparator_0.vnn.n14 por_ana_0.comparator_0.vnn.t22 16.5305
R29127 por_ana_0.comparator_0.vnn.n14 por_ana_0.comparator_0.vnn.t28 16.5305
R29128 por_ana_0.comparator_0.vnn.n13 por_ana_0.comparator_0.vnn.t16 16.5305
R29129 por_ana_0.comparator_0.vnn.n13 por_ana_0.comparator_0.vnn.t26 16.5305
R29130 por_ana_0.comparator_0.vnn.n12 por_ana_0.comparator_0.vnn.t18 16.5305
R29131 por_ana_0.comparator_0.vnn.n12 por_ana_0.comparator_0.vnn.t24 16.5305
R29132 por_ana_0.comparator_0.vnn.n11 por_ana_0.comparator_0.vnn.t21 16.5305
R29133 por_ana_0.comparator_0.vnn.n11 por_ana_0.comparator_0.vnn.t29 16.5305
R29134 por_ana_0.comparator_0.vnn.n10 por_ana_0.comparator_0.vnn.t17 16.5305
R29135 por_ana_0.comparator_0.vnn.n10 por_ana_0.comparator_0.vnn.t25 16.5305
R29136 por_ana_0.comparator_0.vnn.n9 por_ana_0.comparator_0.vnn.t20 16.5305
R29137 por_ana_0.comparator_0.vnn.n9 por_ana_0.comparator_0.vnn.t30 16.5305
R29138 por_ana_0.comparator_0.vnn.n8 por_ana_0.comparator_0.vnn.t15 16.5305
R29139 por_ana_0.comparator_0.vnn.n8 por_ana_0.comparator_0.vnn.t27 16.5305
R29140 por_ana_0.comparator_0.vnn.n1 por_ana_0.comparator_0.vnn.t54 16.4779
R29141 por_ana_0.comparator_0.vnn.n3 por_ana_0.comparator_0.vnn.t56 16.4779
R29142 por_ana_0.comparator_0.vnn.n4 por_ana_0.comparator_0.vnn.t55 16.4779
R29143 por_ana_0.comparator_0.vnn.n2 por_ana_0.comparator_0.vnn.t62 16.4779
R29144 por_ana_0.comparator_0.vnn.n1 por_ana_0.comparator_0.vnn.t57 16.4779
R29145 por_ana_0.comparator_0.vnn.n1 por_ana_0.comparator_0.vnn.t51 16.4779
R29146 por_ana_0.comparator_0.vnn.n1 por_ana_0.comparator_0.vnn.t52 16.4779
R29147 por_ana_0.comparator_0.vnn.n5 por_ana_0.comparator_0.vnn.t61 16.4779
R29148 por_ana_0.comparator_0.vnn.n6 por_ana_0.comparator_0.vnn.t33 14.2251
R29149 por_ana_0.comparator_0.vnn.n6 por_ana_0.comparator_0.vnn.t31 14.2251
R29150 por_ana_0.comparator_0.vnn.n6 por_ana_0.comparator_0.vnn.t39 14.2251
R29151 por_ana_0.comparator_0.vnn.n6 por_ana_0.comparator_0.vnn.t35 14.2251
R29152 por_ana_0.comparator_0.vnn.n6 por_ana_0.comparator_0.vnn.t41 14.2251
R29153 por_ana_0.comparator_0.vnn.n6 por_ana_0.comparator_0.vnn.t37 14.2251
R29154 por_ana_0.comparator_0.vnn.n6 por_ana_0.comparator_0.vnn.t43 14.2251
R29155 por_ana_0.comparator_0.vnn.n6 por_ana_0.comparator_0.vnn.t45 14.2251
R29156 por_ana_0.comparator_0.vnn por_ana_0.comparator_0.vnn.n1 13.4051
R29157 por_ana_0.comparator_0.vnn por_ana_0.comparator_0.vnn.n0 11.9816
R29158 por_ana_0.comparator_0.vnn.n1 por_ana_0.comparator_0.vnn.t48 11.9724
R29159 por_ana_0.comparator_0.vnn.n3 por_ana_0.comparator_0.vnn.t50 11.9724
R29160 por_ana_0.comparator_0.vnn.n4 por_ana_0.comparator_0.vnn.t49 11.9724
R29161 por_ana_0.comparator_0.vnn.n2 por_ana_0.comparator_0.vnn.t58 11.9724
R29162 por_ana_0.comparator_0.vnn.n1 por_ana_0.comparator_0.vnn.t53 11.9724
R29163 por_ana_0.comparator_0.vnn.n1 por_ana_0.comparator_0.vnn.t59 11.9724
R29164 por_ana_0.comparator_0.vnn.n1 por_ana_0.comparator_0.vnn.t60 11.9724
R29165 por_ana_0.comparator_0.vnn.n5 por_ana_0.comparator_0.vnn.t47 11.9724
R29166 por_ana_0.comparator_0.vnn por_ana_0.comparator_0.vnn.n7 9.57847
R29167 por_ana_0.comparator_0.vnn.n1 por_ana_0.comparator_0.vnn.n4 9.23963
R29168 por_ana_0.comparator_0.vnn.n1 por_ana_0.comparator_0.vnn.n3 9.23963
R29169 por_ana_0.comparator_0.vnn.n1 por_ana_0.comparator_0.vnn.n2 9.23963
R29170 por_ana_0.comparator_0.vnn.n1 por_ana_0.comparator_0.vnn.n5 9.22553
R29171 por_ana_0.comparator_0.vnn.n7 por_ana_0.comparator_0.vnn.n6 8.84171
R29172 por_ana_0.comparator_0.vinn.n6 por_ana_0.comparator_0.vinn.t27 51.0275
R29173 por_ana_0.comparator_0.vinn.n0 por_ana_0.comparator_0.vinn.n17 48.371
R29174 por_ana_0.comparator_0.vinn.n1 por_ana_0.comparator_0.vinn.n20 48.371
R29175 por_ana_0.comparator_0.vinn.n2 por_ana_0.comparator_0.vinn.n23 48.371
R29176 por_ana_0.comparator_0.vinn.n3 por_ana_0.comparator_0.vinn.n26 48.371
R29177 por_ana_0.comparator_0.vinn.n29 por_ana_0.comparator_0.vinn.n4 48.371
R29178 por_ana_0.comparator_0.vinn.n5 por_ana_0.comparator_0.vinn.n9 48.371
R29179 por_ana_0.comparator_0.vinn.n6 por_ana_0.comparator_0.vinn.n11 48.371
R29180 por_ana_0.comparator_0.vinn.n7 por_ana_0.comparator_0.vinn.n14 48.371
R29181 por_ana_0.comparator_0.vinn.n10 por_ana_0.comparator_0.vinn.n7 45.4885
R29182 por_ana_0.comparator_0.vinn.n13 por_ana_0.comparator_0.vinn.n0 45.4885
R29183 por_ana_0.comparator_0.vinn.n16 por_ana_0.comparator_0.vinn.n1 45.4885
R29184 por_ana_0.comparator_0.vinn.n19 por_ana_0.comparator_0.vinn.n2 45.4885
R29185 por_ana_0.comparator_0.vinn.n22 por_ana_0.comparator_0.vinn.n3 45.4885
R29186 por_ana_0.comparator_0.vinn.n25 por_ana_0.comparator_0.vinn.n4 45.4885
R29187 por_ana_0.comparator_0.vinn.n5 por_ana_0.comparator_0.vinn.n30 45.4885
R29188 por_ana_0.comparator_0.vinn.n47 por_ana_0.comparator_0.vinn.n46 45.3881
R29189 por_ana_0.comparator_0.vinn.n12 por_ana_0.comparator_0.vinn.t46 20.2802
R29190 por_ana_0.comparator_0.vinn.n66 por_ana_0.comparator_0.vinn.n65 17.7666
R29191 por_ana_0.comparator_0.vinn.n63 por_ana_0.comparator_0.vinn.n62 17.7666
R29192 por_ana_0.comparator_0.vinn.n60 por_ana_0.comparator_0.vinn.n59 17.7666
R29193 por_ana_0.comparator_0.vinn.n57 por_ana_0.comparator_0.vinn.n56 17.7666
R29194 por_ana_0.comparator_0.vinn.n54 por_ana_0.comparator_0.vinn.n53 17.7666
R29195 por_ana_0.comparator_0.vinn.n51 por_ana_0.comparator_0.vinn.n50 17.7666
R29196 por_ana_0.comparator_0.vinn.n12 por_ana_0.comparator_0.vinn.n8 17.7666
R29197 por_ana_0.comparator_0.vinn.n47 por_ana_0.comparator_0.vinn.n31 17.6963
R29198 por_ana_0.comparator_0.vinn.n64 por_ana_0.comparator_0.vinn.n63 16.9742
R29199 por_ana_0.comparator_0.vinn.n61 por_ana_0.comparator_0.vinn.n60 16.9742
R29200 por_ana_0.comparator_0.vinn.n58 por_ana_0.comparator_0.vinn.n57 16.9742
R29201 por_ana_0.comparator_0.vinn.n55 por_ana_0.comparator_0.vinn.n54 16.9742
R29202 por_ana_0.comparator_0.vinn.n52 por_ana_0.comparator_0.vinn.n51 16.9742
R29203 por_ana_0.comparator_0.vinn.n49 por_ana_0.comparator_0.vinn.n48 16.9742
R29204 por_ana_0.comparator_0.vinn.n67 por_ana_0.comparator_0.vinn.n66 16.9742
R29205 por_ana_0.comparator_0.vinn.n39 por_ana_0.comparator_0.vinn.t57 9.72783
R29206 por_ana_0.comparator_0.vinn.n32 por_ana_0.comparator_0.vinn.t49 9.65028
R29207 por_ana_0.comparator_0.vinn.n46 por_ana_0.comparator_0.vinn.n38 8.96563
R29208 por_ana_0.comparator_0.vinn.n45 por_ana_0.comparator_0.vinn.t50 8.73727
R29209 por_ana_0.comparator_0.vinn.n44 por_ana_0.comparator_0.vinn.t58 8.73727
R29210 por_ana_0.comparator_0.vinn.n43 por_ana_0.comparator_0.vinn.t56 8.73727
R29211 por_ana_0.comparator_0.vinn.n42 por_ana_0.comparator_0.vinn.t51 8.73727
R29212 por_ana_0.comparator_0.vinn.n41 por_ana_0.comparator_0.vinn.t60 8.73727
R29213 por_ana_0.comparator_0.vinn.n40 por_ana_0.comparator_0.vinn.t52 8.73727
R29214 por_ana_0.comparator_0.vinn.n39 por_ana_0.comparator_0.vinn.t61 8.73727
R29215 por_ana_0.comparator_0.vinn.n38 por_ana_0.comparator_0.vinn.t59 8.65985
R29216 por_ana_0.comparator_0.vinn.n37 por_ana_0.comparator_0.vinn.t53 8.65985
R29217 por_ana_0.comparator_0.vinn.n36 por_ana_0.comparator_0.vinn.t48 8.65985
R29218 por_ana_0.comparator_0.vinn.n35 por_ana_0.comparator_0.vinn.t62 8.65985
R29219 por_ana_0.comparator_0.vinn.n34 por_ana_0.comparator_0.vinn.t54 8.65985
R29220 por_ana_0.comparator_0.vinn.n33 por_ana_0.comparator_0.vinn.t63 8.65985
R29221 por_ana_0.comparator_0.vinn.n32 por_ana_0.comparator_0.vinn.t55 8.65985
R29222 por_ana_0.comparator_0.vinn.n46 por_ana_0.comparator_0.vinn.n45 5.98511
R29223 por_ana_0.comparator_0.vinn.t6 por_ana_0.comparator_0.vinn.n10 5.5395
R29224 por_ana_0.comparator_0.vinn.n10 por_ana_0.comparator_0.vinn.t41 5.5395
R29225 por_ana_0.comparator_0.vinn.t1 por_ana_0.comparator_0.vinn.n13 5.5395
R29226 por_ana_0.comparator_0.vinn.n13 por_ana_0.comparator_0.vinn.t28 5.5395
R29227 por_ana_0.comparator_0.vinn.n17 por_ana_0.comparator_0.vinn.t29 5.5395
R29228 por_ana_0.comparator_0.vinn.n17 por_ana_0.comparator_0.vinn.t0 5.5395
R29229 por_ana_0.comparator_0.vinn.t0 por_ana_0.comparator_0.vinn.n16 5.5395
R29230 por_ana_0.comparator_0.vinn.n16 por_ana_0.comparator_0.vinn.t33 5.5395
R29231 por_ana_0.comparator_0.vinn.n20 por_ana_0.comparator_0.vinn.t32 5.5395
R29232 por_ana_0.comparator_0.vinn.n20 por_ana_0.comparator_0.vinn.t2 5.5395
R29233 por_ana_0.comparator_0.vinn.t2 por_ana_0.comparator_0.vinn.n19 5.5395
R29234 por_ana_0.comparator_0.vinn.n19 por_ana_0.comparator_0.vinn.t11 5.5395
R29235 por_ana_0.comparator_0.vinn.n23 por_ana_0.comparator_0.vinn.t10 5.5395
R29236 por_ana_0.comparator_0.vinn.n23 por_ana_0.comparator_0.vinn.t5 5.5395
R29237 por_ana_0.comparator_0.vinn.t5 por_ana_0.comparator_0.vinn.n22 5.5395
R29238 por_ana_0.comparator_0.vinn.n22 por_ana_0.comparator_0.vinn.t45 5.5395
R29239 por_ana_0.comparator_0.vinn.n26 por_ana_0.comparator_0.vinn.t44 5.5395
R29240 por_ana_0.comparator_0.vinn.n26 por_ana_0.comparator_0.vinn.t4 5.5395
R29241 por_ana_0.comparator_0.vinn.t4 por_ana_0.comparator_0.vinn.n25 5.5395
R29242 por_ana_0.comparator_0.vinn.n25 por_ana_0.comparator_0.vinn.t31 5.5395
R29243 por_ana_0.comparator_0.vinn.n29 por_ana_0.comparator_0.vinn.t30 5.5395
R29244 por_ana_0.comparator_0.vinn.t3 por_ana_0.comparator_0.vinn.n29 5.5395
R29245 por_ana_0.comparator_0.vinn.n30 por_ana_0.comparator_0.vinn.t3 5.5395
R29246 por_ana_0.comparator_0.vinn.n30 por_ana_0.comparator_0.vinn.t25 5.5395
R29247 por_ana_0.comparator_0.vinn.n9 por_ana_0.comparator_0.vinn.t24 5.5395
R29248 por_ana_0.comparator_0.vinn.n9 por_ana_0.comparator_0.vinn.t7 5.5395
R29249 por_ana_0.comparator_0.vinn.n11 por_ana_0.comparator_0.vinn.t26 5.5395
R29250 por_ana_0.comparator_0.vinn.n11 por_ana_0.comparator_0.vinn.t6 5.5395
R29251 por_ana_0.comparator_0.vinn.n14 por_ana_0.comparator_0.vinn.t40 5.5395
R29252 por_ana_0.comparator_0.vinn.n14 por_ana_0.comparator_0.vinn.t1 5.5395
R29253 por_ana_0.comparator_0.vinn.n28 por_ana_0.comparator_0.vinn.n5 3.79433
R29254 por_ana_0.comparator_0.vinn.n15 por_ana_0.comparator_0.vinn.n6 3.79433
R29255 por_ana_0.comparator_0.vinn.n4 por_ana_0.comparator_0.vinn.n28 3.4105
R29256 por_ana_0.comparator_0.vinn.n27 por_ana_0.comparator_0.vinn.n3 3.4105
R29257 por_ana_0.comparator_0.vinn.n24 por_ana_0.comparator_0.vinn.n2 3.4105
R29258 por_ana_0.comparator_0.vinn.n21 por_ana_0.comparator_0.vinn.n1 3.4105
R29259 por_ana_0.comparator_0.vinn.n18 por_ana_0.comparator_0.vinn.n0 3.4105
R29260 por_ana_0.comparator_0.vinn.n15 por_ana_0.comparator_0.vinn.n7 3.4105
R29261 por_ana_0.comparator_0.vinn.n65 por_ana_0.comparator_0.vinn.t20 3.3065
R29262 por_ana_0.comparator_0.vinn.n65 por_ana_0.comparator_0.vinn.t13 3.3065
R29263 por_ana_0.comparator_0.vinn.t13 por_ana_0.comparator_0.vinn.n64 3.3065
R29264 por_ana_0.comparator_0.vinn.n64 por_ana_0.comparator_0.vinn.t37 3.3065
R29265 por_ana_0.comparator_0.vinn.n62 por_ana_0.comparator_0.vinn.t36 3.3065
R29266 por_ana_0.comparator_0.vinn.n62 por_ana_0.comparator_0.vinn.t12 3.3065
R29267 por_ana_0.comparator_0.vinn.t12 por_ana_0.comparator_0.vinn.n61 3.3065
R29268 por_ana_0.comparator_0.vinn.n61 por_ana_0.comparator_0.vinn.t42 3.3065
R29269 por_ana_0.comparator_0.vinn.n59 por_ana_0.comparator_0.vinn.t43 3.3065
R29270 por_ana_0.comparator_0.vinn.n59 por_ana_0.comparator_0.vinn.t14 3.3065
R29271 por_ana_0.comparator_0.vinn.t14 por_ana_0.comparator_0.vinn.n58 3.3065
R29272 por_ana_0.comparator_0.vinn.n58 por_ana_0.comparator_0.vinn.t9 3.3065
R29273 por_ana_0.comparator_0.vinn.n56 por_ana_0.comparator_0.vinn.t8 3.3065
R29274 por_ana_0.comparator_0.vinn.n56 por_ana_0.comparator_0.vinn.t17 3.3065
R29275 por_ana_0.comparator_0.vinn.t17 por_ana_0.comparator_0.vinn.n55 3.3065
R29276 por_ana_0.comparator_0.vinn.n55 por_ana_0.comparator_0.vinn.t35 3.3065
R29277 por_ana_0.comparator_0.vinn.n53 por_ana_0.comparator_0.vinn.t34 3.3065
R29278 por_ana_0.comparator_0.vinn.n53 por_ana_0.comparator_0.vinn.t16 3.3065
R29279 por_ana_0.comparator_0.vinn.t16 por_ana_0.comparator_0.vinn.n52 3.3065
R29280 por_ana_0.comparator_0.vinn.n52 por_ana_0.comparator_0.vinn.t39 3.3065
R29281 por_ana_0.comparator_0.vinn.n50 por_ana_0.comparator_0.vinn.t38 3.3065
R29282 por_ana_0.comparator_0.vinn.n50 por_ana_0.comparator_0.vinn.t15 3.3065
R29283 por_ana_0.comparator_0.vinn.t15 por_ana_0.comparator_0.vinn.n49 3.3065
R29284 por_ana_0.comparator_0.vinn.n49 por_ana_0.comparator_0.vinn.t23 3.3065
R29285 por_ana_0.comparator_0.vinn.n31 por_ana_0.comparator_0.vinn.t22 3.3065
R29286 por_ana_0.comparator_0.vinn.n31 por_ana_0.comparator_0.vinn.t19 3.3065
R29287 por_ana_0.comparator_0.vinn.n8 por_ana_0.comparator_0.vinn.t47 3.3065
R29288 por_ana_0.comparator_0.vinn.t18 por_ana_0.comparator_0.vinn.n8 3.3065
R29289 por_ana_0.comparator_0.vinn.t18 por_ana_0.comparator_0.vinn.n67 3.3065
R29290 por_ana_0.comparator_0.vinn.n67 por_ana_0.comparator_0.vinn.t21 3.3065
R29291 por_ana_0.comparator_0.vinn.n66 por_ana_0.comparator_0.vinn.n7 1.98488
R29292 por_ana_0.comparator_0.vinn.n6 por_ana_0.comparator_0.vinn.n12 1.98488
R29293 por_ana_0.comparator_0.vinn.n48 por_ana_0.comparator_0.vinn.n5 1.98488
R29294 por_ana_0.comparator_0.vinn.n51 por_ana_0.comparator_0.vinn.n4 1.98488
R29295 por_ana_0.comparator_0.vinn.n54 por_ana_0.comparator_0.vinn.n3 1.98488
R29296 por_ana_0.comparator_0.vinn.n57 por_ana_0.comparator_0.vinn.n2 1.98488
R29297 por_ana_0.comparator_0.vinn.n60 por_ana_0.comparator_0.vinn.n1 1.98488
R29298 por_ana_0.comparator_0.vinn.n63 por_ana_0.comparator_0.vinn.n0 1.98488
R29299 por_ana_0.comparator_0.vinn.n45 por_ana_0.comparator_0.vinn.n44 0.99106
R29300 por_ana_0.comparator_0.vinn.n44 por_ana_0.comparator_0.vinn.n43 0.99106
R29301 por_ana_0.comparator_0.vinn.n43 por_ana_0.comparator_0.vinn.n42 0.99106
R29302 por_ana_0.comparator_0.vinn.n42 por_ana_0.comparator_0.vinn.n41 0.99106
R29303 por_ana_0.comparator_0.vinn.n41 por_ana_0.comparator_0.vinn.n40 0.99106
R29304 por_ana_0.comparator_0.vinn.n40 por_ana_0.comparator_0.vinn.n39 0.99106
R29305 por_ana_0.comparator_0.vinn.n38 por_ana_0.comparator_0.vinn.n37 0.99093
R29306 por_ana_0.comparator_0.vinn.n37 por_ana_0.comparator_0.vinn.n36 0.99093
R29307 por_ana_0.comparator_0.vinn.n36 por_ana_0.comparator_0.vinn.n35 0.99093
R29308 por_ana_0.comparator_0.vinn.n35 por_ana_0.comparator_0.vinn.n34 0.99093
R29309 por_ana_0.comparator_0.vinn.n34 por_ana_0.comparator_0.vinn.n33 0.99093
R29310 por_ana_0.comparator_0.vinn.n33 por_ana_0.comparator_0.vinn.n32 0.99093
R29311 por_ana_0.comparator_0.vinn.n28 por_ana_0.comparator_0.vinn.n27 0.384333
R29312 por_ana_0.comparator_0.vinn.n27 por_ana_0.comparator_0.vinn.n24 0.384333
R29313 por_ana_0.comparator_0.vinn.n24 por_ana_0.comparator_0.vinn.n21 0.384333
R29314 por_ana_0.comparator_0.vinn.n21 por_ana_0.comparator_0.vinn.n18 0.384333
R29315 por_ana_0.comparator_0.vinn.n18 por_ana_0.comparator_0.vinn.n15 0.384333
R29316 por_ana_0.comparator_0.vinn.n48 por_ana_0.comparator_0.vinn.n47 0.0708125
R29317 por_dig_0.cnt_por\[0\] por_dig_0.cnt_por\[0\].n10 439.457
R29318 por_dig_0.cnt_por\[0\].t22 por_dig_0.cnt_por\[0\].t13 395.01
R29319 por_dig_0.cnt_por\[0\].n17 por_dig_0.cnt_por\[0\].t11 334.723
R29320 por_dig_0.cnt_por\[0\].n11 por_dig_0.cnt_por\[0\].t24 329.902
R29321 por_dig_0.cnt_por\[0\] por_dig_0.cnt_por\[0\].t22 320.745
R29322 por_dig_0.cnt_por\[0\].n10 por_dig_0.cnt_por\[0\].t14 272.062
R29323 por_dig_0.cnt_por\[0\].n2 por_dig_0.cnt_por\[0\].n1 248.085
R29324 por_dig_0.cnt_por\[0\].n25 por_dig_0.cnt_por\[0\].t26 241.536
R29325 por_dig_0.cnt_por\[0\].n22 por_dig_0.cnt_por\[0\].t18 241.536
R29326 por_dig_0.cnt_por\[0\].n15 por_dig_0.cnt_por\[0\].t25 241.536
R29327 por_dig_0.cnt_por\[0\].n8 por_dig_0.cnt_por\[0\].t20 241.536
R29328 por_dig_0.cnt_por\[0\].n3 por_dig_0.cnt_por\[0\].t23 237.787
R29329 por_dig_0.cnt_por\[0\].n5 por_dig_0.cnt_por\[0\].t19 221.72
R29330 por_dig_0.cnt_por\[0\].n2 por_dig_0.cnt_por\[0\].n0 208.507
R29331 por_dig_0.cnt_por\[0\].n17 por_dig_0.cnt_por\[0\].t16 206.19
R29332 por_dig_0.cnt_por\[0\].n10 por_dig_0.cnt_por\[0\].t21 206.19
R29333 por_dig_0.cnt_por\[0\].n6 por_dig_0.cnt_por\[0\].t12 192.264
R29334 por_dig_0.cnt_por\[0\].n16 por_dig_0.cnt_por\[0\].n15 190.109
R29335 por_dig_0.cnt_por\[0\].n9 por_dig_0.cnt_por\[0\].n8 180.948
R29336 por_dig_0.cnt_por\[0\].n25 por_dig_0.cnt_por\[0\].t15 169.237
R29337 por_dig_0.cnt_por\[0\].n22 por_dig_0.cnt_por\[0\].t27 169.237
R29338 por_dig_0.cnt_por\[0\].n15 por_dig_0.cnt_por\[0\].t9 169.237
R29339 por_dig_0.cnt_por\[0\].n8 por_dig_0.cnt_por\[0\].t8 169.237
R29340 por_dig_0.cnt_por\[0\].n23 por_dig_0.cnt_por\[0\].n22 159.952
R29341 por_dig_0.cnt_por\[0\] por_dig_0.cnt_por\[0\].n25 157.166
R29342 por_dig_0.cnt_por\[0\].n3 por_dig_0.cnt_por\[0\] 155.201
R29343 por_dig_0.cnt_por\[0\].n18 por_dig_0.cnt_por\[0\].n17 152
R29344 por_dig_0.cnt_por\[0\].n12 por_dig_0.cnt_por\[0\].n11 152
R29345 por_dig_0.cnt_por\[0\].n7 por_dig_0.cnt_por\[0\].n6 152
R29346 por_dig_0.cnt_por\[0\].n4 por_dig_0.cnt_por\[0\].t10 149.421
R29347 por_dig_0.cnt_por\[0\].n11 por_dig_0.cnt_por\[0\].t17 148.35
R29348 por_dig_0.cnt_por\[0\].n33 por_dig_0.cnt_por\[0\].n31 137.576
R29349 por_dig_0.cnt_por\[0\].n33 por_dig_0.cnt_por\[0\].n32 99.1759
R29350 por_dig_0.cnt_por\[0\].n4 por_dig_0.cnt_por\[0\].n3 55.3412
R29351 por_dig_0.cnt_por\[0\].n6 por_dig_0.cnt_por\[0\].n5 28.5635
R29352 por_dig_0.cnt_por\[0\].n7 por_dig_0.cnt_por\[0\] 28.1605
R29353 por_dig_0.cnt_por\[0\].n14 por_dig_0.cnt_por\[0\].n9 27.1384
R29354 por_dig_0.cnt_por\[0\].n0 por_dig_0.cnt_por\[0\].t4 26.5955
R29355 por_dig_0.cnt_por\[0\].n0 por_dig_0.cnt_por\[0\].t6 26.5955
R29356 por_dig_0.cnt_por\[0\].n1 por_dig_0.cnt_por\[0\].t5 26.5955
R29357 por_dig_0.cnt_por\[0\].n1 por_dig_0.cnt_por\[0\].t7 26.5955
R29358 por_dig_0.cnt_por\[0\].n19 por_dig_0.cnt_por\[0\] 26.1855
R29359 por_dig_0.cnt_por\[0\].n31 por_dig_0.cnt_por\[0\].t2 24.9236
R29360 por_dig_0.cnt_por\[0\].n31 por_dig_0.cnt_por\[0\].t0 24.9236
R29361 por_dig_0.cnt_por\[0\].n32 por_dig_0.cnt_por\[0\].t1 24.9236
R29362 por_dig_0.cnt_por\[0\].n32 por_dig_0.cnt_por\[0\].t3 24.9236
R29363 por_dig_0.cnt_por\[0\] por_dig_0.cnt_por\[0\].n33 22.8275
R29364 por_dig_0.cnt_por\[0\].n12 por_dig_0.cnt_por\[0\] 20.211
R29365 por_dig_0.cnt_por\[0\].n30 por_dig_0.cnt_por\[0\].n2 17.2539
R29366 por_dig_0.cnt_por\[0\].n30 por_dig_0.cnt_por\[0\].n29 16.5768
R29367 por_dig_0.cnt_por\[0\].n28 por_dig_0.cnt_por\[0\].n24 16.0972
R29368 por_dig_0.cnt_por\[0\].n21 por_dig_0.cnt_por\[0\] 15.364
R29369 por_dig_0.cnt_por\[0\].n16 por_dig_0.cnt_por\[0\] 14.8762
R29370 por_dig_0.cnt_por\[0\].n24 por_dig_0.cnt_por\[0\] 14.1918
R29371 por_dig_0.cnt_por\[0\].n27 por_dig_0.cnt_por\[0\].n26 13.734
R29372 por_dig_0.cnt_por\[0\] por_dig_0.cnt_por\[0\].n23 12.8005
R29373 por_dig_0.cnt_por\[0\].n27 por_dig_0.cnt_por\[0\] 12.5005
R29374 por_dig_0.cnt_por\[0\].n26 por_dig_0.cnt_por\[0\] 11.4531
R29375 por_dig_0.cnt_por\[0\].n21 por_dig_0.cnt_por\[0\].n20 11.1694
R29376 por_dig_0.cnt_por\[0\].n19 por_dig_0.cnt_por\[0\].n18 10.3976
R29377 por_dig_0.cnt_por\[0\].n14 por_dig_0.cnt_por\[0\].n13 9.3005
R29378 por_dig_0.cnt_por\[0\].n18 por_dig_0.cnt_por\[0\] 8.22907
R29379 por_dig_0.cnt_por\[0\].n13 por_dig_0.cnt_por\[0\] 6.06366
R29380 por_dig_0.cnt_por\[0\].n29 por_dig_0.cnt_por\[0\].n28 5.88649
R29381 por_dig_0.cnt_por\[0\].n28 por_dig_0.cnt_por\[0\].n27 4.79462
R29382 por_dig_0.cnt_por\[0\].n24 por_dig_0.cnt_por\[0\] 4.73093
R29383 por_dig_0.cnt_por\[0\].n13 por_dig_0.cnt_por\[0\].n12 4.71629
R29384 por_dig_0.cnt_por\[0\].n26 por_dig_0.cnt_por\[0\] 3.81804
R29385 por_dig_0.cnt_por\[0\].n5 por_dig_0.cnt_por\[0\].n4 3.57087
R29386 por_dig_0.cnt_por\[0\].n23 por_dig_0.cnt_por\[0\] 3.29747
R29387 por_dig_0.cnt_por\[0\].n9 por_dig_0.cnt_por\[0\] 3.10907
R29388 por_dig_0.cnt_por\[0\] por_dig_0.cnt_por\[0\].n30 2.65416
R29389 por_dig_0.cnt_por\[0\].n29 por_dig_0.cnt_por\[0\].n21 2.33292
R29390 por_dig_0.cnt_por\[0\] por_dig_0.cnt_por\[0\].n16 1.73023
R29391 por_dig_0.cnt_por\[0\] por_dig_0.cnt_por\[0\].n7 1.2805
R29392 por_dig_0.cnt_por\[0\].n20 por_dig_0.cnt_por\[0\] 1.02729
R29393 por_dig_0.cnt_por\[0\] por_dig_0.cnt_por\[0\].n19 0.976626
R29394 por_dig_0.cnt_por\[0\].n20 por_dig_0.cnt_por\[0\].n14 0.960321
R29395 pwup_filt.n15 pwup_filt.t33 260.322
R29396 pwup_filt.n2 pwup_filt.n0 243.458
R29397 pwup_filt.n2 pwup_filt.n1 205.059
R29398 pwup_filt.n4 pwup_filt.n3 205.059
R29399 pwup_filt.n6 pwup_filt.n5 205.059
R29400 pwup_filt.n8 pwup_filt.n7 205.059
R29401 pwup_filt.n10 pwup_filt.n9 205.059
R29402 pwup_filt.n12 pwup_filt.n11 205.059
R29403 pwup_filt.n14 pwup_filt.n13 205.059
R29404 pwup_filt.n15 pwup_filt.t32 175.169
R29405 pwup_filt.n16 pwup_filt.n15 153.385
R29406 pwup_filt.n22 pwup_filt.n20 133.534
R29407 pwup_filt.n22 pwup_filt.n21 99.1759
R29408 pwup_filt.n24 pwup_filt.n23 99.1759
R29409 pwup_filt.n26 pwup_filt.n25 99.1759
R29410 pwup_filt.n28 pwup_filt.n27 99.1759
R29411 pwup_filt.n30 pwup_filt.n29 99.1759
R29412 pwup_filt.n32 pwup_filt.n31 99.1759
R29413 pwup_filt pwup_filt.n33 97.4305
R29414 pwup_filt.n4 pwup_filt.n2 38.4005
R29415 pwup_filt.n6 pwup_filt.n4 38.4005
R29416 pwup_filt.n8 pwup_filt.n6 38.4005
R29417 pwup_filt.n10 pwup_filt.n8 38.4005
R29418 pwup_filt.n12 pwup_filt.n10 38.4005
R29419 pwup_filt.n14 pwup_filt.n12 38.4005
R29420 pwup_filt.n24 pwup_filt.n22 34.3584
R29421 pwup_filt.n26 pwup_filt.n24 34.3584
R29422 pwup_filt.n28 pwup_filt.n26 34.3584
R29423 pwup_filt.n30 pwup_filt.n28 34.3584
R29424 pwup_filt.n32 pwup_filt.n30 34.3584
R29425 pwup_filt.n34 pwup_filt.n32 34.3584
R29426 pwup_filt.n13 pwup_filt.t26 26.5955
R29427 pwup_filt.n13 pwup_filt.t29 26.5955
R29428 pwup_filt.n0 pwup_filt.t21 26.5955
R29429 pwup_filt.n0 pwup_filt.t25 26.5955
R29430 pwup_filt.n1 pwup_filt.t16 26.5955
R29431 pwup_filt.n1 pwup_filt.t24 26.5955
R29432 pwup_filt.n3 pwup_filt.t23 26.5955
R29433 pwup_filt.n3 pwup_filt.t19 26.5955
R29434 pwup_filt.n5 pwup_filt.t22 26.5955
R29435 pwup_filt.n5 pwup_filt.t20 26.5955
R29436 pwup_filt.n7 pwup_filt.t18 26.5955
R29437 pwup_filt.n7 pwup_filt.t31 26.5955
R29438 pwup_filt.n9 pwup_filt.t30 26.5955
R29439 pwup_filt.n9 pwup_filt.t28 26.5955
R29440 pwup_filt.n11 pwup_filt.t27 26.5955
R29441 pwup_filt.n11 pwup_filt.t17 26.5955
R29442 pwup_filt pwup_filt.n16 26.2517
R29443 pwup_filt.n33 pwup_filt.t0 24.9236
R29444 pwup_filt.n33 pwup_filt.t3 24.9236
R29445 pwup_filt.n20 pwup_filt.t11 24.9236
R29446 pwup_filt.n20 pwup_filt.t15 24.9236
R29447 pwup_filt.n21 pwup_filt.t6 24.9236
R29448 pwup_filt.n21 pwup_filt.t14 24.9236
R29449 pwup_filt.n23 pwup_filt.t13 24.9236
R29450 pwup_filt.n23 pwup_filt.t9 24.9236
R29451 pwup_filt.n25 pwup_filt.t12 24.9236
R29452 pwup_filt.n25 pwup_filt.t10 24.9236
R29453 pwup_filt.n27 pwup_filt.t8 24.9236
R29454 pwup_filt.n27 pwup_filt.t5 24.9236
R29455 pwup_filt.n29 pwup_filt.t4 24.9236
R29456 pwup_filt.n29 pwup_filt.t2 24.9236
R29457 pwup_filt.n31 pwup_filt.t1 24.9236
R29458 pwup_filt.n31 pwup_filt.t7 24.9236
R29459 pwup_filt.n18 pwup_filt.n17 13.9767
R29460 pwup_filt.n19 pwup_filt.n14 12.6066
R29461 pwup_filt pwup_filt.n34 11.4429
R29462 pwup_filt.n19 pwup_filt.n18 10.4495
R29463 pwup_filt.n18 pwup_filt 9.99427
R29464 pwup_filt pwup_filt.n19 5.81868
R29465 pwup_filt.n16 pwup_filt 2.94104
R29466 pwup_filt.n34 pwup_filt 1.74595
R29467 pwup_filt.n17 pwup_filt 0.203775
R29468 pwup_filt.n17 pwup_filt 0.162258
R29469 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n37 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n35 271.065
R29470 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n26 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n24 205.059
R29471 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n37 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n36 180.583
R29472 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n32 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n31 156.462
R29473 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n14 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n0 69.6745
R29474 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n20 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n22 69.6745
R29475 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n9 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n21 69.6745
R29476 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n18 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n19 69.6745
R29477 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n4 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A 69.6745
R29478 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n29 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n23 155.492
R29479 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n30 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.t22 113.543
R29480 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n26 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n25 98.5495
R29481 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n27 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.t39 93.5093
R29482 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n1 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.t21 92.5445
R29483 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n2 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.t20 92.5445
R29484 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n3 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.t16 92.5445
R29485 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n5 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.t15 92.5445
R29486 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n6 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.t12 92.5445
R29487 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n7 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.t24 92.5445
R29488 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n8 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.t11 92.5445
R29489 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n10 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.t19 92.5445
R29490 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n11 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.t18 92.5445
R29491 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n12 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.t14 92.5445
R29492 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n13 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.t13 92.5445
R29493 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n15 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.t37 92.5445
R29494 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n16 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.t28 92.5445
R29495 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n17 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.t8 92.5445
R29496 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n2 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n3 84.8982
R29497 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n6 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n5 84.8982
R29498 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n7 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n8 84.8982
R29499 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n11 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n10 84.8982
R29500 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n12 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n13 84.8982
R29501 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n17 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n15 84.8982
R29502 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n0 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n28 69.8017
R29503 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n27 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.t17 67.9625
R29504 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n30 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.t36 67.7525
R29505 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n31 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n29 61.8937
R29506 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n1 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n30 57.5119
R29507 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n16 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n27 57.5119
R29508 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n1 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.t35 46.7545
R29509 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n2 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.t9 46.7545
R29510 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n3 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.t31 46.7545
R29511 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n5 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.t30 46.7545
R29512 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n6 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.t26 46.7545
R29513 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n7 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.t38 46.7545
R29514 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n8 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.t34 46.7545
R29515 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n10 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.t33 46.7545
R29516 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n11 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.t32 46.7545
R29517 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n12 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.t29 46.7545
R29518 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n13 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.t27 46.7545
R29519 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n15 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.t25 46.7545
R29520 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n16 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.t10 46.7545
R29521 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n17 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.t23 46.7545
R29522 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n13 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n14 37.9969
R29523 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n11 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n22 37.9969
R29524 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n8 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n9 37.9969
R29525 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n6 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n19 37.9969
R29526 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n3 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n4 37.9969
R29527 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n28 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n17 37.9906
R29528 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n28 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n16 37.9727
R29529 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n15 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n14 37.9654
R29530 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n22 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n12 37.9654
R29531 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n10 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n9 37.9654
R29532 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n19 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n7 37.9654
R29533 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n5 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n4 37.9654
R29534 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n25 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.t7 21.2805
R29535 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n25 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.t6 21.2805
R29536 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n24 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.t5 21.2805
R29537 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n24 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.t4 21.2805
R29538 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n35 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.t1 17.8272
R29539 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n35 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.t0 17.8272
R29540 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n36 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.t3 17.8272
R29541 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n36 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.t2 17.8272
R29542 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n32 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n23 13.9641
R29543 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n34 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n26 13.1544
R29544 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n29 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n2 12.0505
R29545 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n31 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n1 12.0505
R29546 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n23 9.3005
R29547 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n32 9.3005
R29548 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n37 6.86595
R29549 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n34 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n33 6.51686
R29550 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n0 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A 6.20638
R29551 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n33 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A 5.52042
R29552 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n0 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A 5.08202
R29553 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n20 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A 5.05932
R29554 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n0 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A 4.2342
R29555 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n21 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A 3.91226
R29556 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n20 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A 3.38637
R29557 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n33 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A 3.14232
R29558 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n18 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A 2.76521
R29559 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n21 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A 2.53854
R29560 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n0 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n20 1.692
R29561 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n18 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A 1.69072
R29562 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n34 1.51323
R29563 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n21 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n20 1.02288
R29564 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n21 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n18 1.02288
R29565 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n18 1.02288
R29566 por_dig_0.clknet_1_0__leaf_osc_ck.n18 por_dig_0.clknet_1_0__leaf_osc_ck.n16 333.392
R29567 por_dig_0.clknet_1_0__leaf_osc_ck.n18 por_dig_0.clknet_1_0__leaf_osc_ck.n17 301.392
R29568 por_dig_0.clknet_1_0__leaf_osc_ck.n20 por_dig_0.clknet_1_0__leaf_osc_ck.n19 301.392
R29569 por_dig_0.clknet_1_0__leaf_osc_ck.n22 por_dig_0.clknet_1_0__leaf_osc_ck.n21 301.392
R29570 por_dig_0.clknet_1_0__leaf_osc_ck.n24 por_dig_0.clknet_1_0__leaf_osc_ck.n23 301.392
R29571 por_dig_0.clknet_1_0__leaf_osc_ck.n57 por_dig_0.clknet_1_0__leaf_osc_ck.n15 301.392
R29572 por_dig_0.clknet_1_0__leaf_osc_ck por_dig_0.clknet_1_0__leaf_osc_ck.n58 297.752
R29573 por_dig_0.clknet_1_0__leaf_osc_ck.n52 por_dig_0.clknet_1_0__leaf_osc_ck.t48 294.557
R29574 por_dig_0.clknet_1_0__leaf_osc_ck.n47 por_dig_0.clknet_1_0__leaf_osc_ck.t41 294.557
R29575 por_dig_0.clknet_1_0__leaf_osc_ck.n43 por_dig_0.clknet_1_0__leaf_osc_ck.t43 294.557
R29576 por_dig_0.clknet_1_0__leaf_osc_ck.n31 por_dig_0.clknet_1_0__leaf_osc_ck.t39 294.557
R29577 por_dig_0.clknet_1_0__leaf_osc_ck.n37 por_dig_0.clknet_1_0__leaf_osc_ck.t33 294.557
R29578 por_dig_0.clknet_1_0__leaf_osc_ck.n35 por_dig_0.clknet_1_0__leaf_osc_ck.t45 294.557
R29579 por_dig_0.clknet_1_0__leaf_osc_ck.n33 por_dig_0.clknet_1_0__leaf_osc_ck.t46 294.557
R29580 por_dig_0.clknet_1_0__leaf_osc_ck.n28 por_dig_0.clknet_1_0__leaf_osc_ck.t40 294.557
R29581 por_dig_0.clknet_1_0__leaf_osc_ck.n26 por_dig_0.clknet_1_0__leaf_osc_ck.t32 294.557
R29582 por_dig_0.clknet_1_0__leaf_osc_ck.n55 por_dig_0.clknet_1_0__leaf_osc_ck.n25 293.348
R29583 por_dig_0.clknet_1_0__leaf_osc_ck.n2 por_dig_0.clknet_1_0__leaf_osc_ck.n0 248.638
R29584 por_dig_0.clknet_1_0__leaf_osc_ck.n52 por_dig_0.clknet_1_0__leaf_osc_ck.t37 211.01
R29585 por_dig_0.clknet_1_0__leaf_osc_ck.n47 por_dig_0.clknet_1_0__leaf_osc_ck.t42 211.01
R29586 por_dig_0.clknet_1_0__leaf_osc_ck.n43 por_dig_0.clknet_1_0__leaf_osc_ck.t44 211.01
R29587 por_dig_0.clknet_1_0__leaf_osc_ck.n31 por_dig_0.clknet_1_0__leaf_osc_ck.t47 211.01
R29588 por_dig_0.clknet_1_0__leaf_osc_ck.n37 por_dig_0.clknet_1_0__leaf_osc_ck.t34 211.01
R29589 por_dig_0.clknet_1_0__leaf_osc_ck.n35 por_dig_0.clknet_1_0__leaf_osc_ck.t35 211.01
R29590 por_dig_0.clknet_1_0__leaf_osc_ck.n33 por_dig_0.clknet_1_0__leaf_osc_ck.t36 211.01
R29591 por_dig_0.clknet_1_0__leaf_osc_ck.n28 por_dig_0.clknet_1_0__leaf_osc_ck.t49 211.01
R29592 por_dig_0.clknet_1_0__leaf_osc_ck.n26 por_dig_0.clknet_1_0__leaf_osc_ck.t38 211.01
R29593 por_dig_0.clknet_1_0__leaf_osc_ck.n2 por_dig_0.clknet_1_0__leaf_osc_ck.n1 203.463
R29594 por_dig_0.clknet_1_0__leaf_osc_ck.n4 por_dig_0.clknet_1_0__leaf_osc_ck.n3 203.463
R29595 por_dig_0.clknet_1_0__leaf_osc_ck.n8 por_dig_0.clknet_1_0__leaf_osc_ck.n7 203.463
R29596 por_dig_0.clknet_1_0__leaf_osc_ck.n10 por_dig_0.clknet_1_0__leaf_osc_ck.n9 203.463
R29597 por_dig_0.clknet_1_0__leaf_osc_ck.n12 por_dig_0.clknet_1_0__leaf_osc_ck.n11 203.463
R29598 por_dig_0.clknet_1_0__leaf_osc_ck.n6 por_dig_0.clknet_1_0__leaf_osc_ck.n5 202.456
R29599 por_dig_0.clknet_1_0__leaf_osc_ck.n14 por_dig_0.clknet_1_0__leaf_osc_ck.n13 200.212
R29600 por_dig_0.clknet_1_0__leaf_osc_ck por_dig_0.clknet_1_0__leaf_osc_ck.n35 156.207
R29601 por_dig_0.clknet_1_0__leaf_osc_ck por_dig_0.clknet_1_0__leaf_osc_ck.n33 156.207
R29602 por_dig_0.clknet_1_0__leaf_osc_ck por_dig_0.clknet_1_0__leaf_osc_ck.n28 156.207
R29603 por_dig_0.clknet_1_0__leaf_osc_ck.n32 por_dig_0.clknet_1_0__leaf_osc_ck.n31 153.097
R29604 por_dig_0.clknet_1_0__leaf_osc_ck.n53 por_dig_0.clknet_1_0__leaf_osc_ck.n52 152
R29605 por_dig_0.clknet_1_0__leaf_osc_ck.n48 por_dig_0.clknet_1_0__leaf_osc_ck.n47 152
R29606 por_dig_0.clknet_1_0__leaf_osc_ck.n44 por_dig_0.clknet_1_0__leaf_osc_ck.n43 152
R29607 por_dig_0.clknet_1_0__leaf_osc_ck.n38 por_dig_0.clknet_1_0__leaf_osc_ck.n37 152
R29608 por_dig_0.clknet_1_0__leaf_osc_ck.n27 por_dig_0.clknet_1_0__leaf_osc_ck.n26 152
R29609 por_dig_0.clknet_1_0__leaf_osc_ck.n4 por_dig_0.clknet_1_0__leaf_osc_ck.n2 45.177
R29610 por_dig_0.clknet_1_0__leaf_osc_ck.n10 por_dig_0.clknet_1_0__leaf_osc_ck.n8 45.177
R29611 por_dig_0.clknet_1_0__leaf_osc_ck.n12 por_dig_0.clknet_1_0__leaf_osc_ck.n10 45.177
R29612 por_dig_0.clknet_1_0__leaf_osc_ck.n6 por_dig_0.clknet_1_0__leaf_osc_ck.n4 44.0476
R29613 por_dig_0.clknet_1_0__leaf_osc_ck.n8 por_dig_0.clknet_1_0__leaf_osc_ck.n6 44.0476
R29614 por_dig_0.clknet_1_0__leaf_osc_ck.n0 por_dig_0.clknet_1_0__leaf_osc_ck.t5 40.0005
R29615 por_dig_0.clknet_1_0__leaf_osc_ck.n0 por_dig_0.clknet_1_0__leaf_osc_ck.t8 40.0005
R29616 por_dig_0.clknet_1_0__leaf_osc_ck.n1 por_dig_0.clknet_1_0__leaf_osc_ck.t14 40.0005
R29617 por_dig_0.clknet_1_0__leaf_osc_ck.n1 por_dig_0.clknet_1_0__leaf_osc_ck.t4 40.0005
R29618 por_dig_0.clknet_1_0__leaf_osc_ck.n3 por_dig_0.clknet_1_0__leaf_osc_ck.t12 40.0005
R29619 por_dig_0.clknet_1_0__leaf_osc_ck.n3 por_dig_0.clknet_1_0__leaf_osc_ck.t1 40.0005
R29620 por_dig_0.clknet_1_0__leaf_osc_ck.n5 por_dig_0.clknet_1_0__leaf_osc_ck.t10 40.0005
R29621 por_dig_0.clknet_1_0__leaf_osc_ck.n5 por_dig_0.clknet_1_0__leaf_osc_ck.t0 40.0005
R29622 por_dig_0.clknet_1_0__leaf_osc_ck.n7 por_dig_0.clknet_1_0__leaf_osc_ck.t9 40.0005
R29623 por_dig_0.clknet_1_0__leaf_osc_ck.n7 por_dig_0.clknet_1_0__leaf_osc_ck.t15 40.0005
R29624 por_dig_0.clknet_1_0__leaf_osc_ck.n9 por_dig_0.clknet_1_0__leaf_osc_ck.t6 40.0005
R29625 por_dig_0.clknet_1_0__leaf_osc_ck.n9 por_dig_0.clknet_1_0__leaf_osc_ck.t13 40.0005
R29626 por_dig_0.clknet_1_0__leaf_osc_ck.n11 por_dig_0.clknet_1_0__leaf_osc_ck.t3 40.0005
R29627 por_dig_0.clknet_1_0__leaf_osc_ck.n11 por_dig_0.clknet_1_0__leaf_osc_ck.t11 40.0005
R29628 por_dig_0.clknet_1_0__leaf_osc_ck.n13 por_dig_0.clknet_1_0__leaf_osc_ck.t2 40.0005
R29629 por_dig_0.clknet_1_0__leaf_osc_ck.n13 por_dig_0.clknet_1_0__leaf_osc_ck.t7 40.0005
R29630 por_dig_0.clknet_1_0__leaf_osc_ck.n20 por_dig_0.clknet_1_0__leaf_osc_ck.n18 32.0005
R29631 por_dig_0.clknet_1_0__leaf_osc_ck.n22 por_dig_0.clknet_1_0__leaf_osc_ck.n20 32.0005
R29632 por_dig_0.clknet_1_0__leaf_osc_ck.n57 por_dig_0.clknet_1_0__leaf_osc_ck.n56 32.0005
R29633 por_dig_0.clknet_1_0__leaf_osc_ck.n56 por_dig_0.clknet_1_0__leaf_osc_ck.n24 32.0005
R29634 por_dig_0.clknet_1_0__leaf_osc_ck.n24 por_dig_0.clknet_1_0__leaf_osc_ck.n22 31.2005
R29635 por_dig_0.clknet_1_0__leaf_osc_ck.n16 por_dig_0.clknet_1_0__leaf_osc_ck.t30 27.5805
R29636 por_dig_0.clknet_1_0__leaf_osc_ck.n16 por_dig_0.clknet_1_0__leaf_osc_ck.t17 27.5805
R29637 por_dig_0.clknet_1_0__leaf_osc_ck.n17 por_dig_0.clknet_1_0__leaf_osc_ck.t23 27.5805
R29638 por_dig_0.clknet_1_0__leaf_osc_ck.n17 por_dig_0.clknet_1_0__leaf_osc_ck.t29 27.5805
R29639 por_dig_0.clknet_1_0__leaf_osc_ck.n19 por_dig_0.clknet_1_0__leaf_osc_ck.t21 27.5805
R29640 por_dig_0.clknet_1_0__leaf_osc_ck.n19 por_dig_0.clknet_1_0__leaf_osc_ck.t26 27.5805
R29641 por_dig_0.clknet_1_0__leaf_osc_ck.n21 por_dig_0.clknet_1_0__leaf_osc_ck.t19 27.5805
R29642 por_dig_0.clknet_1_0__leaf_osc_ck.n21 por_dig_0.clknet_1_0__leaf_osc_ck.t25 27.5805
R29643 por_dig_0.clknet_1_0__leaf_osc_ck.n23 por_dig_0.clknet_1_0__leaf_osc_ck.t18 27.5805
R29644 por_dig_0.clknet_1_0__leaf_osc_ck.n23 por_dig_0.clknet_1_0__leaf_osc_ck.t24 27.5805
R29645 por_dig_0.clknet_1_0__leaf_osc_ck.n15 por_dig_0.clknet_1_0__leaf_osc_ck.t28 27.5805
R29646 por_dig_0.clknet_1_0__leaf_osc_ck.n15 por_dig_0.clknet_1_0__leaf_osc_ck.t20 27.5805
R29647 por_dig_0.clknet_1_0__leaf_osc_ck.n58 por_dig_0.clknet_1_0__leaf_osc_ck.t27 27.5805
R29648 por_dig_0.clknet_1_0__leaf_osc_ck.n58 por_dig_0.clknet_1_0__leaf_osc_ck.t16 27.5805
R29649 por_dig_0.clknet_1_0__leaf_osc_ck.n25 por_dig_0.clknet_1_0__leaf_osc_ck.t31 27.5805
R29650 por_dig_0.clknet_1_0__leaf_osc_ck.n25 por_dig_0.clknet_1_0__leaf_osc_ck.t22 27.5805
R29651 por_dig_0.clknet_1_0__leaf_osc_ck.n54 por_dig_0.clknet_1_0__leaf_osc_ck 24.6249
R29652 por_dig_0.clknet_1_0__leaf_osc_ck.n40 por_dig_0.clknet_1_0__leaf_osc_ck.n36 19.2663
R29653 por_dig_0.clknet_1_0__leaf_osc_ck.n46 por_dig_0.clknet_1_0__leaf_osc_ck.n42 14.3618
R29654 por_dig_0.clknet_1_0__leaf_osc_ck.n42 por_dig_0.clknet_1_0__leaf_osc_ck.n41 14.1296
R29655 por_dig_0.clknet_1_0__leaf_osc_ck.n55 por_dig_0.clknet_1_0__leaf_osc_ck.n54 14.0387
R29656 por_dig_0.clknet_1_0__leaf_osc_ck.n40 por_dig_0.clknet_1_0__leaf_osc_ck.n39 13.8005
R29657 por_dig_0.clknet_1_0__leaf_osc_ck.n14 por_dig_0.clknet_1_0__leaf_osc_ck.n12 13.177
R29658 por_dig_0.clknet_1_0__leaf_osc_ck.n51 por_dig_0.clknet_1_0__leaf_osc_ck.n50 11.9371
R29659 por_dig_0.clknet_1_0__leaf_osc_ck.n41 por_dig_0.clknet_1_0__leaf_osc_ck.n34 11.369
R29660 por_dig_0.clknet_1_0__leaf_osc_ck por_dig_0.clknet_1_0__leaf_osc_ck.n53 10.4234
R29661 por_dig_0.clknet_1_0__leaf_osc_ck por_dig_0.clknet_1_0__leaf_osc_ck.n27 10.4234
R29662 por_dig_0.clknet_1_0__leaf_osc_ck.n50 por_dig_0.clknet_1_0__leaf_osc_ck.n46 10.2297
R29663 por_dig_0.clknet_1_0__leaf_osc_ck por_dig_0.clknet_1_0__leaf_osc_ck.n57 10.2022
R29664 por_dig_0.clknet_1_0__leaf_osc_ck.n42 por_dig_0.clknet_1_0__leaf_osc_ck.n32 9.73846
R29665 por_dig_0.clknet_1_0__leaf_osc_ck.n49 por_dig_0.clknet_1_0__leaf_osc_ck 9.32621
R29666 por_dig_0.clknet_1_0__leaf_osc_ck.n45 por_dig_0.clknet_1_0__leaf_osc_ck 9.32621
R29667 por_dig_0.clknet_1_0__leaf_osc_ck.n39 por_dig_0.clknet_1_0__leaf_osc_ck 9.32621
R29668 por_dig_0.clknet_1_0__leaf_osc_ck.n36 por_dig_0.clknet_1_0__leaf_osc_ck 9.32621
R29669 por_dig_0.clknet_1_0__leaf_osc_ck.n34 por_dig_0.clknet_1_0__leaf_osc_ck 9.32621
R29670 por_dig_0.clknet_1_0__leaf_osc_ck.n29 por_dig_0.clknet_1_0__leaf_osc_ck 9.32621
R29671 por_dig_0.clknet_1_0__leaf_osc_ck.n46 por_dig_0.clknet_1_0__leaf_osc_ck.n45 9.3005
R29672 por_dig_0.clknet_1_0__leaf_osc_ck.n50 por_dig_0.clknet_1_0__leaf_osc_ck.n49 9.3005
R29673 por_dig_0.clknet_1_0__leaf_osc_ck.n30 por_dig_0.clknet_1_0__leaf_osc_ck.n29 9.3005
R29674 por_dig_0.clknet_1_0__leaf_osc_ck.n56 por_dig_0.clknet_1_0__leaf_osc_ck.n55 8.04533
R29675 por_dig_0.clknet_1_0__leaf_osc_ck.n41 por_dig_0.clknet_1_0__leaf_osc_ck.n40 7.40435
R29676 por_dig_0.clknet_1_0__leaf_osc_ck.n51 por_dig_0.clknet_1_0__leaf_osc_ck.n30 5.63391
R29677 por_dig_0.clknet_1_0__leaf_osc_ck.n54 por_dig_0.clknet_1_0__leaf_osc_ck.n51 3.75599
R29678 por_dig_0.clknet_1_0__leaf_osc_ck.n32 por_dig_0.clknet_1_0__leaf_osc_ck 3.10907
R29679 por_dig_0.clknet_1_0__leaf_osc_ck.n36 por_dig_0.clknet_1_0__leaf_osc_ck 3.10907
R29680 por_dig_0.clknet_1_0__leaf_osc_ck.n34 por_dig_0.clknet_1_0__leaf_osc_ck 3.10907
R29681 por_dig_0.clknet_1_0__leaf_osc_ck.n29 por_dig_0.clknet_1_0__leaf_osc_ck 3.10907
R29682 por_dig_0.clknet_1_0__leaf_osc_ck.n53 por_dig_0.clknet_1_0__leaf_osc_ck 2.01193
R29683 por_dig_0.clknet_1_0__leaf_osc_ck.n48 por_dig_0.clknet_1_0__leaf_osc_ck 2.01193
R29684 por_dig_0.clknet_1_0__leaf_osc_ck.n44 por_dig_0.clknet_1_0__leaf_osc_ck 2.01193
R29685 por_dig_0.clknet_1_0__leaf_osc_ck.n38 por_dig_0.clknet_1_0__leaf_osc_ck 2.01193
R29686 por_dig_0.clknet_1_0__leaf_osc_ck.n27 por_dig_0.clknet_1_0__leaf_osc_ck 2.01193
R29687 por_dig_0.clknet_1_0__leaf_osc_ck por_dig_0.clknet_1_0__leaf_osc_ck.n14 1.26402
R29688 por_dig_0.clknet_1_0__leaf_osc_ck.n49 por_dig_0.clknet_1_0__leaf_osc_ck.n48 1.09764
R29689 por_dig_0.clknet_1_0__leaf_osc_ck.n45 por_dig_0.clknet_1_0__leaf_osc_ck.n44 1.09764
R29690 por_dig_0.clknet_1_0__leaf_osc_ck.n39 por_dig_0.clknet_1_0__leaf_osc_ck.n38 1.09764
R29691 por_dig_0.clknet_1_0__leaf_osc_ck.n30 por_dig_0.clknet_1_0__leaf_osc_ck 0.565912
R29692 por_ana_0.schmitt_trigger_0.out.n8 por_ana_0.schmitt_trigger_0.out.t10 248.236
R29693 por_ana_0.schmitt_trigger_0.out.n6 por_ana_0.schmitt_trigger_0.out.t12 240.778
R29694 por_ana_0.schmitt_trigger_0.out.n7 por_ana_0.schmitt_trigger_0.out.t4 240.613
R29695 por_ana_0.schmitt_trigger_0.out.n6 por_ana_0.schmitt_trigger_0.out.t5 240.349
R29696 por_ana_0.schmitt_trigger_0.out.n5 por_ana_0.schmitt_trigger_0.out.t1 236.369
R29697 por_ana_0.schmitt_trigger_0.out.n0 por_ana_0.schmitt_trigger_0.out.t9 212.081
R29698 por_ana_0.schmitt_trigger_0.out.n2 por_ana_0.schmitt_trigger_0.out.t6 212.081
R29699 por_ana_0.schmitt_trigger_0.out.n15 por_ana_0.schmitt_trigger_0.out.t7 212.081
R29700 por_ana_0.schmitt_trigger_0.out.n3 por_ana_0.schmitt_trigger_0.out.t8 212.081
R29701 por_ana_0.schmitt_trigger_0.out.n5 por_ana_0.schmitt_trigger_0.out.n4 207.585
R29702 por_ana_0.schmitt_trigger_0.out.n12 por_ana_0.schmitt_trigger_0.out.n3 188.516
R29703 por_ana_0.sky130_fd_sc_hd__inv_4_0.A por_ana_0.schmitt_trigger_0.out.n1 154.304
R29704 por_ana_0.schmitt_trigger_0.out.n14 por_ana_0.schmitt_trigger_0.out.n13 152
R29705 por_ana_0.schmitt_trigger_0.out.n17 por_ana_0.schmitt_trigger_0.out.n16 152
R29706 por_ana_0.schmitt_trigger_0.out.n0 por_ana_0.schmitt_trigger_0.out.t15 139.78
R29707 por_ana_0.schmitt_trigger_0.out.n2 por_ana_0.schmitt_trigger_0.out.t11 139.78
R29708 por_ana_0.schmitt_trigger_0.out.n15 por_ana_0.schmitt_trigger_0.out.t13 139.78
R29709 por_ana_0.schmitt_trigger_0.out.n3 por_ana_0.schmitt_trigger_0.out.t14 139.78
R29710 por_ana_0.schmitt_trigger_0.out.n10 por_ana_0.schmitt_trigger_0.out.t0 91.727
R29711 por_ana_0.schmitt_trigger_0.out.n1 por_ana_0.schmitt_trigger_0.out.n0 30.6732
R29712 por_ana_0.schmitt_trigger_0.out.n2 por_ana_0.schmitt_trigger_0.out.n1 30.6732
R29713 por_ana_0.schmitt_trigger_0.out.n16 por_ana_0.schmitt_trigger_0.out.n2 30.6732
R29714 por_ana_0.schmitt_trigger_0.out.n16 por_ana_0.schmitt_trigger_0.out.n15 30.6732
R29715 por_ana_0.schmitt_trigger_0.out.n15 por_ana_0.schmitt_trigger_0.out.n14 30.6732
R29716 por_ana_0.schmitt_trigger_0.out.n14 por_ana_0.schmitt_trigger_0.out.n3 30.6732
R29717 por_ana_0.schmitt_trigger_0.out.n4 por_ana_0.schmitt_trigger_0.out.t2 28.5655
R29718 por_ana_0.schmitt_trigger_0.out.n4 por_ana_0.schmitt_trigger_0.out.t3 28.5655
R29719 por_ana_0.schmitt_trigger_0.out.n11 por_ana_0.schmitt_trigger_0.out.n10 20.1312
R29720 por_ana_0.sky130_fd_sc_hd__inv_4_0.A por_ana_0.schmitt_trigger_0.out.n17 19.2005
R29721 por_ana_0.sky130_fd_sc_hd__inv_4_0.A por_ana_0.schmitt_trigger_0.out.n12 17.1525
R29722 por_ana_0.schmitt_trigger_0.out.n11 por_ana_0.sky130_fd_sc_hd__inv_4_0.A 12.8005
R29723 por_ana_0.schmitt_trigger_0.out.n9 por_ana_0.schmitt_trigger_0.out.n5 8.66251
R29724 por_ana_0.schmitt_trigger_0.out.n13 por_ana_0.sky130_fd_sc_hd__inv_4_0.A 6.4005
R29725 por_ana_0.schmitt_trigger_0.out.n12 por_ana_0.sky130_fd_sc_hd__inv_4_0.A 6.4005
R29726 por_ana_0.schmitt_trigger_0.out.n8 por_ana_0.schmitt_trigger_0.out.n7 4.94425
R29727 por_ana_0.schmitt_trigger_0.out.n17 por_ana_0.sky130_fd_sc_hd__inv_4_0.A 4.3525
R29728 por_ana_0.schmitt_trigger_0.out.n13 por_ana_0.schmitt_trigger_0.out.n11 4.3525
R29729 por_ana_0.schmitt_trigger_0.out.n9 por_ana_0.schmitt_trigger_0.out.n8 4.05633
R29730 por_ana_0.schmitt_trigger_0.out.n10 por_ana_0.schmitt_trigger_0.out.n9 0.230017
R29731 por_ana_0.schmitt_trigger_0.out.n7 por_ana_0.schmitt_trigger_0.out.n6 0.117348
R29732 por_dig_0.por_unbuf.n32 por_dig_0.por_unbuf.n29 585.503
R29733 por_dig_0.por_unbuf.n33 por_dig_0.por_unbuf.n32 585
R29734 por_dig_0.por_unbuf.n1 por_dig_0.por_unbuf.t8 212.081
R29735 por_dig_0.por_unbuf.n3 por_dig_0.por_unbuf.t21 212.081
R29736 por_dig_0.por_unbuf.n0 por_dig_0.por_unbuf.t4 212.081
R29737 por_dig_0.por_unbuf.n8 por_dig_0.por_unbuf.t7 212.081
R29738 por_dig_0.por_unbuf.n12 por_dig_0.por_unbuf.t6 212.081
R29739 por_dig_0.por_unbuf.n14 por_dig_0.por_unbuf.t19 212.081
R29740 por_dig_0.por_unbuf.n11 por_dig_0.por_unbuf.t20 212.081
R29741 por_dig_0.por_unbuf.n19 por_dig_0.por_unbuf.t5 212.081
R29742 por_dig_0.por_unbuf.n9 por_dig_0.por_unbuf.n8 188.516
R29743 por_dig_0.por_unbuf.n20 por_dig_0.por_unbuf.n19 188.516
R29744 por_dig_0.por_unbuf.n23 por_dig_0.por_unbuf.t9 186.374
R29745 por_dig_0.por_unbuf.n31 por_dig_0.por_unbuf.n30 185
R29746 por_dig_0.por_unbuf.n23 por_dig_0.por_unbuf.t18 170.308
R29747 por_dig_0.por_unbuf.n24 por_dig_0.por_unbuf 155.511
R29748 por_dig_0.por_unbuf.n2 por_dig_0.por_unbuf 154.304
R29749 por_dig_0.por_unbuf.n13 por_dig_0.por_unbuf 154.304
R29750 por_dig_0.por_unbuf.n25 por_dig_0.por_unbuf.n24 153.462
R29751 por_dig_0.por_unbuf.n7 por_dig_0.por_unbuf.n6 152
R29752 por_dig_0.por_unbuf.n5 por_dig_0.por_unbuf.n4 152
R29753 por_dig_0.por_unbuf.n18 por_dig_0.por_unbuf.n17 152
R29754 por_dig_0.por_unbuf.n16 por_dig_0.por_unbuf.n15 152
R29755 por_dig_0.por_unbuf.n1 por_dig_0.por_unbuf.t17 139.78
R29756 por_dig_0.por_unbuf.n3 por_dig_0.por_unbuf.t12 139.78
R29757 por_dig_0.por_unbuf.n0 por_dig_0.por_unbuf.t13 139.78
R29758 por_dig_0.por_unbuf.n8 por_dig_0.por_unbuf.t16 139.78
R29759 por_dig_0.por_unbuf.n12 por_dig_0.por_unbuf.t15 139.78
R29760 por_dig_0.por_unbuf.n14 por_dig_0.por_unbuf.t10 139.78
R29761 por_dig_0.por_unbuf.n11 por_dig_0.por_unbuf.t11 139.78
R29762 por_dig_0.por_unbuf.n19 por_dig_0.por_unbuf.t14 139.78
R29763 por_dig_0.por_unbuf.n24 por_dig_0.por_unbuf.n23 101.513
R29764 por_dig_0.por_unbuf por_dig_0.por_unbuf.n31 81.3181
R29765 por_dig_0.por_unbuf.n2 por_dig_0.por_unbuf.n1 30.6732
R29766 por_dig_0.por_unbuf.n3 por_dig_0.por_unbuf.n2 30.6732
R29767 por_dig_0.por_unbuf.n4 por_dig_0.por_unbuf.n3 30.6732
R29768 por_dig_0.por_unbuf.n4 por_dig_0.por_unbuf.n0 30.6732
R29769 por_dig_0.por_unbuf.n7 por_dig_0.por_unbuf.n0 30.6732
R29770 por_dig_0.por_unbuf.n8 por_dig_0.por_unbuf.n7 30.6732
R29771 por_dig_0.por_unbuf.n13 por_dig_0.por_unbuf.n12 30.6732
R29772 por_dig_0.por_unbuf.n14 por_dig_0.por_unbuf.n13 30.6732
R29773 por_dig_0.por_unbuf.n15 por_dig_0.por_unbuf.n14 30.6732
R29774 por_dig_0.por_unbuf.n15 por_dig_0.por_unbuf.n11 30.6732
R29775 por_dig_0.por_unbuf.n18 por_dig_0.por_unbuf.n11 30.6732
R29776 por_dig_0.por_unbuf.n19 por_dig_0.por_unbuf.n18 30.6732
R29777 por_dig_0.por_unbuf.n32 por_dig_0.por_unbuf.t2 26.5955
R29778 por_dig_0.por_unbuf.n32 por_dig_0.por_unbuf.t3 26.5955
R29779 por_dig_0.por_unbuf.n30 por_dig_0.por_unbuf.t1 24.9236
R29780 por_dig_0.por_unbuf.n30 por_dig_0.por_unbuf.t0 24.9236
R29781 por_dig_0.por_unbuf.n28 por_dig_0.por_unbuf.n27 24.6442
R29782 por_dig_0.por_unbuf.n22 por_dig_0.por_unbuf.n10 21.5696
R29783 por_dig_0.por_unbuf.n22 por_dig_0.por_unbuf.n21 20.7505
R29784 por_dig_0.por_unbuf.n5 por_dig_0.por_unbuf 19.2005
R29785 por_dig_0.por_unbuf.n16 por_dig_0.por_unbuf 19.2005
R29786 por_dig_0.por_unbuf.n6 por_dig_0.por_unbuf 17.1525
R29787 por_dig_0.por_unbuf.n17 por_dig_0.por_unbuf 17.1525
R29788 por_dig_0.por_unbuf por_dig_0.por_unbuf.n33 15.5613
R29789 por_dig_0.por_unbuf.n27 por_dig_0.por_unbuf.n26 13.8005
R29790 por_dig_0.por_unbuf.n21 por_dig_0.por_unbuf 12.5445
R29791 por_dig_0.por_unbuf.n27 por_dig_0.por_unbuf.n22 11.5344
R29792 por_dig_0.por_unbuf.n29 por_dig_0.por_unbuf 10.6873
R29793 por_dig_0.por_unbuf.n10 por_dig_0.por_unbuf.n9 10.4965
R29794 por_dig_0.por_unbuf por_dig_0.por_unbuf.n28 7.02042
R29795 por_dig_0.por_unbuf.n10 por_dig_0.por_unbuf 6.6565
R29796 por_dig_0.por_unbuf.n6 por_dig_0.por_unbuf 6.4005
R29797 por_dig_0.por_unbuf.n9 por_dig_0.por_unbuf 6.4005
R29798 por_dig_0.por_unbuf.n17 por_dig_0.por_unbuf 6.4005
R29799 por_dig_0.por_unbuf.n20 por_dig_0.por_unbuf 6.4005
R29800 por_dig_0.por_unbuf.n26 por_dig_0.por_unbuf.n25 5.9876
R29801 por_dig_0.por_unbuf.n28 por_dig_0.por_unbuf 5.54059
R29802 por_dig_0.por_unbuf.n31 por_dig_0.por_unbuf 5.27109
R29803 por_dig_0.por_unbuf.n25 por_dig_0.por_unbuf 4.74889
R29804 por_dig_0.por_unbuf.n21 por_dig_0.por_unbuf.n20 4.6085
R29805 por_dig_0.por_unbuf.n26 por_dig_0.por_unbuf 4.54244
R29806 por_dig_0.por_unbuf por_dig_0.por_unbuf.n5 4.3525
R29807 por_dig_0.por_unbuf por_dig_0.por_unbuf.n16 4.3525
R29808 por_dig_0.por_unbuf por_dig_0.por_unbuf.n29 4.26717
R29809 por_dig_0.por_unbuf.n33 por_dig_0.por_unbuf 1.50638
R29810 isrc_sel.n0 isrc_sel.t3 186.374
R29811 isrc_sel.n0 isrc_sel.t2 170.308
R29812 isrc_sel.n1 isrc_sel 154.56
R29813 isrc_sel.n2 isrc_sel.n1 153.462
R29814 isrc_sel.n1 isrc_sel.n0 101.513
R29815 isrc_sel.n5 isrc_sel.n4 79.0476
R29816 isrc_sel.n4 isrc_sel.t1 16.5305
R29817 isrc_sel.n4 isrc_sel.t0 16.5305
R29818 isrc_sel.n6 isrc_sel.n3 11.611
R29819 isrc_sel.n6 isrc_sel.n5 6.24886
R29820 isrc_sel.n3 isrc_sel.n2 4.96991
R29821 isrc_sel.n2 isrc_sel 3.46403
R29822 isrc_sel.n3 isrc_sel 2.71109
R29823 isrc_sel.n5 isrc_sel 0.710641
R29824 isrc_sel isrc_sel.n6 0.189953
R29825 por_ana_0.rstring_mux_0.vtop.n4 por_ana_0.rstring_mux_0.vtop.t16 87.3599
R29826 por_ana_0.rstring_mux_0.vtop.n2 por_ana_0.rstring_mux_0.vtop.n0 48.5415
R29827 por_ana_0.rstring_mux_0.vtop.n13 por_ana_0.rstring_mux_0.vtop.n12 48.4284
R29828 por_ana_0.rstring_mux_0.vtop.n11 por_ana_0.rstring_mux_0.vtop.n10 48.4284
R29829 por_ana_0.rstring_mux_0.vtop.n9 por_ana_0.rstring_mux_0.vtop.n8 48.4284
R29830 por_ana_0.rstring_mux_0.vtop.n7 por_ana_0.rstring_mux_0.vtop.n6 48.4284
R29831 por_ana_0.rstring_mux_0.vtop.n2 por_ana_0.rstring_mux_0.vtop.n1 48.4284
R29832 por_ana_0.rstring_mux_0.vtop.n15 por_ana_0.rstring_mux_0.vtop.n14 45.0184
R29833 por_ana_0.rstring_mux_0.vtop.n4 por_ana_0.rstring_mux_0.vtop.n3 45.0184
R29834 por_ana_0.rstring_mux_0.vtop por_ana_0.rstring_mux_0.vtop.t17 19.1879
R29835 por_ana_0.rstring_mux_0.vtop.n14 por_ana_0.rstring_mux_0.vtop.t1 5.5395
R29836 por_ana_0.rstring_mux_0.vtop.n14 por_ana_0.rstring_mux_0.vtop.t14 5.5395
R29837 por_ana_0.rstring_mux_0.vtop.n12 por_ana_0.rstring_mux_0.vtop.t8 5.5395
R29838 por_ana_0.rstring_mux_0.vtop.n12 por_ana_0.rstring_mux_0.vtop.t7 5.5395
R29839 por_ana_0.rstring_mux_0.vtop.n10 por_ana_0.rstring_mux_0.vtop.t9 5.5395
R29840 por_ana_0.rstring_mux_0.vtop.n10 por_ana_0.rstring_mux_0.vtop.t12 5.5395
R29841 por_ana_0.rstring_mux_0.vtop.n8 por_ana_0.rstring_mux_0.vtop.t3 5.5395
R29842 por_ana_0.rstring_mux_0.vtop.n8 por_ana_0.rstring_mux_0.vtop.t10 5.5395
R29843 por_ana_0.rstring_mux_0.vtop.n6 por_ana_0.rstring_mux_0.vtop.t6 5.5395
R29844 por_ana_0.rstring_mux_0.vtop.n6 por_ana_0.rstring_mux_0.vtop.t4 5.5395
R29845 por_ana_0.rstring_mux_0.vtop.n3 por_ana_0.rstring_mux_0.vtop.t11 5.5395
R29846 por_ana_0.rstring_mux_0.vtop.n3 por_ana_0.rstring_mux_0.vtop.t5 5.5395
R29847 por_ana_0.rstring_mux_0.vtop.n1 por_ana_0.rstring_mux_0.vtop.t15 5.5395
R29848 por_ana_0.rstring_mux_0.vtop.n1 por_ana_0.rstring_mux_0.vtop.t13 5.5395
R29849 por_ana_0.rstring_mux_0.vtop.n0 por_ana_0.rstring_mux_0.vtop.t0 5.5395
R29850 por_ana_0.rstring_mux_0.vtop.n0 por_ana_0.rstring_mux_0.vtop.t2 5.5395
R29851 por_ana_0.rstring_mux_0.vtop.n15 por_ana_0.rstring_mux_0.vtop.n13 3.5118
R29852 por_ana_0.rstring_mux_0.vtop.n5 por_ana_0.rstring_mux_0.vtop.n4 3.4105
R29853 por_ana_0.rstring_mux_0.vtop por_ana_0.rstring_mux_0.vtop.n15 0.829892
R29854 por_ana_0.rstring_mux_0.vtop.n5 por_ana_0.rstring_mux_0.vtop.n2 0.113554
R29855 por_ana_0.rstring_mux_0.vtop.n7 por_ana_0.rstring_mux_0.vtop.n5 0.113554
R29856 por_ana_0.rstring_mux_0.vtop.n9 por_ana_0.rstring_mux_0.vtop.n7 0.113554
R29857 por_ana_0.rstring_mux_0.vtop.n11 por_ana_0.rstring_mux_0.vtop.n9 0.113554
R29858 por_ana_0.rstring_mux_0.vtop.n13 por_ana_0.rstring_mux_0.vtop.n11 0.113554
R29859 por_dig_0.clknet_0_osc_ck.n34 por_dig_0.clknet_0_osc_ck.n32 333.392
R29860 por_dig_0.clknet_0_osc_ck.n38 por_dig_0.clknet_0_osc_ck.n28 301.392
R29861 por_dig_0.clknet_0_osc_ck.n37 por_dig_0.clknet_0_osc_ck.n29 301.392
R29862 por_dig_0.clknet_0_osc_ck.n36 por_dig_0.clknet_0_osc_ck.n30 301.392
R29863 por_dig_0.clknet_0_osc_ck.n35 por_dig_0.clknet_0_osc_ck.n31 301.392
R29864 por_dig_0.clknet_0_osc_ck.n34 por_dig_0.clknet_0_osc_ck.n33 301.392
R29865 por_dig_0.clknet_0_osc_ck por_dig_0.clknet_0_osc_ck.n40 297.752
R29866 por_dig_0.clknet_0_osc_ck.n27 por_dig_0.clknet_0_osc_ck.n26 287.303
R29867 por_dig_0.clknet_0_osc_ck.n2 por_dig_0.clknet_0_osc_ck.n0 248.638
R29868 por_dig_0.clknet_0_osc_ck.n2 por_dig_0.clknet_0_osc_ck.n1 203.463
R29869 por_dig_0.clknet_0_osc_ck.n4 por_dig_0.clknet_0_osc_ck.n3 203.463
R29870 por_dig_0.clknet_0_osc_ck.n8 por_dig_0.clknet_0_osc_ck.n7 203.463
R29871 por_dig_0.clknet_0_osc_ck.n10 por_dig_0.clknet_0_osc_ck.n9 203.463
R29872 por_dig_0.clknet_0_osc_ck.n12 por_dig_0.clknet_0_osc_ck.n11 203.463
R29873 por_dig_0.clknet_0_osc_ck.n6 por_dig_0.clknet_0_osc_ck.n5 202.456
R29874 por_dig_0.clknet_0_osc_ck.n14 por_dig_0.clknet_0_osc_ck.n13 200.212
R29875 por_dig_0.clknet_0_osc_ck.n15 por_dig_0.clknet_0_osc_ck.t42 184.768
R29876 por_dig_0.clknet_0_osc_ck.n16 por_dig_0.clknet_0_osc_ck.t35 184.768
R29877 por_dig_0.clknet_0_osc_ck.n17 por_dig_0.clknet_0_osc_ck.t46 184.768
R29878 por_dig_0.clknet_0_osc_ck.n18 por_dig_0.clknet_0_osc_ck.t36 184.768
R29879 por_dig_0.clknet_0_osc_ck.n23 por_dig_0.clknet_0_osc_ck.t44 184.768
R29880 por_dig_0.clknet_0_osc_ck.n22 por_dig_0.clknet_0_osc_ck.t38 184.768
R29881 por_dig_0.clknet_0_osc_ck.n21 por_dig_0.clknet_0_osc_ck.t33 184.768
R29882 por_dig_0.clknet_0_osc_ck.n20 por_dig_0.clknet_0_osc_ck.t40 184.768
R29883 por_dig_0.clknet_0_osc_ck por_dig_0.clknet_0_osc_ck.n18 173.609
R29884 por_dig_0.clknet_0_osc_ck.n24 por_dig_0.clknet_0_osc_ck.n23 171.375
R29885 por_dig_0.clknet_0_osc_ck.n15 por_dig_0.clknet_0_osc_ck.t45 146.208
R29886 por_dig_0.clknet_0_osc_ck.n16 por_dig_0.clknet_0_osc_ck.t39 146.208
R29887 por_dig_0.clknet_0_osc_ck.n17 por_dig_0.clknet_0_osc_ck.t34 146.208
R29888 por_dig_0.clknet_0_osc_ck.n18 por_dig_0.clknet_0_osc_ck.t41 146.208
R29889 por_dig_0.clknet_0_osc_ck.n23 por_dig_0.clknet_0_osc_ck.t37 146.208
R29890 por_dig_0.clknet_0_osc_ck.n22 por_dig_0.clknet_0_osc_ck.t47 146.208
R29891 por_dig_0.clknet_0_osc_ck.n21 por_dig_0.clknet_0_osc_ck.t43 146.208
R29892 por_dig_0.clknet_0_osc_ck.n20 por_dig_0.clknet_0_osc_ck.t32 146.208
R29893 por_dig_0.clknet_0_osc_ck.n4 por_dig_0.clknet_0_osc_ck.n2 45.177
R29894 por_dig_0.clknet_0_osc_ck.n10 por_dig_0.clknet_0_osc_ck.n8 45.177
R29895 por_dig_0.clknet_0_osc_ck.n12 por_dig_0.clknet_0_osc_ck.n10 45.177
R29896 por_dig_0.clknet_0_osc_ck.n6 por_dig_0.clknet_0_osc_ck.n4 44.0476
R29897 por_dig_0.clknet_0_osc_ck.n8 por_dig_0.clknet_0_osc_ck.n6 44.0476
R29898 por_dig_0.clknet_0_osc_ck.n16 por_dig_0.clknet_0_osc_ck.n15 40.6397
R29899 por_dig_0.clknet_0_osc_ck.n17 por_dig_0.clknet_0_osc_ck.n16 40.6397
R29900 por_dig_0.clknet_0_osc_ck.n18 por_dig_0.clknet_0_osc_ck.n17 40.6397
R29901 por_dig_0.clknet_0_osc_ck.n23 por_dig_0.clknet_0_osc_ck.n22 40.6397
R29902 por_dig_0.clknet_0_osc_ck.n22 por_dig_0.clknet_0_osc_ck.n21 40.6397
R29903 por_dig_0.clknet_0_osc_ck.n21 por_dig_0.clknet_0_osc_ck.n20 40.6397
R29904 por_dig_0.clknet_0_osc_ck.n0 por_dig_0.clknet_0_osc_ck.t1 40.0005
R29905 por_dig_0.clknet_0_osc_ck.n0 por_dig_0.clknet_0_osc_ck.t4 40.0005
R29906 por_dig_0.clknet_0_osc_ck.n1 por_dig_0.clknet_0_osc_ck.t2 40.0005
R29907 por_dig_0.clknet_0_osc_ck.n1 por_dig_0.clknet_0_osc_ck.t11 40.0005
R29908 por_dig_0.clknet_0_osc_ck.n3 por_dig_0.clknet_0_osc_ck.t8 40.0005
R29909 por_dig_0.clknet_0_osc_ck.n3 por_dig_0.clknet_0_osc_ck.t14 40.0005
R29910 por_dig_0.clknet_0_osc_ck.n5 por_dig_0.clknet_0_osc_ck.t9 40.0005
R29911 por_dig_0.clknet_0_osc_ck.n5 por_dig_0.clknet_0_osc_ck.t15 40.0005
R29912 por_dig_0.clknet_0_osc_ck.n7 por_dig_0.clknet_0_osc_ck.t10 40.0005
R29913 por_dig_0.clknet_0_osc_ck.n7 por_dig_0.clknet_0_osc_ck.t0 40.0005
R29914 por_dig_0.clknet_0_osc_ck.n9 por_dig_0.clknet_0_osc_ck.t12 40.0005
R29915 por_dig_0.clknet_0_osc_ck.n9 por_dig_0.clknet_0_osc_ck.t3 40.0005
R29916 por_dig_0.clknet_0_osc_ck.n11 por_dig_0.clknet_0_osc_ck.t13 40.0005
R29917 por_dig_0.clknet_0_osc_ck.n11 por_dig_0.clknet_0_osc_ck.t5 40.0005
R29918 por_dig_0.clknet_0_osc_ck.n13 por_dig_0.clknet_0_osc_ck.t6 40.0005
R29919 por_dig_0.clknet_0_osc_ck.n13 por_dig_0.clknet_0_osc_ck.t7 40.0005
R29920 por_dig_0.clknet_0_osc_ck.n39 por_dig_0.clknet_0_osc_ck.n38 32.0005
R29921 por_dig_0.clknet_0_osc_ck.n38 por_dig_0.clknet_0_osc_ck.n37 32.0005
R29922 por_dig_0.clknet_0_osc_ck.n36 por_dig_0.clknet_0_osc_ck.n35 32.0005
R29923 por_dig_0.clknet_0_osc_ck.n35 por_dig_0.clknet_0_osc_ck.n34 32.0005
R29924 por_dig_0.clknet_0_osc_ck.n37 por_dig_0.clknet_0_osc_ck.n36 31.2005
R29925 por_dig_0.clknet_0_osc_ck.n27 por_dig_0.clknet_0_osc_ck.n25 28.6283
R29926 por_dig_0.clknet_0_osc_ck.n26 por_dig_0.clknet_0_osc_ck.t26 27.5805
R29927 por_dig_0.clknet_0_osc_ck.n26 por_dig_0.clknet_0_osc_ck.t18 27.5805
R29928 por_dig_0.clknet_0_osc_ck.n40 por_dig_0.clknet_0_osc_ck.t19 27.5805
R29929 por_dig_0.clknet_0_osc_ck.n40 por_dig_0.clknet_0_osc_ck.t20 27.5805
R29930 por_dig_0.clknet_0_osc_ck.n28 por_dig_0.clknet_0_osc_ck.t25 27.5805
R29931 por_dig_0.clknet_0_osc_ck.n28 por_dig_0.clknet_0_osc_ck.t16 27.5805
R29932 por_dig_0.clknet_0_osc_ck.n29 por_dig_0.clknet_0_osc_ck.t23 27.5805
R29933 por_dig_0.clknet_0_osc_ck.n29 por_dig_0.clknet_0_osc_ck.t29 27.5805
R29934 por_dig_0.clknet_0_osc_ck.n30 por_dig_0.clknet_0_osc_ck.t22 27.5805
R29935 por_dig_0.clknet_0_osc_ck.n30 por_dig_0.clknet_0_osc_ck.t28 27.5805
R29936 por_dig_0.clknet_0_osc_ck.n31 por_dig_0.clknet_0_osc_ck.t21 27.5805
R29937 por_dig_0.clknet_0_osc_ck.n31 por_dig_0.clknet_0_osc_ck.t27 27.5805
R29938 por_dig_0.clknet_0_osc_ck.n32 por_dig_0.clknet_0_osc_ck.t30 27.5805
R29939 por_dig_0.clknet_0_osc_ck.n32 por_dig_0.clknet_0_osc_ck.t17 27.5805
R29940 por_dig_0.clknet_0_osc_ck.n33 por_dig_0.clknet_0_osc_ck.t31 27.5805
R29941 por_dig_0.clknet_0_osc_ck.n33 por_dig_0.clknet_0_osc_ck.t24 27.5805
R29942 por_dig_0.clknet_0_osc_ck.n25 por_dig_0.clknet_0_osc_ck.n19 22.3735
R29943 por_dig_0.clknet_0_osc_ck.n39 por_dig_0.clknet_0_osc_ck.n27 14.0898
R29944 por_dig_0.clknet_0_osc_ck.n14 por_dig_0.clknet_0_osc_ck.n12 13.177
R29945 por_dig_0.clknet_0_osc_ck.n19 por_dig_0.clknet_0_osc_ck 10.3624
R29946 por_dig_0.clknet_0_osc_ck por_dig_0.clknet_0_osc_ck.n39 10.2022
R29947 por_dig_0.clknet_0_osc_ck por_dig_0.clknet_0_osc_ck.n24 9.14336
R29948 por_dig_0.clknet_0_osc_ck.n24 por_dig_0.clknet_0_osc_ck 4.67352
R29949 por_dig_0.clknet_0_osc_ck.n25 por_dig_0.clknet_0_osc_ck 4.18457
R29950 por_dig_0.clknet_0_osc_ck.n19 por_dig_0.clknet_0_osc_ck 3.45447
R29951 por_dig_0.clknet_0_osc_ck por_dig_0.clknet_0_osc_ck.n14 1.26402
R29952 por_dig_0.net5.t12 por_dig_0.net5.t4 403.274
R29953 por_dig_0.net5.n1 por_dig_0.net5.t10 323.55
R29954 por_dig_0.net5.n0 por_dig_0.net5.t1 319.171
R29955 por_dig_0.net5.n12 por_dig_0.net5.t12 306.14
R29956 por_dig_0.net5.n16 por_dig_0.net5.t5 241.536
R29957 por_dig_0.net5.n20 por_dig_0.net5.t19 241.536
R29958 por_dig_0.net5.n7 por_dig_0.net5.t9 231.017
R29959 por_dig_0.net5 por_dig_0.net5.t0 209.923
R29960 por_dig_0.net5.n4 por_dig_0.net5.t6 204.656
R29961 por_dig_0.net5.n22 por_dig_0.net5.t15 201.369
R29962 por_dig_0.net5.n11 por_dig_0.net5.t11 196.549
R29963 por_dig_0.net5.n1 por_dig_0.net5.t7 195.017
R29964 por_dig_0.net5.n9 por_dig_0.net5.t18 173.34
R29965 por_dig_0.net5.n16 por_dig_0.net5.t14 169.237
R29966 por_dig_0.net5.n20 por_dig_0.net5.t8 169.237
R29967 por_dig_0.net5.n10 por_dig_0.net5.n9 162.862
R29968 por_dig_0.net5.n9 por_dig_0.net5.t3 162.81
R29969 por_dig_0.net5 por_dig_0.net5.n11 159.024
R29970 por_dig_0.net5.n7 por_dig_0.net5.t17 158.716
R29971 por_dig_0.net5 por_dig_0.net5.n20 158.133
R29972 por_dig_0.net5 por_dig_0.net5.n1 153.409
R29973 por_dig_0.net5.n6 por_dig_0.net5.n3 153.13
R29974 por_dig_0.net5.n23 por_dig_0.net5.n22 152.827
R29975 por_dig_0.net5.n17 por_dig_0.net5.n16 152
R29976 por_dig_0.net5.n8 por_dig_0.net5.n7 152
R29977 por_dig_0.net5.n5 por_dig_0.net5.n4 152
R29978 por_dig_0.net5.n11 por_dig_0.net5.t13 148.35
R29979 por_dig_0.net5.n22 por_dig_0.net5.t16 132.282
R29980 por_dig_0.net5.n3 por_dig_0.net5.t2 121.109
R29981 por_dig_0.net5.n4 por_dig_0.net5.n3 40.9982
R29982 por_dig_0.net5.n21 por_dig_0.net5 23.1946
R29983 por_dig_0.net5 por_dig_0.net5.n26 16.7116
R29984 por_dig_0.net5.n26 por_dig_0.net5 16.0005
R29985 por_dig_0.net5.n19 por_dig_0.net5.n18 14.9842
R29986 por_dig_0.net5.n25 por_dig_0.net5.n24 14.5232
R29987 por_dig_0.net5.n19 por_dig_0.net5.n6 13.291
R29988 por_dig_0.net5.n13 por_dig_0.net5.n12 12.7357
R29989 por_dig_0.net5.n13 por_dig_0.net5 11.9542
R29990 por_dig_0.net5.n24 por_dig_0.net5.n21 11.2972
R29991 por_dig_0.net5.n15 por_dig_0.net5.n8 10.6521
R29992 por_dig_0.net5 por_dig_0.net5.n5 9.6005
R29993 por_dig_0.net5 por_dig_0.net5.n10 9.49091
R29994 por_dig_0.net5.n18 por_dig_0.net5.n17 9.3005
R29995 por_dig_0.net5.n24 por_dig_0.net5.n23 9.3005
R29996 por_dig_0.net5.n14 por_dig_0.net5 8.00812
R29997 por_dig_0.net5.n15 por_dig_0.net5.n14 7.73961
R29998 por_dig_0.net5 por_dig_0.net5.n0 7.73474
R29999 por_dig_0.net5 por_dig_0.net5.n2 6.34564
R30000 por_dig_0.net5.n26 por_dig_0.net5 5.7605
R30001 por_dig_0.net5.n14 por_dig_0.net5.n13 4.5005
R30002 por_dig_0.net5.n18 por_dig_0.net5.n15 4.24604
R30003 por_dig_0.net5.n12 por_dig_0.net5 3.2005
R30004 por_dig_0.net5.n6 por_dig_0.net5 3.2005
R30005 por_dig_0.net5.n5 por_dig_0.net5 3.2005
R30006 por_dig_0.net5.n26 por_dig_0.net5.n25 3.2005
R30007 por_dig_0.net5.n25 por_dig_0.net5 2.8165
R30008 por_dig_0.net5.n21 por_dig_0.net5.n19 2.52385
R30009 por_dig_0.net5.n0 por_dig_0.net5 2.48634
R30010 por_dig_0.net5.n10 por_dig_0.net5 2.32777
R30011 por_dig_0.net5.n8 por_dig_0.net5 2.32777
R30012 por_dig_0.net5.n2 por_dig_0.net5 2.19479
R30013 por_dig_0.net5.n2 por_dig_0.net5 1.80756
R30014 por_dig_0.net5.n23 por_dig_0.net5 1.75534
R30015 por_dig_0.net5.n17 por_dig_0.net5 1.75534
R30016 vin.n94 vin.n93 74.2619
R30017 vin.n92 vin.n60 60.2207
R30018 vin.n59 vin.t22 53.91
R30019 vin.n56 vin.n55 48.371
R30020 vin.n52 vin.n51 48.371
R30021 vin.n48 vin.n8 48.371
R30022 vin.n45 vin.n44 48.371
R30023 vin.n41 vin.n40 48.371
R30024 vin.n37 vin.n21 48.371
R30025 vin.n34 vin.n19 48.371
R30026 vin.n58 vin.n57 45.4885
R30027 vin.n54 vin.n53 45.4885
R30028 vin.n7 vin.n5 45.4885
R30029 vin.n47 vin.n46 45.4885
R30030 vin.n43 vin.n42 45.4885
R30031 vin.n20 vin.n18 45.4885
R30032 vin.n36 vin.n35 45.4885
R30033 vin.n28 vin.n27 45.4885
R30034 vin.n1 vin.t35 21.0726
R30035 vin.n4 vin.n3 17.7666
R30036 vin.n11 vin.n10 17.7666
R30037 vin.n14 vin.n13 17.7666
R30038 vin.n17 vin.n16 17.7666
R30039 vin.n24 vin.n23 17.7666
R30040 vin.n33 vin.n26 17.7666
R30041 vin.n31 vin.n30 17.7666
R30042 vin.n2 vin.n1 16.9742
R30043 vin.n9 vin.n4 16.9742
R30044 vin.n12 vin.n11 16.9742
R30045 vin.n15 vin.n14 16.9742
R30046 vin.n22 vin.n17 16.9742
R30047 vin.n25 vin.n24 16.9742
R30048 vin.n33 vin.n32 16.9742
R30049 vin.n30 vin.n29 16.9742
R30050 vin.n93 vin.t39 16.5305
R30051 vin.n93 vin.t38 16.5305
R30052 vin.n90 vin.t53 14.8978
R30053 vin.n89 vin.t53 14.8978
R30054 vin.n86 vin.t62 14.8978
R30055 vin.n85 vin.t62 14.8978
R30056 vin.n82 vin.t54 14.8978
R30057 vin.n81 vin.t54 14.8978
R30058 vin.n78 vin.t57 14.8978
R30059 vin.n77 vin.t57 14.8978
R30060 vin.n74 vin.t55 14.8978
R30061 vin.n73 vin.t55 14.8978
R30062 vin.n70 vin.t63 14.8978
R30063 vin.n69 vin.t63 14.8978
R30064 vin.n66 vin.t56 14.8978
R30065 vin.n65 vin.t56 14.8978
R30066 vin.n62 vin.t64 14.8978
R30067 vin.t64 vin.n61 14.8978
R30068 vin.t58 vin.n89 12.9902
R30069 vin.n90 vin.t58 12.9902
R30070 vin.t50 vin.n85 12.9902
R30071 vin.n86 vin.t50 12.9902
R30072 vin.t59 vin.n81 12.9902
R30073 vin.n82 vin.t59 12.9902
R30074 vin.t65 vin.n77 12.9902
R30075 vin.n78 vin.t65 12.9902
R30076 vin.t60 vin.n73 12.9902
R30077 vin.n74 vin.t60 12.9902
R30078 vin.t51 vin.n69 12.9902
R30079 vin.n70 vin.t51 12.9902
R30080 vin.t61 vin.n65 12.9902
R30081 vin.n66 vin.t61 12.9902
R30082 vin.t52 vin.n61 12.9902
R30083 vin.n62 vin.t52 12.9902
R30084 vin.n94 vin.n92 6.26717
R30085 vin.n92 vin.n91 6.1004
R30086 vin.n57 vin.t4 5.5395
R30087 vin.n57 vin.t23 5.5395
R30088 vin.n53 vin.t6 5.5395
R30089 vin.n53 vin.t11 5.5395
R30090 vin.n56 vin.t10 5.5395
R30091 vin.t4 vin.n56 5.5395
R30092 vin.t3 vin.n7 5.5395
R30093 vin.n7 vin.t36 5.5395
R30094 vin.n52 vin.t37 5.5395
R30095 vin.t6 vin.n52 5.5395
R30096 vin.n46 vin.t7 5.5395
R30097 vin.n46 vin.t28 5.5395
R30098 vin.n8 vin.t29 5.5395
R30099 vin.n8 vin.t3 5.5395
R30100 vin.n42 vin.t9 5.5395
R30101 vin.n42 vin.t41 5.5395
R30102 vin.n45 vin.t40 5.5395
R30103 vin.t7 vin.n45 5.5395
R30104 vin.t5 vin.n20 5.5395
R30105 vin.n20 vin.t33 5.5395
R30106 vin.n41 vin.t32 5.5395
R30107 vin.t9 vin.n41 5.5395
R30108 vin.n35 vin.t8 5.5395
R30109 vin.n35 vin.t45 5.5395
R30110 vin.n21 vin.t44 5.5395
R30111 vin.n21 vin.t5 5.5395
R30112 vin.n27 vin.t2 5.5395
R30113 vin.n27 vin.t48 5.5395
R30114 vin.n34 vin.t49 5.5395
R30115 vin.t8 vin.n34 5.5395
R30116 vin.n63 vin.n61 5.24569
R30117 vin.n63 vin.n62 4.5005
R30118 vin.n65 vin.n64 4.5005
R30119 vin.n67 vin.n66 4.5005
R30120 vin.n69 vin.n68 4.5005
R30121 vin.n71 vin.n70 4.5005
R30122 vin.n73 vin.n72 4.5005
R30123 vin.n75 vin.n74 4.5005
R30124 vin.n77 vin.n76 4.5005
R30125 vin.n79 vin.n78 4.5005
R30126 vin.n81 vin.n80 4.5005
R30127 vin.n83 vin.n82 4.5005
R30128 vin.n85 vin.n84 4.5005
R30129 vin.n87 vin.n86 4.5005
R30130 vin.n89 vin.n88 4.5005
R30131 vin.n91 vin.n90 4.5005
R30132 vin.n38 vin.n19 3.79433
R30133 vin.n38 vin.n37 3.4105
R30134 vin.n40 vin.n39 3.4105
R30135 vin.n44 vin.n6 3.4105
R30136 vin.n49 vin.n48 3.4105
R30137 vin.n51 vin.n50 3.4105
R30138 vin.n55 vin.n0 3.4105
R30139 vin.n60 vin.n59 3.4105
R30140 vin.t16 vin.n2 3.3065
R30141 vin.n2 vin.t34 3.3065
R30142 vin.t18 vin.n9 3.3065
R30143 vin.n9 vin.t13 3.3065
R30144 vin.n3 vin.t12 3.3065
R30145 vin.n3 vin.t16 3.3065
R30146 vin.t15 vin.n12 3.3065
R30147 vin.n12 vin.t0 3.3065
R30148 vin.n10 vin.t1 3.3065
R30149 vin.n10 vin.t18 3.3065
R30150 vin.t19 vin.n15 3.3065
R30151 vin.n15 vin.t26 3.3065
R30152 vin.n13 vin.t27 3.3065
R30153 vin.n13 vin.t15 3.3065
R30154 vin.t21 vin.n22 3.3065
R30155 vin.n22 vin.t47 3.3065
R30156 vin.n16 vin.t46 3.3065
R30157 vin.n16 vin.t19 3.3065
R30158 vin.t17 vin.n25 3.3065
R30159 vin.n25 vin.t31 3.3065
R30160 vin.n23 vin.t30 3.3065
R30161 vin.n23 vin.t21 3.3065
R30162 vin.n32 vin.t20 3.3065
R30163 vin.n32 vin.t43 3.3065
R30164 vin.n26 vin.t42 3.3065
R30165 vin.n26 vin.t17 3.3065
R30166 vin.n29 vin.t14 3.3065
R30167 vin.n29 vin.t24 3.3065
R30168 vin.n31 vin.t25 3.3065
R30169 vin.t20 vin.n31 3.3065
R30170 vin.n58 vin.n1 1.98319
R30171 vin.n54 vin.n4 1.98319
R30172 vin.n11 vin.n5 1.98319
R30173 vin.n47 vin.n14 1.98319
R30174 vin.n43 vin.n17 1.98319
R30175 vin.n24 vin.n18 1.98319
R30176 vin.n36 vin.n33 1.98319
R30177 vin.n30 vin.n28 1.98319
R30178 vin vin.n94 0.943633
R30179 vin.n91 vin.n88 0.745692
R30180 vin.n87 vin.n84 0.745692
R30181 vin.n83 vin.n80 0.745692
R30182 vin.n79 vin.n76 0.745692
R30183 vin.n75 vin.n72 0.745692
R30184 vin.n71 vin.n68 0.745692
R30185 vin.n67 vin.n64 0.745692
R30186 vin.n39 vin.n38 0.384333
R30187 vin.n39 vin.n6 0.384333
R30188 vin.n49 vin.n6 0.384333
R30189 vin.n50 vin.n49 0.384333
R30190 vin.n50 vin.n0 0.384333
R30191 vin.n60 vin.n0 0.384333
R30192 vin.n88 vin.n87 0.260115
R30193 vin.n84 vin.n83 0.260115
R30194 vin.n80 vin.n79 0.260115
R30195 vin.n76 vin.n75 0.260115
R30196 vin.n72 vin.n71 0.260115
R30197 vin.n68 vin.n67 0.260115
R30198 vin.n64 vin.n63 0.260115
R30199 vin.n59 vin.n58 0.00218919
R30200 vin.n55 vin.n54 0.00218919
R30201 vin.n51 vin.n5 0.00218919
R30202 vin.n48 vin.n47 0.00218919
R30203 vin.n44 vin.n43 0.00218919
R30204 vin.n40 vin.n18 0.00218919
R30205 vin.n37 vin.n36 0.00218919
R30206 vin.n28 vin.n19 0.00218919
R30207 por_ana_0.ibias_gen_0.vstart.n0 por_ana_0.ibias_gen_0.vstart.t10 56.685
R30208 por_ana_0.ibias_gen_0.vstart.n6 por_ana_0.ibias_gen_0.vstart.n5 20.328
R30209 por_ana_0.ibias_gen_0.vstart.n0 por_ana_0.ibias_gen_0.vstart.n1 20.2356
R30210 por_ana_0.ibias_gen_0.vstart.n4 por_ana_0.ibias_gen_0.vstart.n3 20.069
R30211 por_ana_0.ibias_gen_0.vstart.n0 por_ana_0.ibias_gen_0.vstart.n2 20.069
R30212 por_ana_0.ibias_gen_0.vstart.n7 por_ana_0.ibias_gen_0.vstart.n6 20.069
R30213 por_ana_0.ibias_gen_0.vstart.n5 por_ana_0.ibias_gen_0.vstart.t7 3.3065
R30214 por_ana_0.ibias_gen_0.vstart.n5 por_ana_0.ibias_gen_0.vstart.t1 3.3065
R30215 por_ana_0.ibias_gen_0.vstart.n3 por_ana_0.ibias_gen_0.vstart.t0 3.3065
R30216 por_ana_0.ibias_gen_0.vstart.n3 por_ana_0.ibias_gen_0.vstart.t8 3.3065
R30217 por_ana_0.ibias_gen_0.vstart.n2 por_ana_0.ibias_gen_0.vstart.t5 3.3065
R30218 por_ana_0.ibias_gen_0.vstart.n2 por_ana_0.ibias_gen_0.vstart.t3 3.3065
R30219 por_ana_0.ibias_gen_0.vstart.n1 por_ana_0.ibias_gen_0.vstart.t4 3.3065
R30220 por_ana_0.ibias_gen_0.vstart.n1 por_ana_0.ibias_gen_0.vstart.t2 3.3065
R30221 por_ana_0.ibias_gen_0.vstart.n7 por_ana_0.ibias_gen_0.vstart.t6 3.3065
R30222 por_ana_0.ibias_gen_0.vstart.t9 por_ana_0.ibias_gen_0.vstart.n7 3.3065
R30223 por_ana_0.ibias_gen_0.vstart.n4 por_ana_0.ibias_gen_0.vstart.n0 0.280933
R30224 por_ana_0.ibias_gen_0.vstart.n6 por_ana_0.ibias_gen_0.vstart.n4 0.2449
R30225 por_timed_out.n2 por_timed_out 589.769
R30226 por_timed_out.n3 por_timed_out.n2 585
R30227 por_timed_out.n1 por_timed_out.n0 185
R30228 por_timed_out por_timed_out.n1 81.3181
R30229 por_timed_out.n2 por_timed_out.t3 26.5955
R30230 por_timed_out.n2 por_timed_out.t2 26.5955
R30231 por_timed_out.n0 por_timed_out.t1 24.9236
R30232 por_timed_out.n0 por_timed_out.t0 24.9236
R30233 por_timed_out por_timed_out.n4 17.6146
R30234 por_timed_out.n4 por_timed_out 12.8005
R30235 por_timed_out.n1 por_timed_out 5.27109
R30236 por_timed_out.n4 por_timed_out.n3 2.76128
R30237 por_timed_out.n3 por_timed_out 1.50638
R30238 otrip[2].n0 otrip[2].t2 323.55
R30239 otrip[2].n0 otrip[2].t3 195.017
R30240 otrip[2].n1 otrip[2].n0 152
R30241 otrip[2].n4 otrip[2].n3 74.6239
R30242 otrip[2] otrip[2].n2 17.7709
R30243 otrip[2].n3 otrip[2].t0 16.5305
R30244 otrip[2].n3 otrip[2].t1 16.5305
R30245 otrip[2].n5 otrip[2].n4 9.66698
R30246 otrip[2].n2 otrip[2] 6.7304
R30247 otrip[2] otrip[2].n5 4.05854
R30248 otrip[2].n1 otrip[2] 1.45205
R30249 otrip[2].n5 otrip[2] 1.02282
R30250 otrip[2].n2 otrip[2].n1 0.792253
R30251 otrip[2].n4 otrip[2] 0.7431
R30252 por_ana_0.comparator_1.vnn.n7 por_ana_0.comparator_1.vnn.t46 244.34
R30253 por_ana_0.comparator_1.vnn.n7 por_ana_0.comparator_1.vnn.n21 204.284
R30254 por_ana_0.comparator_1.vnn.n7 por_ana_0.comparator_1.vnn.n22 204.284
R30255 por_ana_0.comparator_1.vnn.n7 por_ana_0.comparator_1.vnn.n23 204.284
R30256 por_ana_0.comparator_1.vnn.n7 por_ana_0.comparator_1.vnn.n24 204.284
R30257 por_ana_0.comparator_1.vnn.n7 por_ana_0.comparator_1.vnn.n25 204.284
R30258 por_ana_0.comparator_1.vnn.n7 por_ana_0.comparator_1.vnn.n26 204.284
R30259 por_ana_0.comparator_1.vnn.n7 por_ana_0.comparator_1.vnn.n20 204.284
R30260 por_ana_0.comparator_1.vnn.n6 por_ana_0.comparator_1.vnn.n17 199.784
R30261 por_ana_0.comparator_1.vnn.n6 por_ana_0.comparator_1.vnn.n16 199.65
R30262 por_ana_0.comparator_1.vnn.n6 por_ana_0.comparator_1.vnn.n18 199.65
R30263 por_ana_0.comparator_1.vnn.n6 por_ana_0.comparator_1.vnn.n19 199.65
R30264 por_ana_0.comparator_1.vnn.n0 por_ana_0.comparator_1.vnn.n8 71.9371
R30265 por_ana_0.comparator_1.vnn.n0 por_ana_0.comparator_1.vnn.n15 70.9612
R30266 por_ana_0.comparator_1.vnn.n0 por_ana_0.comparator_1.vnn.n14 70.9612
R30267 por_ana_0.comparator_1.vnn.n0 por_ana_0.comparator_1.vnn.n13 70.9612
R30268 por_ana_0.comparator_1.vnn.n0 por_ana_0.comparator_1.vnn.n12 70.9612
R30269 por_ana_0.comparator_1.vnn.n0 por_ana_0.comparator_1.vnn.n11 70.9612
R30270 por_ana_0.comparator_1.vnn.n0 por_ana_0.comparator_1.vnn.n10 70.9612
R30271 por_ana_0.comparator_1.vnn.n0 por_ana_0.comparator_1.vnn.n9 70.9612
R30272 por_ana_0.comparator_1.vnn.n21 por_ana_0.comparator_1.vnn.t28 27.6955
R30273 por_ana_0.comparator_1.vnn.n21 por_ana_0.comparator_1.vnn.t23 27.6955
R30274 por_ana_0.comparator_1.vnn.n22 por_ana_0.comparator_1.vnn.t27 27.6955
R30275 por_ana_0.comparator_1.vnn.n22 por_ana_0.comparator_1.vnn.t22 27.6955
R30276 por_ana_0.comparator_1.vnn.n23 por_ana_0.comparator_1.vnn.t26 27.6955
R30277 por_ana_0.comparator_1.vnn.n23 por_ana_0.comparator_1.vnn.t21 27.6955
R30278 por_ana_0.comparator_1.vnn.n24 por_ana_0.comparator_1.vnn.t25 27.6955
R30279 por_ana_0.comparator_1.vnn.n24 por_ana_0.comparator_1.vnn.t20 27.6955
R30280 por_ana_0.comparator_1.vnn.n25 por_ana_0.comparator_1.vnn.t18 27.6955
R30281 por_ana_0.comparator_1.vnn.n25 por_ana_0.comparator_1.vnn.t17 27.6955
R30282 por_ana_0.comparator_1.vnn.n26 por_ana_0.comparator_1.vnn.t24 27.6955
R30283 por_ana_0.comparator_1.vnn.n26 por_ana_0.comparator_1.vnn.t19 27.6955
R30284 por_ana_0.comparator_1.vnn.n17 por_ana_0.comparator_1.vnn.t3 27.6955
R30285 por_ana_0.comparator_1.vnn.n17 por_ana_0.comparator_1.vnn.t15 27.6955
R30286 por_ana_0.comparator_1.vnn.n16 por_ana_0.comparator_1.vnn.t11 27.6955
R30287 por_ana_0.comparator_1.vnn.n16 por_ana_0.comparator_1.vnn.t7 27.6955
R30288 por_ana_0.comparator_1.vnn.n18 por_ana_0.comparator_1.vnn.t1 27.6955
R30289 por_ana_0.comparator_1.vnn.n18 por_ana_0.comparator_1.vnn.t13 27.6955
R30290 por_ana_0.comparator_1.vnn.n19 por_ana_0.comparator_1.vnn.t9 27.6955
R30291 por_ana_0.comparator_1.vnn.n19 por_ana_0.comparator_1.vnn.t5 27.6955
R30292 por_ana_0.comparator_1.vnn.n20 por_ana_0.comparator_1.vnn.t16 27.6955
R30293 por_ana_0.comparator_1.vnn.n20 por_ana_0.comparator_1.vnn.t29 27.6955
R30294 por_ana_0.comparator_1.vnn.n15 por_ana_0.comparator_1.vnn.t37 16.5305
R30295 por_ana_0.comparator_1.vnn.n15 por_ana_0.comparator_1.vnn.t41 16.5305
R30296 por_ana_0.comparator_1.vnn.n14 por_ana_0.comparator_1.vnn.t32 16.5305
R30297 por_ana_0.comparator_1.vnn.n14 por_ana_0.comparator_1.vnn.t44 16.5305
R30298 por_ana_0.comparator_1.vnn.n13 por_ana_0.comparator_1.vnn.t36 16.5305
R30299 por_ana_0.comparator_1.vnn.n13 por_ana_0.comparator_1.vnn.t40 16.5305
R30300 por_ana_0.comparator_1.vnn.n12 por_ana_0.comparator_1.vnn.t33 16.5305
R30301 por_ana_0.comparator_1.vnn.n12 por_ana_0.comparator_1.vnn.t45 16.5305
R30302 por_ana_0.comparator_1.vnn.n11 por_ana_0.comparator_1.vnn.t35 16.5305
R30303 por_ana_0.comparator_1.vnn.n11 por_ana_0.comparator_1.vnn.t39 16.5305
R30304 por_ana_0.comparator_1.vnn.n10 por_ana_0.comparator_1.vnn.t31 16.5305
R30305 por_ana_0.comparator_1.vnn.n10 por_ana_0.comparator_1.vnn.t43 16.5305
R30306 por_ana_0.comparator_1.vnn.n9 por_ana_0.comparator_1.vnn.t34 16.5305
R30307 por_ana_0.comparator_1.vnn.n9 por_ana_0.comparator_1.vnn.t38 16.5305
R30308 por_ana_0.comparator_1.vnn.n8 por_ana_0.comparator_1.vnn.t30 16.5305
R30309 por_ana_0.comparator_1.vnn.n8 por_ana_0.comparator_1.vnn.t42 16.5305
R30310 por_ana_0.comparator_1.vnn.n1 por_ana_0.comparator_1.vnn.t56 16.4779
R30311 por_ana_0.comparator_1.vnn.n3 por_ana_0.comparator_1.vnn.t47 16.4779
R30312 por_ana_0.comparator_1.vnn.n4 por_ana_0.comparator_1.vnn.t48 16.4779
R30313 por_ana_0.comparator_1.vnn.n2 por_ana_0.comparator_1.vnn.t49 16.4779
R30314 por_ana_0.comparator_1.vnn.n1 por_ana_0.comparator_1.vnn.t50 16.4779
R30315 por_ana_0.comparator_1.vnn.n1 por_ana_0.comparator_1.vnn.t53 16.4779
R30316 por_ana_0.comparator_1.vnn.n1 por_ana_0.comparator_1.vnn.t51 16.4779
R30317 por_ana_0.comparator_1.vnn.n5 por_ana_0.comparator_1.vnn.t57 16.4779
R30318 por_ana_0.comparator_1.vnn.n6 por_ana_0.comparator_1.vnn.t4 14.2251
R30319 por_ana_0.comparator_1.vnn.n6 por_ana_0.comparator_1.vnn.t8 14.2251
R30320 por_ana_0.comparator_1.vnn.n6 por_ana_0.comparator_1.vnn.t12 14.2251
R30321 por_ana_0.comparator_1.vnn.n6 por_ana_0.comparator_1.vnn.t0 14.2251
R30322 por_ana_0.comparator_1.vnn.n6 por_ana_0.comparator_1.vnn.t6 14.2251
R30323 por_ana_0.comparator_1.vnn.n6 por_ana_0.comparator_1.vnn.t10 14.2251
R30324 por_ana_0.comparator_1.vnn.n6 por_ana_0.comparator_1.vnn.t2 14.2251
R30325 por_ana_0.comparator_1.vnn.n6 por_ana_0.comparator_1.vnn.t14 14.2251
R30326 por_ana_0.comparator_1.vnn por_ana_0.comparator_1.vnn.n1 13.4051
R30327 por_ana_0.comparator_1.vnn por_ana_0.comparator_1.vnn.n0 11.9816
R30328 por_ana_0.comparator_1.vnn.n1 por_ana_0.comparator_1.vnn.t54 11.9724
R30329 por_ana_0.comparator_1.vnn.n3 por_ana_0.comparator_1.vnn.t58 11.9724
R30330 por_ana_0.comparator_1.vnn.n4 por_ana_0.comparator_1.vnn.t59 11.9724
R30331 por_ana_0.comparator_1.vnn.n2 por_ana_0.comparator_1.vnn.t60 11.9724
R30332 por_ana_0.comparator_1.vnn.n1 por_ana_0.comparator_1.vnn.t61 11.9724
R30333 por_ana_0.comparator_1.vnn.n1 por_ana_0.comparator_1.vnn.t52 11.9724
R30334 por_ana_0.comparator_1.vnn.n1 por_ana_0.comparator_1.vnn.t62 11.9724
R30335 por_ana_0.comparator_1.vnn.n5 por_ana_0.comparator_1.vnn.t55 11.9724
R30336 por_ana_0.comparator_1.vnn por_ana_0.comparator_1.vnn.n7 9.57847
R30337 por_ana_0.comparator_1.vnn.n1 por_ana_0.comparator_1.vnn.n4 9.23963
R30338 por_ana_0.comparator_1.vnn.n1 por_ana_0.comparator_1.vnn.n3 9.23963
R30339 por_ana_0.comparator_1.vnn.n1 por_ana_0.comparator_1.vnn.n2 9.23963
R30340 por_ana_0.comparator_1.vnn.n1 por_ana_0.comparator_1.vnn.n5 9.22553
R30341 por_ana_0.comparator_1.vnn.n7 por_ana_0.comparator_1.vnn.n6 8.84171
R30342 por_ana_0.comparator_1.vt.n21 por_ana_0.comparator_1.vt.n20 22508.4
R30343 por_ana_0.comparator_1.vt.n24 por_ana_0.comparator_1.vt.n21 22508.4
R30344 por_ana_0.comparator_1.vt.n24 por_ana_0.comparator_1.vt.n22 22508.4
R30345 por_ana_0.comparator_1.vt.n22 por_ana_0.comparator_1.vt.n20 22508.4
R30346 por_ana_0.comparator_1.vt.n18 por_ana_0.comparator_1.vt.n16 2577.69
R30347 por_ana_0.comparator_1.vt.n18 por_ana_0.comparator_1.vt.n14 2577.69
R30348 por_ana_0.comparator_1.vt.n17 por_ana_0.comparator_1.vt.n16 2577.69
R30349 por_ana_0.comparator_1.vt.n14 por_ana_0.comparator_1.vt.n17 2577.69
R30350 por_ana_0.comparator_1.vt.t36 por_ana_0.comparator_1.vt.t3 1757.46
R30351 por_ana_0.comparator_1.vt.t20 por_ana_0.comparator_1.vt.t36 1757.46
R30352 por_ana_0.comparator_1.vt.t18 por_ana_0.comparator_1.vt.t41 1757.46
R30353 por_ana_0.comparator_1.vt.t41 por_ana_0.comparator_1.vt.t0 1757.46
R30354 por_ana_0.comparator_1.vt.t3 por_ana_0.comparator_1.vt.n22 1032.7
R30355 por_ana_0.comparator_1.vt.t0 por_ana_0.comparator_1.vt.n21 1032.7
R30356 por_ana_0.comparator_1.vt.n23 por_ana_0.comparator_1.vt.t20 878.729
R30357 por_ana_0.comparator_1.vt.n23 por_ana_0.comparator_1.vt.t18 878.729
R30358 por_ana_0.comparator_1.vt.n13 por_ana_0.comparator_1.vt.t7 87.4912
R30359 por_ana_0.comparator_1.vt.n5 por_ana_0.comparator_1.vt.t16 87.4912
R30360 por_ana_0.comparator_1.vt.n5 por_ana_0.comparator_1.vt.t9 87.4912
R30361 por_ana_0.comparator_1.vt.n5 por_ana_0.comparator_1.vt.t15 87.4912
R30362 por_ana_0.comparator_1.vt.n5 por_ana_0.comparator_1.vt.t5 87.4912
R30363 por_ana_0.comparator_1.vt.n4 por_ana_0.comparator_1.vt.t13 87.4912
R30364 por_ana_0.comparator_1.vt.n4 por_ana_0.comparator_1.vt.t4 87.4912
R30365 por_ana_0.comparator_1.vt.n6 por_ana_0.comparator_1.vt.t14 87.4912
R30366 por_ana_0.comparator_1.vt.n6 por_ana_0.comparator_1.vt.t6 87.4912
R30367 por_ana_0.comparator_1.vt.n7 por_ana_0.comparator_1.vt.t12 87.4912
R30368 por_ana_0.comparator_1.vt.n7 por_ana_0.comparator_1.vt.t8 87.4912
R30369 por_ana_0.comparator_1.vt.n7 por_ana_0.comparator_1.vt.t11 87.4912
R30370 por_ana_0.comparator_1.vt.n7 por_ana_0.comparator_1.vt.t2 87.4912
R30371 por_ana_0.comparator_1.vt.n12 por_ana_0.comparator_1.vt.t10 87.4912
R30372 por_ana_0.comparator_1.vt.n12 por_ana_0.comparator_1.vt.t1 87.4912
R30373 por_ana_0.comparator_1.vt.t17 por_ana_0.comparator_1.vt.n13 87.4912
R30374 por_ana_0.comparator_1.vt.n2 por_ana_0.comparator_1.vt.n19 73.2112
R30375 por_ana_0.comparator_1.vt.n9 por_ana_0.comparator_1.vt.n32 70.9612
R30376 por_ana_0.comparator_1.vt.n9 por_ana_0.comparator_1.vt.n31 70.9612
R30377 por_ana_0.comparator_1.vt.n1 por_ana_0.comparator_1.vt.n30 70.9612
R30378 por_ana_0.comparator_1.vt.n1 por_ana_0.comparator_1.vt.n29 70.9612
R30379 por_ana_0.comparator_1.vt.n1 por_ana_0.comparator_1.vt.n28 70.9612
R30380 por_ana_0.comparator_1.vt.n1 por_ana_0.comparator_1.vt.n27 70.9612
R30381 por_ana_0.comparator_1.vt.n0 por_ana_0.comparator_1.vt.n26 70.9612
R30382 por_ana_0.comparator_1.vt.n0 por_ana_0.comparator_1.vt.n25 70.9612
R30383 por_ana_0.comparator_1.vt.n2 por_ana_0.comparator_1.vt.n36 70.9612
R30384 por_ana_0.comparator_1.vt.n2 por_ana_0.comparator_1.vt.n37 70.9612
R30385 por_ana_0.comparator_1.vt.n3 por_ana_0.comparator_1.vt.n38 70.9612
R30386 por_ana_0.comparator_1.vt.n3 por_ana_0.comparator_1.vt.n39 70.9612
R30387 por_ana_0.comparator_1.vt.n3 por_ana_0.comparator_1.vt.n40 70.9612
R30388 por_ana_0.comparator_1.vt.n3 por_ana_0.comparator_1.vt.n41 70.9612
R30389 por_ana_0.comparator_1.vt.n8 por_ana_0.comparator_1.vt.n42 70.9612
R30390 por_ana_0.comparator_1.vt.n8 por_ana_0.comparator_1.vt.n43 70.9612
R30391 por_ana_0.comparator_1.vt.n32 por_ana_0.comparator_1.vt.t33 16.5305
R30392 por_ana_0.comparator_1.vt.n32 por_ana_0.comparator_1.vt.t49 16.5305
R30393 por_ana_0.comparator_1.vt.n31 por_ana_0.comparator_1.vt.t24 16.5305
R30394 por_ana_0.comparator_1.vt.n31 por_ana_0.comparator_1.vt.t42 16.5305
R30395 por_ana_0.comparator_1.vt.n30 por_ana_0.comparator_1.vt.t34 16.5305
R30396 por_ana_0.comparator_1.vt.n30 por_ana_0.comparator_1.vt.t50 16.5305
R30397 por_ana_0.comparator_1.vt.n29 por_ana_0.comparator_1.vt.t25 16.5305
R30398 por_ana_0.comparator_1.vt.n29 por_ana_0.comparator_1.vt.t43 16.5305
R30399 por_ana_0.comparator_1.vt.n28 por_ana_0.comparator_1.vt.t19 16.5305
R30400 por_ana_0.comparator_1.vt.n28 por_ana_0.comparator_1.vt.t53 16.5305
R30401 por_ana_0.comparator_1.vt.n27 por_ana_0.comparator_1.vt.t26 16.5305
R30402 por_ana_0.comparator_1.vt.n27 por_ana_0.comparator_1.vt.t44 16.5305
R30403 por_ana_0.comparator_1.vt.n26 por_ana_0.comparator_1.vt.t35 16.5305
R30404 por_ana_0.comparator_1.vt.n26 por_ana_0.comparator_1.vt.t51 16.5305
R30405 por_ana_0.comparator_1.vt.n25 por_ana_0.comparator_1.vt.t27 16.5305
R30406 por_ana_0.comparator_1.vt.n25 por_ana_0.comparator_1.vt.t45 16.5305
R30407 por_ana_0.comparator_1.vt.n19 por_ana_0.comparator_1.vt.t54 16.5305
R30408 por_ana_0.comparator_1.vt.n19 por_ana_0.comparator_1.vt.t55 16.5305
R30409 por_ana_0.comparator_1.vt.n36 por_ana_0.comparator_1.vt.t40 16.5305
R30410 por_ana_0.comparator_1.vt.n36 por_ana_0.comparator_1.vt.t32 16.5305
R30411 por_ana_0.comparator_1.vt.n37 por_ana_0.comparator_1.vt.t48 16.5305
R30412 por_ana_0.comparator_1.vt.n37 por_ana_0.comparator_1.vt.t23 16.5305
R30413 por_ana_0.comparator_1.vt.n38 por_ana_0.comparator_1.vt.t39 16.5305
R30414 por_ana_0.comparator_1.vt.n38 por_ana_0.comparator_1.vt.t31 16.5305
R30415 por_ana_0.comparator_1.vt.n39 por_ana_0.comparator_1.vt.t52 16.5305
R30416 por_ana_0.comparator_1.vt.n39 por_ana_0.comparator_1.vt.t28 16.5305
R30417 por_ana_0.comparator_1.vt.n40 por_ana_0.comparator_1.vt.t38 16.5305
R30418 por_ana_0.comparator_1.vt.n40 por_ana_0.comparator_1.vt.t30 16.5305
R30419 por_ana_0.comparator_1.vt.n41 por_ana_0.comparator_1.vt.t47 16.5305
R30420 por_ana_0.comparator_1.vt.n41 por_ana_0.comparator_1.vt.t22 16.5305
R30421 por_ana_0.comparator_1.vt.n42 por_ana_0.comparator_1.vt.t37 16.5305
R30422 por_ana_0.comparator_1.vt.n42 por_ana_0.comparator_1.vt.t29 16.5305
R30423 por_ana_0.comparator_1.vt.n43 por_ana_0.comparator_1.vt.t46 16.5305
R30424 por_ana_0.comparator_1.vt.n43 por_ana_0.comparator_1.vt.t21 16.5305
R30425 por_ana_0.comparator_1.vt.n22 por_ana_0.comparator_1.vt.n16 11.9393
R30426 por_ana_0.comparator_1.vt.n14 por_ana_0.comparator_1.vt.n21 11.9393
R30427 por_ana_0.comparator_1.vt.n0 por_ana_0.comparator_1.vt.n2 10.3229
R30428 por_ana_0.comparator_1.vt.n45 por_ana_0.comparator_1.vt.n44 7.14705
R30429 por_ana_0.comparator_1.vt.n34 por_ana_0.comparator_1.vt.n33 7.14705
R30430 por_ana_0.comparator_1.vt.n35 por_ana_0.comparator_1.vt.n15 7.14705
R30431 por_ana_0.comparator_1.vt.n11 por_ana_0.comparator_1.vt.n10 7.14705
R30432 por_ana_0.comparator_1.vt.n6 por_ana_0.comparator_1.vt.n11 5.19386
R30433 por_ana_0.comparator_1.vt.n13 por_ana_0.comparator_1.vt.n15 5.19386
R30434 por_ana_0.comparator_1.vt.n44 por_ana_0.comparator_1.vt.n8 5.04137
R30435 por_ana_0.comparator_1.vt.n33 por_ana_0.comparator_1.vt.n9 5.04137
R30436 por_ana_0.comparator_1.vt.n34 por_ana_0.comparator_1.vt.n12 4.95167
R30437 por_ana_0.comparator_1.vt.n4 por_ana_0.comparator_1.vt.n45 4.95167
R30438 por_ana_0.comparator_1.vt.n8 por_ana_0.comparator_1.vt.n3 4.88031
R30439 por_ana_0.comparator_1.vt.n0 por_ana_0.comparator_1.vt.n10 4.5005
R30440 por_ana_0.comparator_1.vt.n2 por_ana_0.comparator_1.vt.n35 4.5005
R30441 por_ana_0.comparator_1.vt.n16 por_ana_0.comparator_1.vt.n15 4.20915
R30442 por_ana_0.comparator_1.vt.n14 por_ana_0.comparator_1.vt.n11 4.20915
R30443 por_ana_0.comparator_1.vt.n14 por_ana_0.comparator_1.vt.n34 4.01128
R30444 por_ana_0.comparator_1.vt.n45 por_ana_0.comparator_1.vt.n16 4.01128
R30445 por_ana_0.comparator_1.vt.n18 por_ana_0.comparator_1.vt.n20 3.9532
R30446 por_ana_0.comparator_1.vt.n23 por_ana_0.comparator_1.vt.n20 3.9532
R30447 por_ana_0.comparator_1.vt.n17 por_ana_0.comparator_1.vt.n24 3.9532
R30448 por_ana_0.comparator_1.vt.n24 por_ana_0.comparator_1.vt.n23 3.9532
R30449 por_ana_0.comparator_1.vt.n9 por_ana_0.comparator_1.vt.n1 3.90435
R30450 por_ana_0.comparator_1.vt.n1 por_ana_0.comparator_1.vt.n0 3.76733
R30451 por_ana_0.comparator_1.vt.n3 por_ana_0.comparator_1.vt.n2 3.70723
R30452 por_ana_0.comparator_1.vt.n35 por_ana_0.comparator_1.vt.n18 3.6402
R30453 por_ana_0.comparator_1.vt.n44 por_ana_0.comparator_1.vt.n17 3.6402
R30454 por_ana_0.comparator_1.vt.n33 por_ana_0.comparator_1.vt.n17 3.57378
R30455 por_ana_0.comparator_1.vt.n18 por_ana_0.comparator_1.vt.n10 3.57378
R30456 por_ana_0.comparator_1.vt.n12 por_ana_0.comparator_1.vt.n7 3.26612
R30457 por_ana_0.comparator_1.vt.n5 por_ana_0.comparator_1.vt.n4 3.26612
R30458 por_ana_0.comparator_1.vt.n13 por_ana_0.comparator_1.vt.n5 2.44972
R30459 por_ana_0.comparator_1.vt.n7 por_ana_0.comparator_1.vt.n6 2.44972
R30460 por_ana_0.comparator_0.n1.n2 por_ana_0.comparator_0.n1.t8 227.657
R30461 por_ana_0.comparator_0.n1.n2 por_ana_0.comparator_0.n1.t19 227.173
R30462 por_ana_0.comparator_0.n1.n2 por_ana_0.comparator_0.n1.t14 227.173
R30463 por_ana_0.comparator_0.n1.n2 por_ana_0.comparator_0.n1.t13 227.173
R30464 por_ana_0.comparator_0.n1.n2 por_ana_0.comparator_0.n1.t4 227.173
R30465 por_ana_0.comparator_0.n1.n2 por_ana_0.comparator_0.n1.t15 227.173
R30466 por_ana_0.comparator_0.n1.n2 por_ana_0.comparator_0.n1.t9 227.173
R30467 por_ana_0.comparator_0.n1.n2 por_ana_0.comparator_0.n1.t5 227.173
R30468 por_ana_0.comparator_0.n1.n0 por_ana_0.comparator_0.n1.t16 224.042
R30469 por_ana_0.comparator_0.n1.n0 por_ana_0.comparator_0.n1.t10 223.559
R30470 por_ana_0.comparator_0.n1.n0 por_ana_0.comparator_0.n1.t6 223.559
R30471 por_ana_0.comparator_0.n1.n0 por_ana_0.comparator_0.n1.t17 223.559
R30472 por_ana_0.comparator_0.n1.n0 por_ana_0.comparator_0.n1.t12 223.559
R30473 por_ana_0.comparator_0.n1.n0 por_ana_0.comparator_0.n1.t7 223.559
R30474 por_ana_0.comparator_0.n1.n0 por_ana_0.comparator_0.n1.t18 223.559
R30475 por_ana_0.comparator_0.n1.n0 por_ana_0.comparator_0.n1.t11 223.559
R30476 por_ana_0.comparator_0.n1.n1 por_ana_0.comparator_0.n1.n3 204.31
R30477 por_ana_0.comparator_0.n1.n4 por_ana_0.comparator_0.n1.n1 71.6326
R30478 por_ana_0.comparator_0.n1.n3 por_ana_0.comparator_0.n1.t2 27.6955
R30479 por_ana_0.comparator_0.n1.n3 por_ana_0.comparator_0.n1.t0 27.6955
R30480 por_ana_0.comparator_0.n1.t1 por_ana_0.comparator_0.n1.n4 16.5305
R30481 por_ana_0.comparator_0.n1.n4 por_ana_0.comparator_0.n1.t3 16.5305
R30482 por_ana_0.comparator_0.n1.n1 por_ana_0.comparator_0.n1.n0 11.9908
R30483 por_ana_0.comparator_0.n1.n1 por_ana_0.comparator_0.n1.n2 8.13016
R30484 porb_h.n2 porb_h.n1 157.593
R30485 porb_h.n43 porb_h.n42 157.591
R30486 porb_h.n38 porb_h.n37 157.591
R30487 porb_h.n32 porb_h.n31 157.591
R30488 porb_h.n26 porb_h.n25 157.591
R30489 porb_h.n20 porb_h.n19 157.591
R30490 porb_h.n14 porb_h.n13 157.591
R30491 porb_h.n8 porb_h.n7 157.591
R30492 porb_h.n43 porb_h.n41 136.965
R30493 porb_h.n38 porb_h.n36 136.965
R30494 porb_h.n32 porb_h.n30 136.965
R30495 porb_h.n26 porb_h.n24 136.965
R30496 porb_h.n20 porb_h.n18 136.965
R30497 porb_h.n14 porb_h.n12 136.965
R30498 porb_h.n8 porb_h.n6 136.965
R30499 porb_h.n2 porb_h.n0 136.965
R30500 porb_h.n41 porb_h.t29 21.2805
R30501 porb_h.n41 porb_h.t30 21.2805
R30502 porb_h.n36 porb_h.t28 21.2805
R30503 porb_h.n36 porb_h.t27 21.2805
R30504 porb_h.n30 porb_h.t25 21.2805
R30505 porb_h.n30 porb_h.t24 21.2805
R30506 porb_h.n24 porb_h.t21 21.2805
R30507 porb_h.n24 porb_h.t20 21.2805
R30508 porb_h.n18 porb_h.t19 21.2805
R30509 porb_h.n18 porb_h.t16 21.2805
R30510 porb_h.n12 porb_h.t26 21.2805
R30511 porb_h.n12 porb_h.t23 21.2805
R30512 porb_h.n6 porb_h.t22 21.2805
R30513 porb_h.n6 porb_h.t31 21.2805
R30514 porb_h.n0 porb_h.t18 21.2805
R30515 porb_h.n0 porb_h.t17 21.2805
R30516 porb_h.n42 porb_h.t0 17.8272
R30517 porb_h.n42 porb_h.t2 17.8272
R30518 porb_h.n37 porb_h.t15 17.8272
R30519 porb_h.n37 porb_h.t1 17.8272
R30520 porb_h.n31 porb_h.t12 17.8272
R30521 porb_h.n31 porb_h.t11 17.8272
R30522 porb_h.n25 porb_h.t8 17.8272
R30523 porb_h.n25 porb_h.t7 17.8272
R30524 porb_h.n19 porb_h.t14 17.8272
R30525 porb_h.n19 porb_h.t3 17.8272
R30526 porb_h.n13 porb_h.t13 17.8272
R30527 porb_h.n13 porb_h.t10 17.8272
R30528 porb_h.n7 porb_h.t9 17.8272
R30529 porb_h.n7 porb_h.t6 17.8272
R30530 porb_h.n1 porb_h.t5 17.8272
R30531 porb_h.n1 porb_h.t4 17.8272
R30532 porb_h.n44 porb_h.n43 10.1618
R30533 porb_h.n3 porb_h.n2 9.98018
R30534 porb_h.n39 porb_h.n38 9.98018
R30535 porb_h.n33 porb_h.n32 9.98018
R30536 porb_h.n27 porb_h.n26 9.98018
R30537 porb_h.n21 porb_h.n20 9.98018
R30538 porb_h.n15 porb_h.n14 9.98018
R30539 porb_h.n9 porb_h.n8 9.98018
R30540 porb_h.n44 porb_h 8.39491
R30541 porb_h.n40 porb_h 7.09609
R30542 porb_h.n34 porb_h 5.94903
R30543 porb_h.n35 porb_h 5.08746
R30544 porb_h.n28 porb_h 4.80197
R30545 porb_h.n29 porb_h 4.23963
R30546 porb_h porb_h.n45 3.88917
R30547 porb_h.n22 porb_h 3.65491
R30548 porb_h.n23 porb_h 3.3918
R30549 porb_h.n17 porb_h 2.54398
R30550 porb_h.n16 porb_h 2.50785
R30551 porb_h.n11 porb_h 1.69615
R30552 porb_h.n10 porb_h 1.36079
R30553 porb_h.n5 porb_h.n4 0.934324
R30554 porb_h.n11 porb_h.n10 0.934324
R30555 porb_h.n17 porb_h.n16 0.934324
R30556 porb_h.n23 porb_h.n22 0.934324
R30557 porb_h.n29 porb_h.n28 0.934324
R30558 porb_h.n35 porb_h.n34 0.934324
R30559 porb_h.n5 porb_h 0.848326
R30560 porb_h.n45 porb_h.n44 0.252453
R30561 porb_h.n45 porb_h.n40 0.224765
R30562 porb_h.n4 porb_h 0.213735
R30563 porb_h.n4 porb_h.n3 0.0793043
R30564 porb_h.n3 porb_h 0.0793043
R30565 porb_h.n10 porb_h.n9 0.0793043
R30566 porb_h.n9 porb_h.n5 0.0793043
R30567 porb_h.n16 porb_h.n15 0.0793043
R30568 porb_h.n15 porb_h.n11 0.0793043
R30569 porb_h.n22 porb_h.n21 0.0793043
R30570 porb_h.n21 porb_h.n17 0.0793043
R30571 porb_h.n28 porb_h.n27 0.0793043
R30572 porb_h.n27 porb_h.n23 0.0793043
R30573 porb_h.n34 porb_h.n33 0.0793043
R30574 porb_h.n33 porb_h.n29 0.0793043
R30575 porb_h.n40 porb_h.n39 0.0793043
R30576 porb_h.n39 porb_h.n35 0.0793043
R30577 por_dig_0.otrip_decoded[5].n1 por_dig_0.otrip_decoded[5].n0 289.849
R30578 por_dig_0.otrip_decoded[5].n2 por_dig_0.otrip_decoded[5].t4 186.374
R30579 por_dig_0.otrip_decoded[5].n9 por_dig_0.otrip_decoded[5].n8 185
R30580 por_dig_0.otrip_decoded[5].n2 por_dig_0.otrip_decoded[5].t5 170.308
R30581 por_dig_0.otrip_decoded[5].n3 por_dig_0.otrip_decoded[5] 154.56
R30582 por_dig_0.otrip_decoded[5].n4 por_dig_0.otrip_decoded[5].n3 153.462
R30583 por_dig_0.otrip_decoded[5].n3 por_dig_0.otrip_decoded[5].n2 101.513
R30584 por_dig_0.otrip_decoded[5] por_dig_0.otrip_decoded[5].n9 81.3181
R30585 por_dig_0.otrip_decoded[5].n6 por_dig_0.otrip_decoded[5].n5 32.8055
R30586 por_dig_0.otrip_decoded[5].n0 por_dig_0.otrip_decoded[5].t3 26.5955
R30587 por_dig_0.otrip_decoded[5].n0 por_dig_0.otrip_decoded[5].t2 26.5955
R30588 por_dig_0.otrip_decoded[5].n8 por_dig_0.otrip_decoded[5].t1 24.9236
R30589 por_dig_0.otrip_decoded[5].n8 por_dig_0.otrip_decoded[5].t0 24.9236
R30590 por_dig_0.otrip_decoded[5].n7 por_dig_0.otrip_decoded[5] 18.234
R30591 por_dig_0.otrip_decoded[5] por_dig_0.otrip_decoded[5].n1 9.15439
R30592 por_dig_0.otrip_decoded[5].n1 por_dig_0.otrip_decoded[5] 7.71085
R30593 por_dig_0.otrip_decoded[5].n5 por_dig_0.otrip_decoded[5].n4 4.96991
R30594 por_dig_0.otrip_decoded[5].n7 por_dig_0.otrip_decoded[5] 4.26717
R30595 por_dig_0.otrip_decoded[5].n4 por_dig_0.otrip_decoded[5] 3.46403
R30596 por_dig_0.otrip_decoded[5].n5 por_dig_0.otrip_decoded[5] 2.71109
R30597 por_dig_0.otrip_decoded[5] por_dig_0.otrip_decoded[5].n6 2.51389
R30598 por_dig_0.otrip_decoded[5].n6 por_dig_0.otrip_decoded[5] 2.26389
R30599 por_dig_0.otrip_decoded[5].n9 por_dig_0.otrip_decoded[5].n7 1.00442
R30600 por_dig_0.otrip_decoded[3].n2 por_dig_0.otrip_decoded[3].n1 289.849
R30601 por_dig_0.otrip_decoded[3].n3 por_dig_0.otrip_decoded[3].t4 186.374
R30602 por_dig_0.otrip_decoded[3].n9 por_dig_0.otrip_decoded[3].n8 185
R30603 por_dig_0.otrip_decoded[3].n3 por_dig_0.otrip_decoded[3].t5 170.308
R30604 por_dig_0.otrip_decoded[3].n4 por_dig_0.otrip_decoded[3] 154.56
R30605 por_dig_0.otrip_decoded[3].n5 por_dig_0.otrip_decoded[3].n4 153.462
R30606 por_dig_0.otrip_decoded[3].n4 por_dig_0.otrip_decoded[3].n3 101.513
R30607 por_dig_0.otrip_decoded[3] por_dig_0.otrip_decoded[3].n9 81.3181
R30608 por_dig_0.otrip_decoded[3].n0 por_dig_0.otrip_decoded[3].n6 36.0141
R30609 por_dig_0.otrip_decoded[3].n1 por_dig_0.otrip_decoded[3].t3 26.5955
R30610 por_dig_0.otrip_decoded[3].n1 por_dig_0.otrip_decoded[3].t2 26.5955
R30611 por_dig_0.otrip_decoded[3].n8 por_dig_0.otrip_decoded[3].t0 24.9236
R30612 por_dig_0.otrip_decoded[3].n8 por_dig_0.otrip_decoded[3].t1 24.9236
R30613 por_dig_0.otrip_decoded[3].n7 por_dig_0.otrip_decoded[3] 18.234
R30614 por_dig_0.otrip_decoded[3] por_dig_0.otrip_decoded[3].n2 9.15439
R30615 por_dig_0.otrip_decoded[3].n2 por_dig_0.otrip_decoded[3] 7.71085
R30616 por_dig_0.otrip_decoded[3].n6 por_dig_0.otrip_decoded[3].n5 4.96991
R30617 por_dig_0.otrip_decoded[3].n7 por_dig_0.otrip_decoded[3] 4.26717
R30618 por_dig_0.otrip_decoded[3] por_dig_0.otrip_decoded[3].n0 3.50496
R30619 por_dig_0.otrip_decoded[3].n5 por_dig_0.otrip_decoded[3] 3.46403
R30620 por_dig_0.otrip_decoded[3].n6 por_dig_0.otrip_decoded[3] 2.71109
R30621 por_dig_0.otrip_decoded[3].n0 por_dig_0.otrip_decoded[3] 1.49604
R30622 por_dig_0.otrip_decoded[3].n0 por_dig_0.otrip_decoded[3] 1.39633
R30623 por_dig_0.otrip_decoded[3].n0 por_dig_0.otrip_decoded[3] 1.32193
R30624 por_dig_0.otrip_decoded[3].n9 por_dig_0.otrip_decoded[3].n7 1.00442
R30625 por_ana_0.comparator_0.vt.n23 por_ana_0.comparator_0.vt.n21 22508.4
R30626 por_ana_0.comparator_0.vt.n23 por_ana_0.comparator_0.vt.n20 22508.4
R30627 por_ana_0.comparator_0.vt.n20 por_ana_0.comparator_0.vt.n19 22508.4
R30628 por_ana_0.comparator_0.vt.n21 por_ana_0.comparator_0.vt.n19 22508.4
R30629 por_ana_0.comparator_0.vt.n12 por_ana_0.comparator_0.vt.n13 2577.69
R30630 por_ana_0.comparator_0.vt.n14 por_ana_0.comparator_0.vt.n13 2577.69
R30631 por_ana_0.comparator_0.vt.n15 por_ana_0.comparator_0.vt.n14 2577.69
R30632 por_ana_0.comparator_0.vt.n12 por_ana_0.comparator_0.vt.n15 2577.69
R30633 por_ana_0.comparator_0.vt.t3 por_ana_0.comparator_0.vt.t21 1757.46
R30634 por_ana_0.comparator_0.vt.t36 por_ana_0.comparator_0.vt.t3 1757.46
R30635 por_ana_0.comparator_0.vt.t0 por_ana_0.comparator_0.vt.t40 1757.46
R30636 por_ana_0.comparator_0.vt.t18 por_ana_0.comparator_0.vt.t0 1757.46
R30637 por_ana_0.comparator_0.vt.t21 por_ana_0.comparator_0.vt.n19 1032.7
R30638 por_ana_0.comparator_0.vt.n23 por_ana_0.comparator_0.vt.t18 1032.7
R30639 por_ana_0.comparator_0.vt.n22 por_ana_0.comparator_0.vt.t36 878.729
R30640 por_ana_0.comparator_0.vt.t40 por_ana_0.comparator_0.vt.n22 878.729
R30641 por_ana_0.comparator_0.vt.n10 por_ana_0.comparator_0.vt.t29 87.4912
R30642 por_ana_0.comparator_0.vt.n10 por_ana_0.comparator_0.vt.t35 87.4912
R30643 por_ana_0.comparator_0.vt.n7 por_ana_0.comparator_0.vt.t23 87.4912
R30644 por_ana_0.comparator_0.vt.n7 por_ana_0.comparator_0.vt.t28 87.4912
R30645 por_ana_0.comparator_0.vt.n7 por_ana_0.comparator_0.vt.t34 87.4912
R30646 por_ana_0.comparator_0.vt.n7 por_ana_0.comparator_0.vt.t27 87.4912
R30647 por_ana_0.comparator_0.vt.n6 por_ana_0.comparator_0.vt.t33 87.4912
R30648 por_ana_0.comparator_0.vt.n6 por_ana_0.comparator_0.vt.t22 87.4912
R30649 por_ana_0.comparator_0.vt.n4 por_ana_0.comparator_0.vt.t26 87.4912
R30650 por_ana_0.comparator_0.vt.n4 por_ana_0.comparator_0.vt.t32 87.4912
R30651 por_ana_0.comparator_0.vt.n5 por_ana_0.comparator_0.vt.t20 87.4912
R30652 por_ana_0.comparator_0.vt.n5 por_ana_0.comparator_0.vt.t25 87.4912
R30653 por_ana_0.comparator_0.vt.n5 por_ana_0.comparator_0.vt.t31 87.4912
R30654 por_ana_0.comparator_0.vt.n5 por_ana_0.comparator_0.vt.t24 87.4912
R30655 por_ana_0.comparator_0.vt.n11 por_ana_0.comparator_0.vt.t30 87.4912
R30656 por_ana_0.comparator_0.vt.n11 por_ana_0.comparator_0.vt.t19 87.4912
R30657 por_ana_0.comparator_0.vt.n1 por_ana_0.comparator_0.vt.n17 73.2112
R30658 por_ana_0.comparator_0.vt.n9 por_ana_0.comparator_0.vt.n44 70.9612
R30659 por_ana_0.comparator_0.vt.n9 por_ana_0.comparator_0.vt.n43 70.9612
R30660 por_ana_0.comparator_0.vt.n0 por_ana_0.comparator_0.vt.n42 70.9612
R30661 por_ana_0.comparator_0.vt.n0 por_ana_0.comparator_0.vt.n41 70.9612
R30662 por_ana_0.comparator_0.vt.n0 por_ana_0.comparator_0.vt.n40 70.9612
R30663 por_ana_0.comparator_0.vt.n1 por_ana_0.comparator_0.vt.n18 70.9612
R30664 por_ana_0.comparator_0.vt.n1 por_ana_0.comparator_0.vt.n24 70.9612
R30665 por_ana_0.comparator_0.vt.n2 por_ana_0.comparator_0.vt.n25 70.9612
R30666 por_ana_0.comparator_0.vt.n2 por_ana_0.comparator_0.vt.n26 70.9612
R30667 por_ana_0.comparator_0.vt.n2 por_ana_0.comparator_0.vt.n27 70.9612
R30668 por_ana_0.comparator_0.vt.n2 por_ana_0.comparator_0.vt.n28 70.9612
R30669 por_ana_0.comparator_0.vt.n8 por_ana_0.comparator_0.vt.n29 70.9612
R30670 por_ana_0.comparator_0.vt.n8 por_ana_0.comparator_0.vt.n30 70.9612
R30671 por_ana_0.comparator_0.vt.n3 por_ana_0.comparator_0.vt.n35 70.9612
R30672 por_ana_0.comparator_0.vt.n3 por_ana_0.comparator_0.vt.n16 70.9612
R30673 por_ana_0.comparator_0.vt.n45 por_ana_0.comparator_0.vt.n9 70.9612
R30674 por_ana_0.comparator_0.vt.n44 por_ana_0.comparator_0.vt.t52 16.5305
R30675 por_ana_0.comparator_0.vt.n44 por_ana_0.comparator_0.vt.t2 16.5305
R30676 por_ana_0.comparator_0.vt.n43 por_ana_0.comparator_0.vt.t42 16.5305
R30677 por_ana_0.comparator_0.vt.n43 por_ana_0.comparator_0.vt.t11 16.5305
R30678 por_ana_0.comparator_0.vt.n42 por_ana_0.comparator_0.vt.t51 16.5305
R30679 por_ana_0.comparator_0.vt.n42 por_ana_0.comparator_0.vt.t1 16.5305
R30680 por_ana_0.comparator_0.vt.n41 por_ana_0.comparator_0.vt.t41 16.5305
R30681 por_ana_0.comparator_0.vt.n41 por_ana_0.comparator_0.vt.t10 16.5305
R30682 por_ana_0.comparator_0.vt.n40 por_ana_0.comparator_0.vt.t46 16.5305
R30683 por_ana_0.comparator_0.vt.n40 por_ana_0.comparator_0.vt.t16 16.5305
R30684 por_ana_0.comparator_0.vt.n17 por_ana_0.comparator_0.vt.t54 16.5305
R30685 por_ana_0.comparator_0.vt.n17 por_ana_0.comparator_0.vt.t55 16.5305
R30686 por_ana_0.comparator_0.vt.n18 por_ana_0.comparator_0.vt.t15 16.5305
R30687 por_ana_0.comparator_0.vt.n18 por_ana_0.comparator_0.vt.t50 16.5305
R30688 por_ana_0.comparator_0.vt.n24 por_ana_0.comparator_0.vt.t7 16.5305
R30689 por_ana_0.comparator_0.vt.n24 por_ana_0.comparator_0.vt.t39 16.5305
R30690 por_ana_0.comparator_0.vt.n25 por_ana_0.comparator_0.vt.t9 16.5305
R30691 por_ana_0.comparator_0.vt.n25 por_ana_0.comparator_0.vt.t45 16.5305
R30692 por_ana_0.comparator_0.vt.n26 por_ana_0.comparator_0.vt.t14 16.5305
R30693 por_ana_0.comparator_0.vt.n26 por_ana_0.comparator_0.vt.t49 16.5305
R30694 por_ana_0.comparator_0.vt.n27 por_ana_0.comparator_0.vt.t5 16.5305
R30695 por_ana_0.comparator_0.vt.n27 por_ana_0.comparator_0.vt.t38 16.5305
R30696 por_ana_0.comparator_0.vt.n28 por_ana_0.comparator_0.vt.t13 16.5305
R30697 por_ana_0.comparator_0.vt.n28 por_ana_0.comparator_0.vt.t48 16.5305
R30698 por_ana_0.comparator_0.vt.n29 por_ana_0.comparator_0.vt.t4 16.5305
R30699 por_ana_0.comparator_0.vt.n29 por_ana_0.comparator_0.vt.t37 16.5305
R30700 por_ana_0.comparator_0.vt.n30 por_ana_0.comparator_0.vt.t8 16.5305
R30701 por_ana_0.comparator_0.vt.n30 por_ana_0.comparator_0.vt.t44 16.5305
R30702 por_ana_0.comparator_0.vt.n35 por_ana_0.comparator_0.vt.t53 16.5305
R30703 por_ana_0.comparator_0.vt.n35 por_ana_0.comparator_0.vt.t6 16.5305
R30704 por_ana_0.comparator_0.vt.n16 por_ana_0.comparator_0.vt.t43 16.5305
R30705 por_ana_0.comparator_0.vt.n16 por_ana_0.comparator_0.vt.t12 16.5305
R30706 por_ana_0.comparator_0.vt.n45 por_ana_0.comparator_0.vt.t47 16.5305
R30707 por_ana_0.comparator_0.vt.t17 por_ana_0.comparator_0.vt.n45 16.5305
R30708 por_ana_0.comparator_0.vt.n14 por_ana_0.comparator_0.vt.n23 11.9393
R30709 por_ana_0.comparator_0.vt.n12 por_ana_0.comparator_0.vt.n19 11.9393
R30710 por_ana_0.comparator_0.vt.n3 por_ana_0.comparator_0.vt.n1 10.3229
R30711 por_ana_0.comparator_0.vt.n34 por_ana_0.comparator_0.vt.n33 7.14705
R30712 por_ana_0.comparator_0.vt.n37 por_ana_0.comparator_0.vt.n36 7.14705
R30713 por_ana_0.comparator_0.vt.n32 por_ana_0.comparator_0.vt.n31 7.14705
R30714 por_ana_0.comparator_0.vt.n39 por_ana_0.comparator_0.vt.n38 7.14705
R30715 por_ana_0.comparator_0.vt.n33 por_ana_0.comparator_0.vt.n10 5.19386
R30716 por_ana_0.comparator_0.vt.n4 por_ana_0.comparator_0.vt.n37 5.19386
R30717 por_ana_0.comparator_0.vt.n31 por_ana_0.comparator_0.vt.n8 5.04137
R30718 por_ana_0.comparator_0.vt.n0 por_ana_0.comparator_0.vt.n39 5.04137
R30719 por_ana_0.comparator_0.vt.n6 por_ana_0.comparator_0.vt.n32 4.95167
R30720 por_ana_0.comparator_0.vt.n38 por_ana_0.comparator_0.vt.n11 4.95167
R30721 por_ana_0.comparator_0.vt.n8 por_ana_0.comparator_0.vt.n2 4.88031
R30722 por_ana_0.comparator_0.vt.n36 por_ana_0.comparator_0.vt.n3 4.5005
R30723 por_ana_0.comparator_0.vt.n1 por_ana_0.comparator_0.vt.n34 4.5005
R30724 por_ana_0.comparator_0.vt.n37 por_ana_0.comparator_0.vt.n14 4.20915
R30725 por_ana_0.comparator_0.vt.n33 por_ana_0.comparator_0.vt.n12 4.20915
R30726 por_ana_0.comparator_0.vt.n32 por_ana_0.comparator_0.vt.n12 4.01128
R30727 por_ana_0.comparator_0.vt.n38 por_ana_0.comparator_0.vt.n14 4.01128
R30728 por_ana_0.comparator_0.vt.n21 por_ana_0.comparator_0.vt.n13 3.9532
R30729 por_ana_0.comparator_0.vt.n22 por_ana_0.comparator_0.vt.n21 3.9532
R30730 por_ana_0.comparator_0.vt.n15 por_ana_0.comparator_0.vt.n20 3.9532
R30731 por_ana_0.comparator_0.vt.n22 por_ana_0.comparator_0.vt.n20 3.9532
R30732 por_ana_0.comparator_0.vt.n9 por_ana_0.comparator_0.vt.n0 3.90435
R30733 por_ana_0.comparator_0.vt.n9 por_ana_0.comparator_0.vt.n3 3.76733
R30734 por_ana_0.comparator_0.vt.n2 por_ana_0.comparator_0.vt.n1 3.70723
R30735 por_ana_0.comparator_0.vt.n31 por_ana_0.comparator_0.vt.n15 3.6402
R30736 por_ana_0.comparator_0.vt.n34 por_ana_0.comparator_0.vt.n13 3.6402
R30737 por_ana_0.comparator_0.vt.n36 por_ana_0.comparator_0.vt.n13 3.57378
R30738 por_ana_0.comparator_0.vt.n39 por_ana_0.comparator_0.vt.n15 3.57378
R30739 por_ana_0.comparator_0.vt.n7 por_ana_0.comparator_0.vt.n6 3.26612
R30740 por_ana_0.comparator_0.vt.n11 por_ana_0.comparator_0.vt.n5 3.26612
R30741 por_ana_0.comparator_0.vt.n5 por_ana_0.comparator_0.vt.n4 2.44972
R30742 por_ana_0.comparator_0.vt.n10 por_ana_0.comparator_0.vt.n7 2.44972
R30743 por_dig_0.otrip_decoded[6].n1 por_dig_0.otrip_decoded[6].n0 289.849
R30744 por_dig_0.otrip_decoded[6].n2 por_dig_0.otrip_decoded[6].t4 186.374
R30745 por_dig_0.otrip_decoded[6].n9 por_dig_0.otrip_decoded[6].n8 185
R30746 por_dig_0.otrip_decoded[6].n2 por_dig_0.otrip_decoded[6].t5 170.308
R30747 por_dig_0.otrip_decoded[6].n3 por_dig_0.otrip_decoded[6] 154.56
R30748 por_dig_0.otrip_decoded[6].n4 por_dig_0.otrip_decoded[6].n3 153.462
R30749 por_dig_0.otrip_decoded[6].n3 por_dig_0.otrip_decoded[6].n2 101.513
R30750 por_dig_0.otrip_decoded[6] por_dig_0.otrip_decoded[6].n9 81.3181
R30751 por_dig_0.otrip_decoded[6].n6 por_dig_0.otrip_decoded[6].n5 34.7028
R30752 por_dig_0.otrip_decoded[6].n0 por_dig_0.otrip_decoded[6].t3 26.5955
R30753 por_dig_0.otrip_decoded[6].n0 por_dig_0.otrip_decoded[6].t2 26.5955
R30754 por_dig_0.otrip_decoded[6].n8 por_dig_0.otrip_decoded[6].t0 24.9236
R30755 por_dig_0.otrip_decoded[6].n8 por_dig_0.otrip_decoded[6].t1 24.9236
R30756 por_dig_0.otrip_decoded[6].n7 por_dig_0.otrip_decoded[6] 15.243
R30757 por_dig_0.otrip_decoded[6] por_dig_0.otrip_decoded[6].n6 10.9291
R30758 por_dig_0.otrip_decoded[6] por_dig_0.otrip_decoded[6].n1 9.15439
R30759 por_dig_0.otrip_decoded[6].n1 por_dig_0.otrip_decoded[6] 7.71085
R30760 por_dig_0.otrip_decoded[6].n5 por_dig_0.otrip_decoded[6].n4 4.96991
R30761 por_dig_0.otrip_decoded[6].n7 por_dig_0.otrip_decoded[6] 4.26717
R30762 por_dig_0.otrip_decoded[6].n4 por_dig_0.otrip_decoded[6] 3.46403
R30763 por_dig_0.otrip_decoded[6].n6 por_dig_0.otrip_decoded[6] 2.89336
R30764 por_dig_0.otrip_decoded[6].n5 por_dig_0.otrip_decoded[6] 2.71109
R30765 por_dig_0.otrip_decoded[6].n9 por_dig_0.otrip_decoded[6].n7 1.00442
R30766 por_ana_0.ibias_gen_0.vn1.n0 por_ana_0.ibias_gen_0.vn1.n1 47.4959
R30767 por_ana_0.ibias_gen_0.vn1.n3 por_ana_0.ibias_gen_0.vn1.t12 27.5855
R30768 por_ana_0.ibias_gen_0.vn1.n2 por_ana_0.ibias_gen_0.vn1.t11 27.5855
R30769 por_ana_0.ibias_gen_0.vn1.n6 por_ana_0.ibias_gen_0.vn1.t17 27.5855
R30770 por_ana_0.ibias_gen_0.vn1.n5 por_ana_0.ibias_gen_0.vn1.t15 27.5855
R30771 por_ana_0.ibias_gen_0.vn1.n10 por_ana_0.ibias_gen_0.vn1.t4 26.004
R30772 por_ana_0.ibias_gen_0.vn1.n0 por_ana_0.ibias_gen_0.vn1.n13 24.5059
R30773 por_ana_0.ibias_gen_0.vn1.n3 por_ana_0.ibias_gen_0.vn1.t10 24.3247
R30774 por_ana_0.ibias_gen_0.vn1.n2 por_ana_0.ibias_gen_0.vn1.t16 24.3247
R30775 por_ana_0.ibias_gen_0.vn1.n6 por_ana_0.ibias_gen_0.vn1.t14 24.3247
R30776 por_ana_0.ibias_gen_0.vn1.n5 por_ana_0.ibias_gen_0.vn1.t13 24.3247
R30777 por_ana_0.ibias_gen_0.vn1.n9 por_ana_0.ibias_gen_0.vn1.t2 24.3247
R30778 por_ana_0.ibias_gen_0.vn1.n14 por_ana_0.ibias_gen_0.vn1.n0 17.1535
R30779 por_ana_0.ibias_gen_0.vn1.n12 por_ana_0.ibias_gen_0.vn1.n11 13.8791
R30780 por_ana_0.ibias_gen_0.vn1.n0 por_ana_0.ibias_gen_0.vn1.n12 12.7397
R30781 por_ana_0.ibias_gen_0.vn1.n1 por_ana_0.ibias_gen_0.vn1.t7 5.5395
R30782 por_ana_0.ibias_gen_0.vn1.n1 por_ana_0.ibias_gen_0.vn1.t0 5.5395
R30783 por_ana_0.ibias_gen_0.vn1.n4 por_ana_0.ibias_gen_0.vn1.n2 4.66645
R30784 por_ana_0.ibias_gen_0.vn1.n7 por_ana_0.ibias_gen_0.vn1.n5 4.66645
R30785 por_ana_0.ibias_gen_0.vn1.n13 por_ana_0.ibias_gen_0.vn1.t6 3.3065
R30786 por_ana_0.ibias_gen_0.vn1.n13 por_ana_0.ibias_gen_0.vn1.t8 3.3065
R30787 por_ana_0.ibias_gen_0.vn1.n11 por_ana_0.ibias_gen_0.vn1.t3 3.3065
R30788 por_ana_0.ibias_gen_0.vn1.n11 por_ana_0.ibias_gen_0.vn1.t5 3.3065
R30789 por_ana_0.ibias_gen_0.vn1.n14 por_ana_0.ibias_gen_0.vn1.t9 3.3065
R30790 por_ana_0.ibias_gen_0.vn1.t1 por_ana_0.ibias_gen_0.vn1.n14 3.3065
R30791 por_ana_0.ibias_gen_0.vn1.n8 por_ana_0.ibias_gen_0.vn1.n4 2.41645
R30792 por_ana_0.ibias_gen_0.vn1.n8 por_ana_0.ibias_gen_0.vn1.n7 2.41645
R30793 por_ana_0.ibias_gen_0.vn1.n4 por_ana_0.ibias_gen_0.vn1.n3 2.2505
R30794 por_ana_0.ibias_gen_0.vn1.n7 por_ana_0.ibias_gen_0.vn1.n6 2.2505
R30795 por_ana_0.ibias_gen_0.vn1.n9 por_ana_0.ibias_gen_0.vn1.n8 2.2505
R30796 por_ana_0.ibias_gen_0.vn1.n10 por_ana_0.ibias_gen_0.vn1.n9 1.58202
R30797 por_ana_0.ibias_gen_0.vn1.n12 por_ana_0.ibias_gen_0.vn1.n10 1.37822
R30798 por_ana_0.ibias_gen_0.vp1.n5 por_ana_0.ibias_gen_0.vp1.n4 53.0003
R30799 por_ana_0.ibias_gen_0.vp1.t10 por_ana_0.ibias_gen_0.vp1.n3 49.8109
R30800 por_ana_0.ibias_gen_0.vp1.n3 por_ana_0.ibias_gen_0.vp1.t12 49.8109
R30801 por_ana_0.ibias_gen_0.vp1.t12 por_ana_0.ibias_gen_0.vp1.n0 49.7878
R30802 por_ana_0.ibias_gen_0.vp1.n0 por_ana_0.ibias_gen_0.vp1.t10 49.6053
R30803 por_ana_0.ibias_gen_0.vp1 por_ana_0.ibias_gen_0.vp1.n6 45.7548
R30804 por_ana_0.ibias_gen_0.vp1.n2 por_ana_0.ibias_gen_0.vp1.n1 42.4505
R30805 por_ana_0.ibias_gen_0.vp1.n9 por_ana_0.ibias_gen_0.vp1.n7 18.5825
R30806 por_ana_0.ibias_gen_0.vp1.n15 por_ana_0.ibias_gen_0.vp1.n14 17.1535
R30807 por_ana_0.ibias_gen_0.vp1.n11 por_ana_0.ibias_gen_0.vp1.n10 16.3247
R30808 por_ana_0.ibias_gen_0.vp1.n9 por_ana_0.ibias_gen_0.vp1.n8 16.3247
R30809 por_ana_0.ibias_gen_0.vp1.n13 por_ana_0.ibias_gen_0.vp1.n12 15.5548
R30810 por_ana_0.ibias_gen_0.vp1.n15 por_ana_0.ibias_gen_0.vp1.n13 11.684
R30811 por_ana_0.ibias_gen_0.vp1.n6 por_ana_0.ibias_gen_0.vp1.t0 5.5395
R30812 por_ana_0.ibias_gen_0.vp1.n6 por_ana_0.ibias_gen_0.vp1.t14 5.5395
R30813 por_ana_0.ibias_gen_0.vp1.n4 por_ana_0.ibias_gen_0.vp1.t17 5.5395
R30814 por_ana_0.ibias_gen_0.vp1.n4 por_ana_0.ibias_gen_0.vp1.t16 5.5395
R30815 por_ana_0.ibias_gen_0.vp1.n1 por_ana_0.ibias_gen_0.vp1.t13 5.5395
R30816 por_ana_0.ibias_gen_0.vp1.n1 por_ana_0.ibias_gen_0.vp1.t11 5.5395
R30817 por_ana_0.ibias_gen_0.vp1.n5 por_ana_0.ibias_gen_0.vp1.n0 4.85318
R30818 por_ana_0.ibias_gen_0.vp1.n11 por_ana_0.ibias_gen_0.vp1.n9 4.51612
R30819 por_ana_0.ibias_gen_0.vp1.n12 por_ana_0.ibias_gen_0.vp1.t3 3.3065
R30820 por_ana_0.ibias_gen_0.vp1.n12 por_ana_0.ibias_gen_0.vp1.t8 3.3065
R30821 por_ana_0.ibias_gen_0.vp1.n10 por_ana_0.ibias_gen_0.vp1.t9 3.3065
R30822 por_ana_0.ibias_gen_0.vp1.n10 por_ana_0.ibias_gen_0.vp1.t7 3.3065
R30823 por_ana_0.ibias_gen_0.vp1.n8 por_ana_0.ibias_gen_0.vp1.t5 3.3065
R30824 por_ana_0.ibias_gen_0.vp1.n8 por_ana_0.ibias_gen_0.vp1.t2 3.3065
R30825 por_ana_0.ibias_gen_0.vp1.n7 por_ana_0.ibias_gen_0.vp1.t6 3.3065
R30826 por_ana_0.ibias_gen_0.vp1.n7 por_ana_0.ibias_gen_0.vp1.t4 3.3065
R30827 por_ana_0.ibias_gen_0.vp1.n14 por_ana_0.ibias_gen_0.vp1.t1 3.3065
R30828 por_ana_0.ibias_gen_0.vp1.n14 por_ana_0.ibias_gen_0.vp1.t15 3.3065
R30829 por_ana_0.ibias_gen_0.vp1.n13 por_ana_0.ibias_gen_0.vp1.n11 2.27562
R30830 por_ana_0.ibias_gen_0.vp1 por_ana_0.ibias_gen_0.vp1.n15 1.87819
R30831 por_ana_0.ibias_gen_0.vp1.n2 por_ana_0.ibias_gen_0.vp1.n0 1.48628
R30832 por_ana_0.ibias_gen_0.vp1.n3 por_ana_0.ibias_gen_0.vp1.n2 1.47061
R30833 por_ana_0.ibias_gen_0.vp1 por_ana_0.ibias_gen_0.vp1.n5 1.36236
R30834 por_ana_0.rstring_mux_0.vtrip0.n5 por_ana_0.rstring_mux_0.vtrip0.n3 50.7022
R30835 por_ana_0.rstring_mux_0.vtrip0.n2 por_ana_0.rstring_mux_0.vtrip0.n0 50.7022
R30836 por_ana_0.rstring_mux_0.vtrip0.n7 por_ana_0.rstring_mux_0.vtrip0.n6 25.1771
R30837 por_ana_0.rstring_mux_0.vtrip0.n5 por_ana_0.rstring_mux_0.vtrip0.n4 13.8791
R30838 por_ana_0.rstring_mux_0.vtrip0.n2 por_ana_0.rstring_mux_0.vtrip0.n1 13.8791
R30839 por_ana_0.rstring_mux_0.vtrip0.n6 por_ana_0.rstring_mux_0.vtrip0.n5 13.7519
R30840 por_ana_0.rstring_mux_0.vtrip0.n7 por_ana_0.rstring_mux_0.vtrip0.t7 10.6303
R30841 por_ana_0.rstring_mux_0.vtrip0.n3 por_ana_0.rstring_mux_0.vtrip0.t4 5.5395
R30842 por_ana_0.rstring_mux_0.vtrip0.n3 por_ana_0.rstring_mux_0.vtrip0.t3 5.5395
R30843 por_ana_0.rstring_mux_0.vtrip0.n0 por_ana_0.rstring_mux_0.vtrip0.t6 5.5395
R30844 por_ana_0.rstring_mux_0.vtrip0.n0 por_ana_0.rstring_mux_0.vtrip0.t5 5.5395
R30845 por_ana_0.rstring_mux_0.vtrip0.n6 por_ana_0.rstring_mux_0.vtrip0.n2 3.60196
R30846 por_ana_0.rstring_mux_0.vtrip0.n4 por_ana_0.rstring_mux_0.vtrip0.t2 3.3065
R30847 por_ana_0.rstring_mux_0.vtrip0.n4 por_ana_0.rstring_mux_0.vtrip0.t1 3.3065
R30848 por_ana_0.rstring_mux_0.vtrip0.n1 por_ana_0.rstring_mux_0.vtrip0.t9 3.3065
R30849 por_ana_0.rstring_mux_0.vtrip0.n1 por_ana_0.rstring_mux_0.vtrip0.t8 3.3065
R30850 por_ana_0.rstring_mux_0.vtrip0 por_ana_0.rstring_mux_0.vtrip0.t0 0.769662
R30851 por_ana_0.rstring_mux_0.vtrip0 por_ana_0.rstring_mux_0.vtrip0.n7 0.0563195
R30852 por_dig_0.net20.n13 por_dig_0.net20 586.646
R30853 por_dig_0.net20.n14 por_dig_0.net20.n13 585
R30854 por_dig_0.net20.n13 por_dig_0.net20.n12 585
R30855 por_dig_0.net20.n6 por_dig_0.net20.t8 276.464
R30856 por_dig_0.net20.n2 por_dig_0.net20.t4 230.155
R30857 por_dig_0.net20.n0 por_dig_0.net20.t9 229.369
R30858 por_dig_0.net20.n9 por_dig_0.net20.t6 224.984
R30859 por_dig_0.net20 por_dig_0.net20.t0 209.923
R30860 por_dig_0.net20.n6 por_dig_0.net20.t5 196.131
R30861 por_dig_0.net20.n9 por_dig_0.net20.t2 187.714
R30862 por_dig_0.net20.n2 por_dig_0.net20.t7 157.856
R30863 por_dig_0.net20.n0 por_dig_0.net20.t3 157.07
R30864 por_dig_0.net20 por_dig_0.net20.n9 153.957
R30865 por_dig_0.net20.n7 por_dig_0.net20.n6 152
R30866 por_dig_0.net20.n3 por_dig_0.net20.n2 152
R30867 por_dig_0.net20.n1 por_dig_0.net20.n0 152
R30868 por_dig_0.net20.n5 por_dig_0.net20.n4 34.824
R30869 por_dig_0.net20.n13 por_dig_0.net20.t1 26.5955
R30870 por_dig_0.net20.n11 por_dig_0.net20.n8 24.6806
R30871 por_dig_0.net20 por_dig_0.net20.n11 19.317
R30872 por_dig_0.net20.n4 por_dig_0.net20 12.8005
R30873 por_dig_0.net20.n5 por_dig_0.net20.n1 12.6224
R30874 por_dig_0.net20.n14 por_dig_0.net20 10.7891
R30875 por_dig_0.net20 por_dig_0.net20.n12 10.7891
R30876 por_dig_0.net20.n8 por_dig_0.net20.n7 10.6843
R30877 por_dig_0.net20 por_dig_0.net20.n10 9.4552
R30878 por_dig_0.net20.n10 por_dig_0.net20 9.06717
R30879 por_dig_0.net20.n8 por_dig_0.net20.n5 8.28724
R30880 por_dig_0.net20.n11 por_dig_0.net20 4.63992
R30881 por_dig_0.net20.n10 por_dig_0.net20 3.02272
R30882 por_dig_0.net20.n3 por_dig_0.net20 2.76128
R30883 por_dig_0.net20.n1 por_dig_0.net20 2.10199
R30884 por_dig_0.net20 por_dig_0.net20.n14 1.64621
R30885 por_dig_0.net20.n12 por_dig_0.net20 1.64621
R30886 por_dig_0.net20.n7 por_dig_0.net20 1.55726
R30887 por_dig_0.net20.n4 por_dig_0.net20.n3 1.50638
R30888 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[7].n1 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[7].n0 873.303
R30889 por_ana_0.sky130_fd_sc_hvl__lsbuflv2hv_1_0[1|7].X por_ana_0.rstring_mux_0.vtrip_decoded_avdd[7].n1 585
R30890 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[7].t0 por_ana_0.sky130_fd_sc_hvl__lsbuflv2hv_1_0[1|7].X 511.971
R30891 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[7].n2 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[7].t2 384.704
R30892 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[7].n2 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[7].t3 384.226
R30893 por_ana_0.sky130_fd_sc_hvl__lsbuflv2hv_1_0[1|7].X por_ana_0.rstring_mux_0.vtrip_decoded_avdd[7].t1 155.607
R30894 por_ana_0.rstring_mux_0.sky130_fd_sc_hvl__inv_1_0[15].A por_ana_0.rstring_mux_0.vtrip_decoded_avdd[7].n3 153.165
R30895 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[7].n1 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[7].t0 147.756
R30896 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[7].n3 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[7].t5 114.031
R30897 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[7].n3 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[7].t4 81.5883
R30898 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[7].n6 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[7].n5 40.5975
R30899 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[7].n5 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[7].n4 13.8005
R30900 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[7].n5 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[7].n2 10.1657
R30901 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[7].n0 por_ana_0.sky130_fd_sc_hvl__lsbuflv2hv_1_0[1|7].X 8.85549
R30902 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[7].n4 por_ana_0.rstring_mux_0.sky130_fd_sc_hvl__inv_1_0[15].A 7.97972
R30903 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[7].n4 por_ana_0.rstring_mux_0.sky130_fd_sc_hvl__inv_1_0[15].A 7.97972
R30904 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[7].n6 por_ana_0.sky130_fd_sc_hvl__lsbuflv2hv_1_0[1|7].X 7.49318
R30905 por_ana_0.sky130_fd_sc_hvl__lsbuflv2hv_1_0[1|7].X por_ana_0.rstring_mux_0.vtrip_decoded_avdd[7].n0 4.05904
R30906 por_ana_0.sky130_fd_sc_hvl__lsbuflv2hv_1_0[1|7].X por_ana_0.rstring_mux_0.vtrip_decoded_avdd[7].n6 4.05904
R30907 por_ana_0.rstring_mux_0.vtrip7.n5 por_ana_0.rstring_mux_0.vtrip7.n3 50.7022
R30908 por_ana_0.rstring_mux_0.vtrip7.n2 por_ana_0.rstring_mux_0.vtrip7.n0 50.7022
R30909 por_ana_0.rstring_mux_0.vtrip7.n6 por_ana_0.rstring_mux_0.vtrip7.n5 15.3935
R30910 por_ana_0.rstring_mux_0.vtrip7.n5 por_ana_0.rstring_mux_0.vtrip7.n4 13.8791
R30911 por_ana_0.rstring_mux_0.vtrip7.n2 por_ana_0.rstring_mux_0.vtrip7.n1 13.8791
R30912 por_ana_0.rstring_mux_0.vtrip7.t6 por_ana_0.rstring_mux_0.vtrip7.n7 10.5857
R30913 por_ana_0.rstring_mux_0.vtrip7.n7 por_ana_0.rstring_mux_0.vtrip7.t7 10.5847
R30914 por_ana_0.rstring_mux_0.vtrip7.n3 por_ana_0.rstring_mux_0.vtrip7.t1 5.5395
R30915 por_ana_0.rstring_mux_0.vtrip7.n3 por_ana_0.rstring_mux_0.vtrip7.t0 5.5395
R30916 por_ana_0.rstring_mux_0.vtrip7.n0 por_ana_0.rstring_mux_0.vtrip7.t8 5.5395
R30917 por_ana_0.rstring_mux_0.vtrip7.n0 por_ana_0.rstring_mux_0.vtrip7.t9 5.5395
R30918 por_ana_0.rstring_mux_0.vtrip7.n6 por_ana_0.rstring_mux_0.vtrip7.n2 5.2741
R30919 por_ana_0.rstring_mux_0.vtrip7.n4 por_ana_0.rstring_mux_0.vtrip7.t5 3.3065
R30920 por_ana_0.rstring_mux_0.vtrip7.n4 por_ana_0.rstring_mux_0.vtrip7.t4 3.3065
R30921 por_ana_0.rstring_mux_0.vtrip7.n1 por_ana_0.rstring_mux_0.vtrip7.t2 3.3065
R30922 por_ana_0.rstring_mux_0.vtrip7.n1 por_ana_0.rstring_mux_0.vtrip7.t3 3.3065
R30923 por_ana_0.rstring_mux_0.vtrip7.n7 por_ana_0.rstring_mux_0.vtrip7.n6 2.48711
R30924 por_dig_0.otrip_decoded[7].n2 por_dig_0.otrip_decoded[7].n1 289.849
R30925 por_dig_0.otrip_decoded[7].n3 por_dig_0.otrip_decoded[7].t4 186.374
R30926 por_dig_0.otrip_decoded[7].n9 por_dig_0.otrip_decoded[7].n8 185
R30927 por_dig_0.otrip_decoded[7].n3 por_dig_0.otrip_decoded[7].t5 170.308
R30928 por_dig_0.otrip_decoded[7].n4 por_dig_0.otrip_decoded[7] 154.56
R30929 por_dig_0.otrip_decoded[7].n5 por_dig_0.otrip_decoded[7].n4 153.462
R30930 por_dig_0.otrip_decoded[7].n4 por_dig_0.otrip_decoded[7].n3 101.513
R30931 por_dig_0.otrip_decoded[7] por_dig_0.otrip_decoded[7].n9 81.3181
R30932 por_dig_0.otrip_decoded[7].n0 por_dig_0.otrip_decoded[7].n6 31.3316
R30933 por_dig_0.otrip_decoded[7].n1 por_dig_0.otrip_decoded[7].t3 26.5955
R30934 por_dig_0.otrip_decoded[7].n1 por_dig_0.otrip_decoded[7].t2 26.5955
R30935 por_dig_0.otrip_decoded[7].n8 por_dig_0.otrip_decoded[7].t1 24.9236
R30936 por_dig_0.otrip_decoded[7].n8 por_dig_0.otrip_decoded[7].t0 24.9236
R30937 por_dig_0.otrip_decoded[7].n7 por_dig_0.otrip_decoded[7] 18.234
R30938 por_dig_0.otrip_decoded[7] por_dig_0.otrip_decoded[7].n2 9.15439
R30939 por_dig_0.otrip_decoded[7].n2 por_dig_0.otrip_decoded[7] 7.71085
R30940 por_dig_0.otrip_decoded[7].n6 por_dig_0.otrip_decoded[7].n5 4.96991
R30941 por_dig_0.otrip_decoded[7].n7 por_dig_0.otrip_decoded[7] 4.26717
R30942 por_dig_0.otrip_decoded[7].n5 por_dig_0.otrip_decoded[7] 3.46403
R30943 por_dig_0.otrip_decoded[7] por_dig_0.otrip_decoded[7].n0 3.25586
R30944 por_dig_0.otrip_decoded[7].n6 por_dig_0.otrip_decoded[7] 2.71109
R30945 por_dig_0.otrip_decoded[7].n0 por_dig_0.otrip_decoded[7] 1.6322
R30946 por_dig_0.otrip_decoded[7].n0 por_dig_0.otrip_decoded[7] 1.60467
R30947 por_dig_0.otrip_decoded[7].n9 por_dig_0.otrip_decoded[7].n7 1.00442
R30948 otrip[1].n0 otrip[1].t2 323.55
R30949 otrip[1].n0 otrip[1].t3 195.017
R30950 otrip[1] otrip[1].n0 155.036
R30951 otrip[1].n3 otrip[1].n2 74.5413
R30952 otrip[1].n4 otrip[1].n1 20.2722
R30953 otrip[1].n2 otrip[1].t0 16.5305
R30954 otrip[1].n2 otrip[1].t1 16.5305
R30955 otrip[1].n4 otrip[1].n3 10.0822
R30956 otrip[1].n1 otrip[1] 6.7304
R30957 otrip[1].n1 otrip[1] 2.2438
R30958 otrip[1] otrip[1].n4 1.35764
R30959 otrip[1].n3 otrip[1] 0.690617
R30960 por_ana_0.comparator_0.vn.n1 por_ana_0.comparator_0.vn.t6 234.096
R30961 por_ana_0.comparator_0.vn.n2 por_ana_0.comparator_0.vn.t5 94.5098
R30962 por_ana_0.comparator_0.vn.n1 por_ana_0.comparator_0.vn.t0 87.5075
R30963 por_ana_0.comparator_0.vn.n0 por_ana_0.comparator_0.vn.n3 66.4612
R30964 por_ana_0.comparator_0.vn.n3 por_ana_0.comparator_0.vn.t2 16.5305
R30965 por_ana_0.comparator_0.vn.n3 por_ana_0.comparator_0.vn.t4 16.5305
R30966 por_ana_0.comparator_0.vn.n0 por_ana_0.comparator_0.vn.t7 16.2067
R30967 por_ana_0.comparator_0.vn.n0 por_ana_0.comparator_0.vn.t3 13.954
R30968 por_ana_0.comparator_0.vn.n0 por_ana_0.comparator_0.vn.t1 11.7013
R30969 por_ana_0.comparator_0.vn.n0 por_ana_0.comparator_0.vn.t8 11.7013
R30970 por_ana_0.comparator_0.vn por_ana_0.comparator_0.vn.n0 11.4244
R30971 por_ana_0.comparator_0.vn por_ana_0.comparator_0.vn.n2 10.7596
R30972 por_ana_0.comparator_0.vn.n2 por_ana_0.comparator_0.vn.n1 8.74658
R30973 por_dig_0.osc_ena.n5 por_dig_0.osc_ena.n4 585
R30974 por_dig_0.osc_ena.n6 por_dig_0.osc_ena.n5 585
R30975 por_dig_0.osc_ena.n1 por_dig_0.osc_ena.t5 413.582
R30976 por_dig_0.osc_ena.n0 por_dig_0.osc_ena.t6 348.789
R30977 por_dig_0.osc_ena.n1 por_dig_0.osc_ena.t4 227.718
R30978 por_dig_0.osc_ena.n0 por_dig_0.osc_ena.t7 224.327
R30979 por_dig_0.osc_ena.n3 por_dig_0.osc_ena.n2 185
R30980 por_dig_0.osc_ena.n4 por_dig_0.osc_ena 79.5613
R30981 por_dig_0.osc_ena.n5 por_dig_0.osc_ena.t3 26.5955
R30982 por_dig_0.osc_ena.n5 por_dig_0.osc_ena.t2 26.5955
R30983 por_dig_0.osc_ena.n2 por_dig_0.osc_ena.t1 24.9236
R30984 por_dig_0.osc_ena.n2 por_dig_0.osc_ena.t0 24.9236
R30985 por_dig_0.osc_ena.n3 por_dig_0.osc_ena 16.0287
R30986 por_dig_0.osc_ena por_dig_0.osc_ena.n0 13.8267
R30987 por_dig_0.osc_ena por_dig_0.osc_ena.n6 13.3025
R30988 por_dig_0.osc_ena por_dig_0.osc_ena.n4 7.02795
R30989 por_dig_0.osc_ena por_dig_0.osc_ena.n1 4.5005
R30990 por_dig_0.osc_ena.n6 por_dig_0.osc_ena 3.76521
R30991 por_dig_0.osc_ena por_dig_0.osc_ena.n3 3.26325
R30992 por_dig_0.otrip_decoded[2].n1 por_dig_0.otrip_decoded[2].n0 289.849
R30993 por_dig_0.otrip_decoded[2].n2 por_dig_0.otrip_decoded[2].t4 186.374
R30994 por_dig_0.otrip_decoded[2].n8 por_dig_0.otrip_decoded[2].n7 185
R30995 por_dig_0.otrip_decoded[2].n2 por_dig_0.otrip_decoded[2].t5 170.308
R30996 por_dig_0.otrip_decoded[2].n3 por_dig_0.otrip_decoded[2] 154.56
R30997 por_dig_0.otrip_decoded[2].n4 por_dig_0.otrip_decoded[2].n3 153.462
R30998 por_dig_0.otrip_decoded[2].n3 por_dig_0.otrip_decoded[2].n2 101.513
R30999 por_dig_0.otrip_decoded[2] por_dig_0.otrip_decoded[2].n8 81.3181
R31000 por_dig_0.otrip_decoded[2] por_dig_0.otrip_decoded[2].n5 36.832
R31001 por_dig_0.otrip_decoded[2].n0 por_dig_0.otrip_decoded[2].t3 26.5955
R31002 por_dig_0.otrip_decoded[2].n0 por_dig_0.otrip_decoded[2].t2 26.5955
R31003 por_dig_0.otrip_decoded[2].n7 por_dig_0.otrip_decoded[2].t1 24.9236
R31004 por_dig_0.otrip_decoded[2].n7 por_dig_0.otrip_decoded[2].t0 24.9236
R31005 por_dig_0.otrip_decoded[2].n6 por_dig_0.otrip_decoded[2] 20.2247
R31006 por_dig_0.otrip_decoded[2] por_dig_0.otrip_decoded[2].n1 9.15439
R31007 por_dig_0.otrip_decoded[2].n1 por_dig_0.otrip_decoded[2] 7.71085
R31008 por_dig_0.otrip_decoded[2].n5 por_dig_0.otrip_decoded[2].n4 4.96991
R31009 por_dig_0.otrip_decoded[2].n6 por_dig_0.otrip_decoded[2] 4.26717
R31010 por_dig_0.otrip_decoded[2].n4 por_dig_0.otrip_decoded[2] 3.46403
R31011 por_dig_0.otrip_decoded[2].n5 por_dig_0.otrip_decoded[2] 2.71109
R31012 por_dig_0.otrip_decoded[2].n8 por_dig_0.otrip_decoded[2].n6 1.00442
R31013 por_ana_0.rstring_mux_0.ena.n5 por_ana_0.rstring_mux_0.ena.n4 873.303
R31014 por_ana_0.sky130_fd_sc_hvl__lsbuflv2hv_1_0[0|8].X por_ana_0.rstring_mux_0.ena.n5 585
R31015 por_ana_0.rstring_mux_0.ena.t0 por_ana_0.sky130_fd_sc_hvl__lsbuflv2hv_1_0[0|8].X 511.971
R31016 por_ana_0.rstring_mux_0.ena.n1 por_ana_0.rstring_mux_0.ena.t4 392.176
R31017 por_ana_0.rstring_mux_0.ena.n0 por_ana_0.rstring_mux_0.ena.t3 220.19
R31018 por_ana_0.rstring_mux_0.ena.n0 por_ana_0.rstring_mux_0.ena.t13 216.667
R31019 por_ana_0.rstring_mux_0.ena.n9 por_ana_0.rstring_mux_0.ena.n8 152
R31020 por_ana_0.rstring_mux_0.ena.n5 por_ana_0.rstring_mux_0.ena.t0 147.756
R31021 por_ana_0.rstring_mux_0.ena.n2 por_ana_0.rstring_mux_0.ena.t5 125.388
R31022 por_ana_0.rstring_mux_0.ena.n2 por_ana_0.rstring_mux_0.ena.t6 124.674
R31023 por_ana_0.rstring_mux_0.ena.n2 por_ana_0.rstring_mux_0.ena.t7 124.674
R31024 por_ana_0.rstring_mux_0.ena.n3 por_ana_0.rstring_mux_0.ena.t10 123.192
R31025 por_ana_0.rstring_mux_0.ena.n3 por_ana_0.rstring_mux_0.ena.t2 122.623
R31026 por_ana_0.rstring_mux_0.ena.n8 por_ana_0.rstring_mux_0.ena.t12 114.031
R31027 por_ana_0.rstring_mux_0.ena.n0 por_ana_0.rstring_mux_0.ena.t8 100.222
R31028 por_ana_0.rstring_mux_0.ena.n8 por_ana_0.rstring_mux_0.ena.t9 81.5883
R31029 por_ana_0.rstring_mux_0.ena.n6 por_ana_0.rstring_mux_0.ena.t1 50.7343
R31030 por_ana_0.rstring_mux_0.ena.n6 por_ana_0.rstring_mux_0.ena.t11 50.112
R31031 por_ana_0.rstring_mux_0.ena.n11 por_ana_0.rstring_mux_0.ena.n10 42.0365
R31032 por_ana_0.rstring_mux_0.ena.n1 por_ana_0.rstring_mux_0.ena.n3 40.3455
R31033 por_ana_0.rstring_mux_0.ena.n1 por_ana_0.rstring_mux_0.ena.n6 31.9476
R31034 por_ana_0.rstring_mux_0.ena.n10 por_ana_0.rstring_mux_0.sky130_fd_sc_hvl__inv_1_1.A 21.1071
R31035 por_ana_0.rstring_mux_0.ena.n10 por_ana_0.rstring_mux_0.ena.n7 18.7092
R31036 por_ana_0.rstring_mux_0.sky130_fd_sc_hvl__inv_1_1.A por_ana_0.rstring_mux_0.ena.n9 11.4706
R31037 por_ana_0.rstring_mux_0.ena.n4 por_ana_0.sky130_fd_sc_hvl__lsbuflv2hv_1_0[0|8].X 8.85549
R31038 por_ana_0.rstring_mux_0.ena.n11 por_ana_0.sky130_fd_sc_hvl__lsbuflv2hv_1_0[0|8].X 7.49318
R31039 por_ana_0.rstring_mux_0.ena.n7 por_ana_0.rstring_mux_0.ena.n1 5.3151
R31040 por_ana_0.rstring_mux_0.ena.n7 por_ana_0.rstring_mux_0.ena.n0 4.82955
R31041 por_ana_0.rstring_mux_0.ena.n3 por_ana_0.rstring_mux_0.ena.n2 4.67042
R31042 por_ana_0.rstring_mux_0.ena.n9 por_ana_0.rstring_mux_0.sky130_fd_sc_hvl__inv_1_1.A 4.48881
R31043 por_ana_0.sky130_fd_sc_hvl__lsbuflv2hv_1_0[0|8].X por_ana_0.rstring_mux_0.ena.n4 4.05904
R31044 por_ana_0.sky130_fd_sc_hvl__lsbuflv2hv_1_0[0|8].X por_ana_0.rstring_mux_0.ena.n11 4.05904
R31045 por_ana_0.rc_osc_0.n.n4 por_ana_0.rc_osc_0.n.t10 244.843
R31046 por_ana_0.rc_osc_0.n.n2 por_ana_0.rc_osc_0.n.t11 240.778
R31047 por_ana_0.rc_osc_0.n.n3 por_ana_0.rc_osc_0.n.t8 240.349
R31048 por_ana_0.rc_osc_0.n.n2 por_ana_0.rc_osc_0.n.t9 240.349
R31049 por_ana_0.rc_osc_0.n.n10 por_ana_0.rc_osc_0.n.n0 211.296
R31050 por_ana_0.rc_osc_0.n.n11 por_ana_0.rc_osc_0.n.n10 204.284
R31051 por_ana_0.rc_osc_0.n.n7 por_ana_0.rc_osc_0.n.t6 123.462
R31052 por_ana_0.rc_osc_0.n.n5 por_ana_0.rc_osc_0.n.t12 120.871
R31053 por_ana_0.rc_osc_0.n.n6 por_ana_0.rc_osc_0.n.t7 120.773
R31054 por_ana_0.rc_osc_0.n.n5 por_ana_0.rc_osc_0.n.t13 120.174
R31055 por_ana_0.rc_osc_0.n.n9 por_ana_0.rc_osc_0.n.n1 72.3553
R31056 por_ana_0.rc_osc_0.n.n0 por_ana_0.rc_osc_0.n.t2 28.5655
R31057 por_ana_0.rc_osc_0.n.n0 por_ana_0.rc_osc_0.n.t1 28.5655
R31058 por_ana_0.rc_osc_0.n.n11 por_ana_0.rc_osc_0.n.t3 28.5655
R31059 por_ana_0.rc_osc_0.n.t5 por_ana_0.rc_osc_0.n.n11 28.5655
R31060 por_ana_0.rc_osc_0.n.n1 por_ana_0.rc_osc_0.n.t4 17.4005
R31061 por_ana_0.rc_osc_0.n.n1 por_ana_0.rc_osc_0.n.t0 17.4005
R31062 por_ana_0.rc_osc_0.n.n4 por_ana_0.rc_osc_0.n.n3 9.0153
R31063 por_ana_0.rc_osc_0.n.n7 por_ana_0.rc_osc_0.n.n6 5.23012
R31064 por_ana_0.rc_osc_0.n.n8 por_ana_0.rc_osc_0.n.n7 3.78258
R31065 por_ana_0.rc_osc_0.n.n9 por_ana_0.rc_osc_0.n.n8 3.4105
R31066 por_ana_0.rc_osc_0.n.n10 por_ana_0.rc_osc_0.n.n9 1.35184
R31067 por_ana_0.rc_osc_0.n.n3 por_ana_0.rc_osc_0.n.n2 0.408448
R31068 por_ana_0.rc_osc_0.n.n8 por_ana_0.rc_osc_0.n.n4 0.147461
R31069 por_ana_0.rc_osc_0.n.n6 por_ana_0.rc_osc_0.n.n5 0.049413
R31070 por_ana_0.comparator_0.vm por_ana_0.comparator_0.vm.n1 205.605
R31071 por_ana_0.comparator_0.vm por_ana_0.comparator_0.vm.t6 97.3098
R31072 por_ana_0.comparator_0.vm por_ana_0.comparator_0.vm.n2 66.4612
R31073 por_ana_0.comparator_0.vm.n1 por_ana_0.comparator_0.vm.t5 27.6955
R31074 por_ana_0.comparator_0.vm.n1 por_ana_0.comparator_0.vm.t4 27.6955
R31075 por_ana_0.comparator_0.vm.n2 por_ana_0.comparator_0.vm.t1 16.5305
R31076 por_ana_0.comparator_0.vm.n2 por_ana_0.comparator_0.vm.t3 16.5305
R31077 por_ana_0.comparator_0.vm.n0 por_ana_0.comparator_0.vm.t7 16.2067
R31078 por_ana_0.comparator_0.vm por_ana_0.comparator_0.vm.t2 13.954
R31079 por_ana_0.comparator_0.vm por_ana_0.comparator_0.vm.n0 12.146
R31080 por_ana_0.comparator_0.vm por_ana_0.comparator_0.vm.t0 11.7013
R31081 por_ana_0.comparator_0.vm.n0 por_ana_0.comparator_0.vm.t8 11.7013
R31082 por_ana_0.comparator_1.vm por_ana_0.comparator_1.vm.n1 205.605
R31083 por_ana_0.comparator_1.vm por_ana_0.comparator_1.vm.t6 97.3098
R31084 por_ana_0.comparator_1.vm por_ana_0.comparator_1.vm.n2 66.4612
R31085 por_ana_0.comparator_1.vm.n1 por_ana_0.comparator_1.vm.t1 27.6955
R31086 por_ana_0.comparator_1.vm.n1 por_ana_0.comparator_1.vm.t0 27.6955
R31087 por_ana_0.comparator_1.vm.n2 por_ana_0.comparator_1.vm.t5 16.5305
R31088 por_ana_0.comparator_1.vm.n2 por_ana_0.comparator_1.vm.t3 16.5305
R31089 por_ana_0.comparator_1.vm.n0 por_ana_0.comparator_1.vm.t7 16.2067
R31090 por_ana_0.comparator_1.vm por_ana_0.comparator_1.vm.t2 13.954
R31091 por_ana_0.comparator_1.vm por_ana_0.comparator_1.vm.n0 12.146
R31092 por_ana_0.comparator_1.vm por_ana_0.comparator_1.vm.t4 11.7013
R31093 por_ana_0.comparator_1.vm.n0 por_ana_0.comparator_1.vm.t8 11.7013
R31094 por_ana_0.comparator_0.ena_b.n0 por_ana_0.comparator_0.ena_b.t0 232.647
R31095 por_ana_0.comparator_0.ena_b.n0 por_ana_0.comparator_0.ena_b.t5 125.588
R31096 por_ana_0.comparator_0.ena_b.n0 por_ana_0.comparator_0.ena_b.t4 123.201
R31097 por_ana_0.comparator_0.ena_b.n0 por_ana_0.comparator_0.ena_b.t2 122.505
R31098 por_ana_0.comparator_0.ena_b.n0 por_ana_0.comparator_0.ena_b.t3 122.505
R31099 por_ana_0.comparator_0.ena_b.n0 por_ana_0.comparator_0.ena_b.t1 91.9743
R31100 por_ana_0.ibias_gen_0.isrc_sel.n2 por_ana_0.ibias_gen_0.isrc_sel.n1 873.303
R31101 por_ana_0.sky130_fd_sc_hvl__lsbuflv2hv_1_0[1|8].X por_ana_0.ibias_gen_0.isrc_sel.n2 585
R31102 por_ana_0.ibias_gen_0.isrc_sel.t0 por_ana_0.sky130_fd_sc_hvl__lsbuflv2hv_1_0[1|8].X 511.971
R31103 por_ana_0.ibias_gen_0.isrc_sel.n3 por_ana_0.ibias_gen_0.isrc_sel.t8 395.779
R31104 por_ana_0.ibias_gen_0.isrc_sel.n4 por_ana_0.ibias_gen_0.isrc_sel.t7 392.36
R31105 por_ana_0.ibias_gen_0.isrc_sel.n3 por_ana_0.ibias_gen_0.isrc_sel.t5 388.736
R31106 por_ana_0.ibias_gen_0.isrc_sel.n6 por_ana_0.ibias_gen_0.isrc_sel.t2 218.921
R31107 por_ana_0.ibias_gen_0.isrc_sel.n6 por_ana_0.ibias_gen_0.isrc_sel.t4 217.906
R31108 por_ana_0.ibias_gen_0.isrc_sel.n5 por_ana_0.ibias_gen_0.isrc_sel.t3 195.367
R31109 por_ana_0.sky130_fd_sc_hvl__lsbuflv2hv_1_0[1|8].X por_ana_0.ibias_gen_0.isrc_sel.t1 155.607
R31110 por_ana_0.ibias_gen_0.isrc_sel.n2 por_ana_0.ibias_gen_0.isrc_sel.t0 147.756
R31111 por_ana_0.ibias_gen_0.isrc_sel.n0 por_ana_0.ibias_gen_0.isrc_sel.t6 109.147
R31112 por_ana_0.ibias_gen_0.isrc_sel.n0 por_ana_0.ibias_gen_0.isrc_sel.t9 106.493
R31113 por_ana_0.ibias_gen_0.isrc_sel.n7 por_ana_0.ibias_gen_0.isrc_sel.n0 39.7612
R31114 por_ana_0.ibias_gen_0.isrc_sel.n1 por_ana_0.sky130_fd_sc_hvl__lsbuflv2hv_1_0[1|8].X 8.85549
R31115 por_ana_0.ibias_gen_0.isrc_sel.n0 por_ana_0.ibias_gen_0.isrc_sel.n6 8.73795
R31116 por_ana_0.ibias_gen_0.isrc_sel.n5 por_ana_0.ibias_gen_0.isrc_sel.n4 8.68564
R31117 por_ana_0.ibias_gen_0.isrc_sel.n4 por_ana_0.ibias_gen_0.isrc_sel.n3 8.5512
R31118 por_ana_0.ibias_gen_0.isrc_sel.n7 por_ana_0.sky130_fd_sc_hvl__lsbuflv2hv_1_0[1|8].X 7.49318
R31119 por_ana_0.ibias_gen_0.isrc_sel.n0 por_ana_0.ibias_gen_0.isrc_sel.n5 6.72285
R31120 por_ana_0.sky130_fd_sc_hvl__lsbuflv2hv_1_0[1|8].X por_ana_0.ibias_gen_0.isrc_sel.n1 4.05904
R31121 por_ana_0.sky130_fd_sc_hvl__lsbuflv2hv_1_0[1|8].X por_ana_0.ibias_gen_0.isrc_sel.n7 4.05904
R31122 por_ana_0.ibias_gen_0.isrc_sel_b.n3 por_ana_0.ibias_gen_0.isrc_sel_b.t4 399.517
R31123 por_ana_0.ibias_gen_0.isrc_sel_b.n0 por_ana_0.ibias_gen_0.isrc_sel_b.t7 392.901
R31124 por_ana_0.ibias_gen_0.isrc_sel_b.n3 por_ana_0.ibias_gen_0.isrc_sel_b.t6 392.341
R31125 por_ana_0.ibias_gen_0.isrc_sel_b.n1 por_ana_0.ibias_gen_0.isrc_sel_b.t8 106.712
R31126 por_ana_0.ibias_gen_0.isrc_sel_b.n1 por_ana_0.ibias_gen_0.isrc_sel_b.t5 105.582
R31127 por_ana_0.ibias_gen_0.isrc_sel_b.n4 por_ana_0.ibias_gen_0.isrc_sel_b.n2 46.6401
R31128 por_ana_0.ibias_gen_0.isrc_sel_b.n5 por_ana_0.ibias_gen_0.isrc_sel_b.n4 18.0932
R31129 por_ana_0.ibias_gen_0.isrc_sel_b.n2 por_ana_0.ibias_gen_0.isrc_sel_b.t2 5.5395
R31130 por_ana_0.ibias_gen_0.isrc_sel_b.n2 por_ana_0.ibias_gen_0.isrc_sel_b.t0 5.5395
R31131 por_ana_0.ibias_gen_0.isrc_sel_b.n4 por_ana_0.ibias_gen_0.isrc_sel_b.n1 4.62075
R31132 por_ana_0.ibias_gen_0.isrc_sel_b.n0 por_ana_0.ibias_gen_0.isrc_sel_b.n3 4.00633
R31133 por_ana_0.ibias_gen_0.isrc_sel_b.n5 por_ana_0.ibias_gen_0.isrc_sel_b.t3 3.3065
R31134 por_ana_0.ibias_gen_0.isrc_sel_b.t1 por_ana_0.ibias_gen_0.isrc_sel_b.n5 3.3065
R31135 por_ana_0.ibias_gen_0.isrc_sel_b.n1 por_ana_0.ibias_gen_0.isrc_sel_b.n0 1.8288
R31136 por_dig_0._036_.n6 por_dig_0._036_.t8 241.439
R31137 por_dig_0._036_.n1 por_dig_0._036_.t6 240.484
R31138 por_dig_0._036_.n3 por_dig_0._036_.t7 233.01
R31139 por_dig_0._036_.n9 por_dig_0._036_.t1 218.572
R31140 por_dig_0._036_.n6 por_dig_0._036_.t5 169.138
R31141 por_dig_0._036_.n1 por_dig_0._036_.t3 168.185
R31142 por_dig_0._036_.n3 por_dig_0._036_.t4 160.709
R31143 por_dig_0._036_ por_dig_0._036_.n6 159.68
R31144 por_dig_0._036_.n4 por_dig_0._036_.n3 152
R31145 por_dig_0._036_.n2 por_dig_0._036_.n1 152
R31146 por_dig_0._036_.n8 por_dig_0._036_.n0 91.5647
R31147 por_dig_0._036_.n9 por_dig_0._036_.n8 88.9533
R31148 por_dig_0._036_.n7 por_dig_0._036_ 74.3729
R31149 por_dig_0._036_.n8 por_dig_0._036_ 27.7737
R31150 por_dig_0._036_.n0 por_dig_0._036_.t0 24.9236
R31151 por_dig_0._036_.n0 por_dig_0._036_.t2 24.9236
R31152 por_dig_0._036_.n5 por_dig_0._036_.n4 20.243
R31153 por_dig_0._036_.n5 por_dig_0._036_ 17.6384
R31154 por_dig_0._036_.n7 por_dig_0._036_.n5 16.1023
R31155 por_dig_0._036_ por_dig_0._036_.n2 13.3631
R31156 por_dig_0._036_ por_dig_0._036_.n9 7.54721
R31157 por_dig_0._036_ por_dig_0._036_.n7 3.0302
R31158 por_dig_0._036_.n4 por_dig_0._036_ 2.13383
R31159 por_dig_0._036_.n2 por_dig_0._036_ 1.82907
R31160 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[4].n1 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[4].n0 873.303
R31161 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[4] por_ana_0.rstring_mux_0.vtrip_decoded_avdd[4].n1 585
R31162 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[4].t0 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[4] 511.971
R31163 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[4].n2 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[4].t3 384.704
R31164 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[4].n2 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[4].t4 384.226
R31165 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[4] por_ana_0.rstring_mux_0.vtrip_decoded_avdd[4].t1 155.607
R31166 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[4] por_ana_0.rstring_mux_0.vtrip_decoded_avdd[4].n3 153.165
R31167 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[4].n1 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[4].t0 147.756
R31168 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[4].n3 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[4].t2 114.031
R31169 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[4].n3 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[4].t5 81.5883
R31170 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[4].n5 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[4] 36.5006
R31171 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[4] por_ana_0.rstring_mux_0.vtrip_decoded_avdd[4].n4 13.8005
R31172 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[4] por_ana_0.rstring_mux_0.vtrip_decoded_avdd[4].n2 9.72818
R31173 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[4].n0 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[4] 8.85549
R31174 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[4].n4 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[4] 7.97972
R31175 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[4].n4 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[4] 7.97972
R31176 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[4].n5 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[4] 7.49318
R31177 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[4] por_ana_0.rstring_mux_0.vtrip_decoded_avdd[4].n0 4.05904
R31178 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[4] por_ana_0.rstring_mux_0.vtrip_decoded_avdd[4].n5 4.05904
R31179 por_ana_0.ibias_gen_0.ena_b.n1 por_ana_0.ibias_gen_0.ena_b.t5 400.171
R31180 por_ana_0.ibias_gen_0.ena_b.n1 por_ana_0.ibias_gen_0.ena_b.t6 392.344
R31181 por_ana_0.ibias_gen_0.ena_b.n2 por_ana_0.ibias_gen_0.ena_b.t4 100.382
R31182 por_ana_0.ibias_gen_0.ena_b.n2 por_ana_0.ibias_gen_0.ena_b.t7 99.138
R31183 por_ana_0.ibias_gen_0.ena_b.n4 por_ana_0.ibias_gen_0.ena_b.n0 46.3607
R31184 por_ana_0.ibias_gen_0.ena_b.n5 por_ana_0.ibias_gen_0.ena_b.n4 18.3117
R31185 por_ana_0.ibias_gen_0.ena_b.n3 por_ana_0.ibias_gen_0.ena_b.n1 7.02575
R31186 por_ana_0.ibias_gen_0.ena_b.n3 por_ana_0.ibias_gen_0.ena_b.n2 6.71284
R31187 por_ana_0.ibias_gen_0.ena_b.n0 por_ana_0.ibias_gen_0.ena_b.t0 5.5395
R31188 por_ana_0.ibias_gen_0.ena_b.n0 por_ana_0.ibias_gen_0.ena_b.t2 5.5395
R31189 por_ana_0.ibias_gen_0.ena_b.n4 por_ana_0.ibias_gen_0.ena_b.n3 5.00928
R31190 por_ana_0.ibias_gen_0.ena_b.t1 por_ana_0.ibias_gen_0.ena_b.n5 3.3065
R31191 por_ana_0.ibias_gen_0.ena_b.n5 por_ana_0.ibias_gen_0.ena_b.t3 3.3065
R31192 force_ena_rc_osc.n0 force_ena_rc_osc.t2 260.322
R31193 force_ena_rc_osc.n0 force_ena_rc_osc.t3 175.169
R31194 force_ena_rc_osc.n1 force_ena_rc_osc.n0 153.165
R31195 force_ena_rc_osc.n3 force_ena_rc_osc.n2 78.4889
R31196 force_ena_rc_osc.n4 force_ena_rc_osc.n3 21.723
R31197 force_ena_rc_osc force_ena_rc_osc.n1 17.7948
R31198 force_ena_rc_osc.n2 force_ena_rc_osc.t1 16.5305
R31199 force_ena_rc_osc.n2 force_ena_rc_osc.t0 16.5305
R31200 force_ena_rc_osc.n3 force_ena_rc_osc 5.28592
R31201 force_ena_rc_osc.n1 force_ena_rc_osc 3.29747
R31202 force_ena_rc_osc.n4 force_ena_rc_osc 0.435642
R31203 force_ena_rc_osc force_ena_rc_osc.n4 0.290725
R31204 por_ana_0.ibias_gen_0.ve.t1 por_ana_0.ibias_gen_0.ve.n0 31123.1
R31205 por_ana_0.ibias_gen_0.ve.n1 por_ana_0.ibias_gen_0.ve.t1 146.25
R31206 por_ana_0.ibias_gen_0.ve.n5 por_ana_0.ibias_gen_0.ve.n4 62.2607
R31207 por_ana_0.ibias_gen_0.ve.n4 por_ana_0.ibias_gen_0.ve.n3 21.4545
R31208 por_ana_0.ibias_gen_0.ve.n4 por_ana_0.ibias_gen_0.ve.n2 20.7025
R31209 por_ana_0.ibias_gen_0.ve.n5 por_ana_0.ibias_gen_0.ve.n1 8.57525
R31210 por_ana_0.sky130_fd_pr__rf_pnp_05v5_W0p68L0p68_0.Emitter por_ana_0.ibias_gen_0.ve.n5 6.71196
R31211 por_ana_0.ibias_gen_0.ve.n3 por_ana_0.ibias_gen_0.ve.t3 3.3065
R31212 por_ana_0.ibias_gen_0.ve.n3 por_ana_0.ibias_gen_0.ve.t0 3.3065
R31213 por_ana_0.ibias_gen_0.ve.n2 por_ana_0.ibias_gen_0.ve.t2 3.3065
R31214 por_ana_0.ibias_gen_0.ve.n2 por_ana_0.ibias_gen_0.ve.t4 3.3065
R31215 por_ana_0.sky130_fd_pr__rf_pnp_05v5_W0p68L0p68_0.Emitter por_ana_0.ibias_gen_0.ve.n1 1.86379
R31216 por_ana_0.rstring_mux_0.vtrip4.n5 por_ana_0.rstring_mux_0.vtrip4.n3 50.7022
R31217 por_ana_0.rstring_mux_0.vtrip4.n2 por_ana_0.rstring_mux_0.vtrip4.n0 50.7022
R31218 por_ana_0.rstring_mux_0.vtrip4.n7 por_ana_0.rstring_mux_0.vtrip4.n6 24.0569
R31219 por_ana_0.rstring_mux_0.vtrip4.n6 por_ana_0.rstring_mux_0.vtrip4.n2 14.0584
R31220 por_ana_0.rstring_mux_0.vtrip4.n5 por_ana_0.rstring_mux_0.vtrip4.n4 13.8791
R31221 por_ana_0.rstring_mux_0.vtrip4.n2 por_ana_0.rstring_mux_0.vtrip4.n1 13.8791
R31222 por_ana_0.rstring_mux_0.vtrip4.n7 por_ana_0.rstring_mux_0.vtrip4.t7 10.6303
R31223 por_ana_0.rstring_mux_0.vtrip4.n3 por_ana_0.rstring_mux_0.vtrip4.t6 5.5395
R31224 por_ana_0.rstring_mux_0.vtrip4.n3 por_ana_0.rstring_mux_0.vtrip4.t5 5.5395
R31225 por_ana_0.rstring_mux_0.vtrip4.n0 por_ana_0.rstring_mux_0.vtrip4.t4 5.5395
R31226 por_ana_0.rstring_mux_0.vtrip4.n0 por_ana_0.rstring_mux_0.vtrip4.t3 5.5395
R31227 por_ana_0.rstring_mux_0.vtrip4.n6 por_ana_0.rstring_mux_0.vtrip4.n5 3.33746
R31228 por_ana_0.rstring_mux_0.vtrip4.n4 por_ana_0.rstring_mux_0.vtrip4.t9 3.3065
R31229 por_ana_0.rstring_mux_0.vtrip4.n4 por_ana_0.rstring_mux_0.vtrip4.t8 3.3065
R31230 por_ana_0.rstring_mux_0.vtrip4.n1 por_ana_0.rstring_mux_0.vtrip4.t2 3.3065
R31231 por_ana_0.rstring_mux_0.vtrip4.n1 por_ana_0.rstring_mux_0.vtrip4.t1 3.3065
R31232 por_ana_0.rstring_mux_0.vtrip4 por_ana_0.rstring_mux_0.vtrip4.t0 0.769662
R31233 por_ana_0.rstring_mux_0.vtrip4 por_ana_0.rstring_mux_0.vtrip4.n7 0.0563195
R31234 por_dig_0.otrip_decoded[0].n2 por_dig_0.otrip_decoded[0].n1 289.849
R31235 por_dig_0.otrip_decoded[0].n3 por_dig_0.otrip_decoded[0].t4 186.374
R31236 por_dig_0.otrip_decoded[0].n9 por_dig_0.otrip_decoded[0].n8 185
R31237 por_dig_0.otrip_decoded[0].n3 por_dig_0.otrip_decoded[0].t5 170.308
R31238 por_dig_0.otrip_decoded[0].n4 por_dig_0.otrip_decoded[0] 154.56
R31239 por_dig_0.otrip_decoded[0].n5 por_dig_0.otrip_decoded[0].n4 153.462
R31240 por_dig_0.otrip_decoded[0].n4 por_dig_0.otrip_decoded[0].n3 101.513
R31241 por_dig_0.otrip_decoded[0] por_dig_0.otrip_decoded[0].n9 81.3181
R31242 por_dig_0.otrip_decoded[0].n0 por_dig_0.otrip_decoded[0].n6 40.7097
R31243 por_dig_0.otrip_decoded[0].n1 por_dig_0.otrip_decoded[0].t2 26.5955
R31244 por_dig_0.otrip_decoded[0].n1 por_dig_0.otrip_decoded[0].t3 26.5955
R31245 por_dig_0.otrip_decoded[0].n8 por_dig_0.otrip_decoded[0].t1 24.9236
R31246 por_dig_0.otrip_decoded[0].n8 por_dig_0.otrip_decoded[0].t0 24.9236
R31247 por_dig_0.otrip_decoded[0].n7 por_dig_0.otrip_decoded[0] 18.234
R31248 por_dig_0.otrip_decoded[0] por_dig_0.otrip_decoded[0].n2 9.15439
R31249 por_dig_0.otrip_decoded[0].n2 por_dig_0.otrip_decoded[0] 7.71085
R31250 por_dig_0.otrip_decoded[0].n6 por_dig_0.otrip_decoded[0].n5 4.96991
R31251 por_dig_0.otrip_decoded[0].n7 por_dig_0.otrip_decoded[0] 4.26717
R31252 por_dig_0.otrip_decoded[0] por_dig_0.otrip_decoded[0].n0 3.85318
R31253 por_dig_0.otrip_decoded[0].n5 por_dig_0.otrip_decoded[0] 3.46403
R31254 por_dig_0.otrip_decoded[0].n6 por_dig_0.otrip_decoded[0] 2.71109
R31255 por_dig_0.otrip_decoded[0].n0 por_dig_0.otrip_decoded[0] 1.14782
R31256 por_dig_0.otrip_decoded[0].n0 por_dig_0.otrip_decoded[0] 1.07133
R31257 por_dig_0.otrip_decoded[0].n9 por_dig_0.otrip_decoded[0].n7 1.00442
R31258 por_dig_0.otrip_decoded[0].n0 por_dig_0.otrip_decoded[0] 0.973714
R31259 ibg_200n.n0 ibg_200n.t1 51.3525
R31260 ibg_200n ibg_200n.n0 41.4648
R31261 ibg_200n.n0 ibg_200n.t0 22.0614
R31262 startup_timed_out.n2 startup_timed_out.n1 585
R31263 startup_timed_out.n1 startup_timed_out.n0 585
R31264 startup_timed_out.n4 startup_timed_out.n3 185
R31265 startup_timed_out startup_timed_out.n2 79.5613
R31266 startup_timed_out.n1 startup_timed_out.t3 26.5955
R31267 startup_timed_out.n1 startup_timed_out.t2 26.5955
R31268 startup_timed_out.n3 startup_timed_out.t1 24.9236
R31269 startup_timed_out.n3 startup_timed_out.t0 24.9236
R31270 startup_timed_out startup_timed_out.n4 17.243
R31271 startup_timed_out.n0 startup_timed_out 13.3025
R31272 startup_timed_out.n2 startup_timed_out 7.02795
R31273 startup_timed_out.n0 startup_timed_out 3.76521
R31274 startup_timed_out.n4 startup_timed_out 3.26325
R31275 otrip[0].n0 otrip[0].t3 323.55
R31276 otrip[0].n0 otrip[0].t2 195.017
R31277 otrip[0].n1 otrip[0].n0 152
R31278 otrip[0].n4 otrip[0].n3 74.301
R31279 otrip[0].n5 otrip[0].n2 17.0381
R31280 otrip[0].n3 otrip[0].t1 16.5305
R31281 otrip[0].n3 otrip[0].t0 16.5305
R31282 otrip[0].n5 otrip[0].n4 11.325
R31283 otrip[0].n2 otrip[0] 6.7304
R31284 otrip[0] otrip[0].n5 2.95139
R31285 otrip[0].n1 otrip[0] 1.45205
R31286 otrip[0].n2 otrip[0].n1 0.792253
R31287 otrip[0].n4 otrip[0] 0.729532
R31288 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[5].n1 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[5].n0 873.303
R31289 por_ana_0.sky130_fd_sc_hvl__lsbuflv2hv_1_0[1|6].X por_ana_0.rstring_mux_0.vtrip_decoded_avdd[5].n1 585
R31290 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[5].t0 por_ana_0.sky130_fd_sc_hvl__lsbuflv2hv_1_0[1|6].X 511.971
R31291 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[5].n2 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[5].t5 384.704
R31292 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[5].n2 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[5].t4 384.226
R31293 por_ana_0.sky130_fd_sc_hvl__lsbuflv2hv_1_0[1|6].X por_ana_0.rstring_mux_0.vtrip_decoded_avdd[5].t1 155.607
R31294 por_ana_0.rstring_mux_0.sky130_fd_sc_hvl__inv_1_0[13].A por_ana_0.rstring_mux_0.vtrip_decoded_avdd[5].n3 153.165
R31295 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[5].n1 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[5].t0 147.756
R31296 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[5].n3 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[5].t3 114.031
R31297 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[5].n3 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[5].t2 81.5883
R31298 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[5].n6 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[5].n5 39.8143
R31299 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[5].n5 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[5].n4 13.8005
R31300 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[5].n5 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[5].n2 9.66019
R31301 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[5].n0 por_ana_0.sky130_fd_sc_hvl__lsbuflv2hv_1_0[1|6].X 8.85549
R31302 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[5].n4 por_ana_0.rstring_mux_0.sky130_fd_sc_hvl__inv_1_0[13].A 7.97972
R31303 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[5].n4 por_ana_0.rstring_mux_0.sky130_fd_sc_hvl__inv_1_0[13].A 7.97972
R31304 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[5].n6 por_ana_0.sky130_fd_sc_hvl__lsbuflv2hv_1_0[1|6].X 7.49318
R31305 por_ana_0.sky130_fd_sc_hvl__lsbuflv2hv_1_0[1|6].X por_ana_0.rstring_mux_0.vtrip_decoded_avdd[5].n0 4.05904
R31306 por_ana_0.sky130_fd_sc_hvl__lsbuflv2hv_1_0[1|6].X por_ana_0.rstring_mux_0.vtrip_decoded_avdd[5].n6 4.05904
R31307 force_dis_rc_osc.n0 force_dis_rc_osc.t2 260.322
R31308 force_dis_rc_osc.n0 force_dis_rc_osc.t3 175.169
R31309 force_dis_rc_osc.n1 force_dis_rc_osc.n0 153.385
R31310 force_dis_rc_osc.n3 force_dis_rc_osc.n2 70.8209
R31311 force_dis_rc_osc force_dis_rc_osc.n1 27.1383
R31312 force_dis_rc_osc.n4 force_dis_rc_osc.n3 16.9931
R31313 force_dis_rc_osc.n2 force_dis_rc_osc.t0 16.5305
R31314 force_dis_rc_osc.n2 force_dis_rc_osc.t1 16.5305
R31315 force_dis_rc_osc.n3 force_dis_rc_osc 12.6078
R31316 force_dis_rc_osc.n1 force_dis_rc_osc 2.94104
R31317 force_dis_rc_osc force_dis_rc_osc.n4 0.218658
R31318 force_dis_rc_osc.n4 force_dis_rc_osc 0.129358
R31319 force_pdn.n0 force_pdn.t2 260.322
R31320 force_pdn.n0 force_pdn.t3 175.169
R31321 force_pdn.n1 force_pdn.n0 153.385
R31322 force_pdn.n3 force_pdn.n2 70.9715
R31323 force_pdn.n4 force_pdn.n3 24.0287
R31324 force_pdn force_pdn.n1 18.4167
R31325 force_pdn.n2 force_pdn.t0 16.5305
R31326 force_pdn.n2 force_pdn.t1 16.5305
R31327 force_pdn.n3 force_pdn 5.28592
R31328 force_pdn.n1 force_pdn 2.94104
R31329 force_pdn.n4 force_pdn 0.433683
R31330 force_pdn force_pdn.n4 0.0717833
R31331 por_ana_0.comparator_0.n0.n2 por_ana_0.comparator_0.n0.t7 227.651
R31332 por_ana_0.comparator_0.n0.n2 por_ana_0.comparator_0.n0.t5 227.173
R31333 por_ana_0.comparator_0.n0.n0 por_ana_0.comparator_0.n0.t8 224.037
R31334 por_ana_0.comparator_0.n0.n0 por_ana_0.comparator_0.n0.t6 223.559
R31335 por_ana_0.comparator_0.n0 por_ana_0.comparator_0.n0.n1 205.605
R31336 por_ana_0.comparator_0.n0 por_ana_0.comparator_0.n0.t4 96.5813
R31337 por_ana_0.comparator_0.n0 por_ana_0.comparator_0.n0.n3 70.9612
R31338 por_ana_0.comparator_0.n0.n1 por_ana_0.comparator_0.n0.t1 27.6955
R31339 por_ana_0.comparator_0.n0.n1 por_ana_0.comparator_0.n0.t0 27.6955
R31340 por_ana_0.comparator_0.n0.n3 por_ana_0.comparator_0.n0.t3 16.5305
R31341 por_ana_0.comparator_0.n0.n3 por_ana_0.comparator_0.n0.t2 16.5305
R31342 por_ana_0.comparator_0.n0.n0 por_ana_0.comparator_0.n0.n2 14.4688
R31343 por_ana_0.comparator_0.n0 por_ana_0.comparator_0.n0.n0 10.4432
R31344 por_ana_0.ibias_gen_0.vr.n2 por_ana_0.ibias_gen_0.vr.n0 21.7373
R31345 por_ana_0.ibias_gen_0.vr.n2 por_ana_0.ibias_gen_0.vr.n1 20.4114
R31346 por_ana_0.ibias_gen_0.vr.t4 por_ana_0.ibias_gen_0.vr.n2 17.6029
R31347 por_ana_0.ibias_gen_0.vr.n1 por_ana_0.ibias_gen_0.vr.t0 3.3065
R31348 por_ana_0.ibias_gen_0.vr.n1 por_ana_0.ibias_gen_0.vr.t3 3.3065
R31349 por_ana_0.ibias_gen_0.vr.n0 por_ana_0.ibias_gen_0.vr.t2 3.3065
R31350 por_ana_0.ibias_gen_0.vr.n0 por_ana_0.ibias_gen_0.vr.t1 3.3065
R31351 por_ana_0.comparator_0.ibias.n0 por_ana_0.comparator_0.ibias.t3 233.487
R31352 por_ana_0.comparator_0.ibias.n1 por_ana_0.comparator_0.ibias.n0 105.507
R31353 por_ana_0.comparator_0.ibias.n0 por_ana_0.comparator_0.ibias.t0 88.1251
R31354 por_ana_0.comparator_0.ibias.t2 por_ana_0.comparator_0.ibias.n1 5.5395
R31355 por_ana_0.comparator_0.ibias.n1 por_ana_0.comparator_0.ibias.t1 5.5395
R31356 por_ana_0.comparator_1.vn.n1 por_ana_0.comparator_1.vn.t2 234.096
R31357 por_ana_0.comparator_1.vn.n2 por_ana_0.comparator_1.vn.t1 94.5098
R31358 por_ana_0.comparator_1.vn.n1 por_ana_0.comparator_1.vn.t0 87.5075
R31359 por_ana_0.comparator_1.vn.n0 por_ana_0.comparator_1.vn.n3 66.4612
R31360 por_ana_0.comparator_1.vn.n3 por_ana_0.comparator_1.vn.t6 16.5305
R31361 por_ana_0.comparator_1.vn.n3 por_ana_0.comparator_1.vn.t4 16.5305
R31362 por_ana_0.comparator_1.vn.n0 por_ana_0.comparator_1.vn.t7 16.2067
R31363 por_ana_0.comparator_1.vn.n0 por_ana_0.comparator_1.vn.t3 13.954
R31364 por_ana_0.comparator_1.vn.n0 por_ana_0.comparator_1.vn.t5 11.7013
R31365 por_ana_0.comparator_1.vn.n0 por_ana_0.comparator_1.vn.t8 11.7013
R31366 por_ana_0.comparator_1.vn por_ana_0.comparator_1.vn.n0 11.4244
R31367 por_ana_0.comparator_1.vn por_ana_0.comparator_1.vn.n2 10.7596
R31368 por_ana_0.comparator_1.vn.n2 por_ana_0.comparator_1.vn.n1 8.74658
R31369 por_ana_0.rstring_mux_0.vtrip1.n5 por_ana_0.rstring_mux_0.vtrip1.n3 50.7022
R31370 por_ana_0.rstring_mux_0.vtrip1.n2 por_ana_0.rstring_mux_0.vtrip1.n0 50.7022
R31371 por_ana_0.rstring_mux_0.vtrip1.n6 por_ana_0.rstring_mux_0.vtrip1.n5 14.0767
R31372 por_ana_0.rstring_mux_0.vtrip1.n5 por_ana_0.rstring_mux_0.vtrip1.n4 13.8791
R31373 por_ana_0.rstring_mux_0.vtrip1.n2 por_ana_0.rstring_mux_0.vtrip1.n1 13.8791
R31374 por_ana_0.rstring_mux_0.vtrip1.t4 por_ana_0.rstring_mux_0.vtrip1.n7 10.5857
R31375 por_ana_0.rstring_mux_0.vtrip1.n7 por_ana_0.rstring_mux_0.vtrip1.t7 10.5847
R31376 por_ana_0.rstring_mux_0.vtrip1.n7 por_ana_0.rstring_mux_0.vtrip1.n6 5.61984
R31377 por_ana_0.rstring_mux_0.vtrip1.n3 por_ana_0.rstring_mux_0.vtrip1.t6 5.5395
R31378 por_ana_0.rstring_mux_0.vtrip1.n3 por_ana_0.rstring_mux_0.vtrip1.t5 5.5395
R31379 por_ana_0.rstring_mux_0.vtrip1.n0 por_ana_0.rstring_mux_0.vtrip1.t1 5.5395
R31380 por_ana_0.rstring_mux_0.vtrip1.n0 por_ana_0.rstring_mux_0.vtrip1.t0 5.5395
R31381 por_ana_0.rstring_mux_0.vtrip1.n6 por_ana_0.rstring_mux_0.vtrip1.n2 3.9186
R31382 por_ana_0.rstring_mux_0.vtrip1.n4 por_ana_0.rstring_mux_0.vtrip1.t9 3.3065
R31383 por_ana_0.rstring_mux_0.vtrip1.n4 por_ana_0.rstring_mux_0.vtrip1.t8 3.3065
R31384 por_ana_0.rstring_mux_0.vtrip1.n1 por_ana_0.rstring_mux_0.vtrip1.t3 3.3065
R31385 por_ana_0.rstring_mux_0.vtrip1.n1 por_ana_0.rstring_mux_0.vtrip1.t2 3.3065
R31386 itest itest.n0 80.4227
R31387 itest.n0 itest.t0 5.5395
R31388 itest.n0 itest.t1 5.5395
C0 por_dig_0.cnt_st\[2\] por_dig_0.cnt_st\[3\] 0.192025f
C1 por_dig_0._025_ por_dig_0.cnt_por\[6\] 0.174846f
C2 a_31908_32909# por_dig_0.net28 0.131599f
C3 a_36880_32915# por_dig_0._002_ 0.609716f
C4 a_29126_6535# a_29882_6535# 0.296258f
C5 a_30070_21903# dvdd 0.176016f
C6 por_ana_0.rstring_mux_0.vtrip_decoded_b_avdd[0] avss 0.36282f
C7 por_ana_0.rstring_mux_0.otrip_decoded_avdd[7] por_ana_0.rstring_mux_0.otrip_decoded_b_avdd[7] 0.572384f
C8 por_ana_0.schmitt_trigger_0.in por_ana_0.rstring_mux_0.otrip_decoded_avdd[3] 0.117015f
C9 a_34418_6535# avss 0.466333f
C10 por_dig_0.net20 a_36381_36691# 0.22392f
C11 a_34510_31277# a_34746_31277# 0.22264f
C12 por_dig_0.net12 dvdd 0.505426f
C13 por_dig_0.net26 dvdd 1.09793f
C14 por_ana_0.rstring_mux_0.otrip_decoded_b_avdd[5] avdd 0.903548f
C15 a_27690_22973# a_28897_22637# 0.28899f
C16 por_dig_0._010_ a_32885_33275# 0.183223f
C17 a_31814_22885# dvdd 0.380879f
C18 por_dig_0.net28 por_dig_0.net8 0.139479f
C19 por_dig_0.net18 por_dig_0.otrip_decoded[5] 0.20913f
C20 por_dig_0.otrip_decoded[4] por_dig_0.otrip_decoded[3] 0.132744f
C21 a_25846_21903# avdd 0.143952f
C22 a_20044_27844# a_20800_27844# 0.296258f
C23 por_dig_0.clknet_1_0__leaf_osc_ck a_31360_31827# 0.333709f
C24 por_dig_0._004_ a_36696_30739# 0.352282f
C25 a_26802_33372# avdd 0.419619f
C26 a_24159_23593# dvdd 0.105303f
C27 a_19676_13935# avss 0.465068f
C28 a_29802_22973# avdd 0.863791f
C29 por_dig_0._007_ a_32610_35603# 0.141526f
C30 por_ana_0.rstring_mux_0.otrip_decoded_avdd[0] por_ana_0.rstring_mux_0.vtrip0 0.50883f
C31 por_dig_0.net24 a_32188_30739# 0.302829f
C32 por_dig_0.net22 por_dig_0._026_ 0.857243f
C33 a_34719_21859# a_34294_21903# 0.460766f
C34 por_dig_0.clknet_1_1__leaf_osc_ck por_dig_0._052_ 0.301336f
C35 a_32004_30189# dvdd 0.239676f
C36 a_32906_36179# a_33256_36551# 0.228946f
C37 por_dig_0.cnt_por\[10\] a_36476_30163# 0.29859f
C38 por_dig_0.net18 dvdd 0.527f
C39 a_14384_13935# a_15140_13935# 0.296258f
C40 por_ana_0.rstring_mux_0.vtrip_decoded_b_avdd[7] avss 0.479446f
C41 por_dig_0._033_ osc_ck 0.118226f
C42 por_dig_0.net27 por_dig_0.cnt_por\[10\] 0.396309f
C43 por_dig_0._018_ dvdd 0.647818f
C44 a_31615_33705# a_31893_33721# 0.125324f
C45 a_38242_31251# dvdd 0.251025f
C46 por_dig_0._005_ a_35921_35629# 0.15568f
C47 por_dig_0.cnt_st\[2\] por_dig_0._030_ 0.521593f
C48 por_dig_0.otrip_decoded[3] a_23366_24619# 0.207798f
C49 por_ana_0.rstring_mux_0.vtrip_decoded_b_avdd[4] avdd 0.903548f
C50 a_22047_21859# dvdd 0.104499f
C51 por_ana_0.vl por_dig_0.otrip_decoded[2] 1.02322f
C52 por_dig_0.force_pdnb por_dig_0.otrip_decoded[6] 0.10144f
C53 por_dig_0.net20 por_dig_0.net23 0.46167f
C54 por_ana_0.sky130_fd_sc_hvl__inv_1_0.A porb 0.423857f
C55 a_38974_34693# por_dig_0.net31 0.135862f
C56 por_ana_0.sky130_fd_sc_hvl__inv_1_0.A por 0.473758f
C57 a_29126_6535# avss 0.466333f
C58 por_ana_0.comparator_1.vnn vin 0.848157f
C59 a_34934_28013# a_35111_28013# 0.159555f
C60 por_dig_0.cnt_por\[5\] a_34387_32909# 0.119299f
C61 a_36831_23593# dvdd 0.107699f
C62 a_36880_33453# dvdd 0.425756f
C63 a_36880_33453# a_37046_33453# 0.906454f
C64 por_dig_0.cnt_por\[9\] a_35000_31795# 0.229052f
C65 por_dig_0.cnt_por\[1\] a_35500_35629# 0.183278f
C66 por_dig_0._048_ por_dig_0._017_ 0.173152f
C67 por_ana_0.rstring_mux_0.otrip_decoded_avdd[2] por_ana_0.rstring_mux_0.otrip_decoded_b_avdd[1] 0.155388f
C68 a_14384_13935# avss 0.465096f
C69 a_2543_22912# a_3299_22912# 0.296258f
C70 por_dig_0.cnt_st\[0\] a_38956_32339# 0.176697f
C71 a_39888_24823# avdd 0.538496f
C72 por_dig_0.net25 a_36480_31251# 0.305396f
C73 por_ana_0.rc_osc_0.m dvdd 2.38557f
C74 por_dig_0.cnt_por\[0\] a_35592_36286# 0.136001f
C75 a_33269_31111# dvdd 0.302575f
C76 por_ana_0.dcomp3v3 avdd 6.668f
C77 por_ana_0.comparator_1.vnn por_ana_0.comparator_1.n0 0.42769f
C78 por_dig_0.net26 a_31893_31545# 0.263898f
C79 a_27590_24619# avdd 0.206171f
C80 a_34633_36147# dvdd 0.200658f
C81 por_dig_0._042_ por_dig_0._003_ 0.231298f
C82 force_ena_rc_osc pwup_filt 0.28199f
C83 a_37614_32883# dvdd 0.203359f
C84 por_ana_0.rstring_mux_0.otrip_decoded_avdd[1] por_ana_0.rstring_mux_0.otrip_decoded_b_avdd[0] 0.176375f
C85 por_ana_0.rc_osc_0.in avdd 1.35364f
C86 por_dig_0.net24 a_37584_35389# 0.280448f
C87 a_22322_6535# a_23078_6535# 0.296258f
C88 por_dig_0._004_ a_37117_31099# 0.17705f
C89 avss isrc_sel 0.230477f
C90 a_22322_6535# avss 0.466333f
C91 por_dig_0.net25 a_37430_30707# 0.16857f
C92 a_32358_28013# a_32535_28013# 0.159555f
C93 por_ana_0.rstring_mux_0.otrip_decoded_b_avdd[2] vin 0.34139f
C94 a_34796_13935# a_35552_13935# 0.296258f
C95 por_ana_0.rstring_mux_0.otrip_decoded_avdd[7] avss 1.37218f
C96 por_dig_0._047_ a_32794_33971# 0.237501f
C97 por_dig_0.net21 a_38957_32883# 0.146155f
C98 por_dig_0.net23 a_36564_32339# 0.183648f
C99 por_dig_0.por_unbuf por_dig_0.otrip_decoded[2] 0.196756f
C100 por_ana_0.vl avss 1.58811f
C101 por_dig_0.clknet_1_0__leaf_osc_ck a_34098_30707# 1.85359f
C102 a_14752_27844# a_15508_27844# 0.296258f
C103 por_dig_0.net24 por_dig_0.cnt_por\[6\] 0.662782f
C104 por_dig_0._009_ dvdd 0.475717f
C105 por_dig_0._053_ dvdd 0.168313f
C106 por_dig_0.osc_ena por_dig_0.otrip_decoded[5] 0.105641f
C107 por_ana_0.comparator_1.vm por_ana_0.comparator_1.n0 2.58153f
C108 a_39728_31527# dvdd 0.249576f
C109 por_dig_0._039_ dvdd 0.569627f
C110 a_36414_32909# dvdd 0.200226f
C111 por_dig_0.cnt_por\[1\] por_dig_0._049_ 0.175577f
C112 a_25478_24619# a_25578_24707# 0.40546f
C113 por_dig_0.clknet_0_osc_ck por_dig_0._018_ 0.632467f
C114 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[2] dvdd 0.279976f
C115 a_35666_35629# a_36016_35629# 0.206984f
C116 por_dig_0.net7 por_dig_0.net17 0.423111f
C117 por_dig_0._035_ por_dig_0._036_ 0.754854f
C118 por_ana_0.rstring_mux_0.otrip_decoded_avdd[3] por_ana_0.rstring_mux_0.otrip_decoded_b_avdd[2] 0.155546f
C119 por_dig_0.net25 a_37706_30431# 0.188233f
C120 avdd otrip[1] 0.225768f
C121 avdd dcomp 0.474805f
C122 por_ana_0.rstring_mux_0.otrip_decoded_avdd[4] avss 1.34995f
C123 por_dig_0.cnt_st\[0\] por_dig_0.net4 0.845085f
C124 por_dig_0.net24 a_33256_35463# 0.156236f
C125 por_dig_0.net9 dvdd 0.369411f
C126 por_dig_0.osc_ena dvdd 7.45726f
C127 a_19094_3138# osc_ck 0.152841f
C128 a_32188_30739# a_32354_30739# 0.614266f
C129 por_ana_0.rstring_mux_0.otrip_decoded_avdd[4] por_ana_0.rstring_mux_0.vtrip4 0.533298f
C130 a_34357_33427# dvdd 0.166696f
C131 por_dig_0._031_ dvdd 0.75531f
C132 a_34728_30189# dvdd 0.203526f
C133 a_17030_6535# avss 0.466333f
C134 por_dig_0.force_pdnb avdd 0.500678f
C135 a_21254_22885# avdd 0.194488f
C136 por_dig_0.cnt_por\[4\] por_dig_0.cnt_por\[8\] 0.119375f
C137 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[2] por_ana_0.dcomp3v3uv 0.359441f
C138 a_24159_21859# a_23734_21903# 0.460766f
C139 a_32740_35091# a_33821_35463# 0.102325f
C140 a_33474_35059# a_33256_35463# 0.209641f
C141 por_dig_0.net34 a_38146_31429# 0.198254f
C142 a_32610_35603# dvdd 0.21733f
C143 por_dig_0.otrip_decoded[2] a_23366_22885# 0.277476f
C144 por_dig_0.net27 a_36328_29645# 0.219834f
C145 a_35390_31277# a_36305_31277# 0.125324f
C146 por_dig_0.net21 dvdd 0.620271f
C147 a_38150_24619# avdd 0.206179f
C148 por_dig_0._025_ por_dig_0._019_ 0.216424f
C149 por_dig_0.net25 dvdd 2.96037f
C150 por_dig_0.net6 a_35030_28557# 0.107171f
C151 a_20422_35244# avss 0.460284f
C152 a_38250_22973# a_39457_22637# 0.28899f
C153 dvdd porb_h 0.231478f
C154 a_28897_22637# por_ana_0.rstring_mux_0.otrip_decoded_avdd[6] 0.136228f
C155 por_dig_0.net28 dvdd 0.474831f
C156 a_41694_1248# a_41694_492# 0.296258f
C157 por_dig_0.clknet_1_0__leaf_osc_ck a_32464_32915# 0.248686f
C158 por_dig_0.net4 por_dig_0._019_ 0.469127f
C159 por_dig_0.otrip_decoded[2] por_ana_0.rstring_mux_0.otrip_decoded_avdd[1] 0.142991f
C160 por_ana_0.vl ibg_200n 0.329198f
C161 por_dig_0.net17 dvdd 0.21063f
C162 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[3] por_ana_0.rstring_mux_0.vtrip_decoded_avdd[2] 1.78143f
C163 a_31566_32909# dvdd 0.2998f
C164 por_dig_0.otrip_decoded[7] por_dig_0.otrip_decoded[3] 4.68124f
C165 por_dig_0.por_unbuf avss 0.800925f
C166 a_39070_34515# a_39328_34515# 0.22264f
C167 por_dig_0.net24 a_31932_33595# 0.507417f
C168 a_33752_28013# por_dig_0.otrip_decoded[2] 0.184193f
C169 a_34719_23593# a_34294_23637# 0.460766f
C170 por_dig_0._046_ dvdd 0.686901f
C171 por_dig_0.net24 por_dig_0._011_ 0.210945f
C172 por_dig_0._023_ a_35040_34317# 0.113663f
C173 a_31526_31827# dvdd 0.360559f
C174 a_37064_34003# a_37580_34375# 0.110816f
C175 a_17030_6535# a_17786_6535# 0.296258f
C176 por_dig_0.clknet_1_1__leaf_osc_ck por_dig_0._048_ 0.189415f
C177 por_dig_0.otrip_decoded[0] dvdd 0.843312f
C178 avdd force_short_oneshot 0.65973f
C179 por_dig_0.por_unbuf vbg_1v2 0.332056f
C180 por_ana_0.rstring_mux_0.otrip_decoded_avdd[6] vin 0.875633f
C181 a_27590_22885# a_27958_21903# 0.138963f
C182 dvdd startup_timed_out 0.63296f
C183 a_29504_13935# a_30260_13935# 0.296258f
C184 a_34294_21903# dvdd 0.176016f
C185 dvdd osc_ck 3.72227f
C186 por_dig_0.net7 a_35130_28673# 0.303836f
C187 por_dig_0.net16 dvdd 0.489588f
C188 por_dig_0._008_ a_32740_35091# 0.22f
C189 por_dig_0._009_ a_35573_33721# 0.762822f
C190 a_25495_33620# a_25595_33708# 0.40546f
C191 por_dig_0.net26 a_32651_31643# 0.161562f
C192 a_31802_32909# por_dig_0.clknet_1_0__leaf_osc_ck 0.11284f
C193 a_34746_31277# a_34852_31277# 0.419086f
C194 por_dig_0._034_ a_35666_35629# 0.31508f
C195 por_dig_0.net20 por_dig_0.cnt_por\[1\] 0.229286f
C196 a_15130_35244# avss 0.460284f
C197 por_dig_0.net18 a_37156_28013# 0.169992f
C198 por_dig_0.net24 por_dig_0.cnt_por\[5\] 0.574351f
C199 a_30070_21903# avdd 0.143952f
C200 por_dig_0.cnt_rsb dvdd 0.681658f
C201 por_ana_0.rstring_mux_0.otrip_decoded_avdd[5] por_ana_0.rstring_mux_0.otrip_decoded_avdd[4] 1.15427f
C202 a_20422_35244# a_21178_35244# 0.296258f
C203 por_dig_0._032_ a_37789_31821# 0.142553f
C204 a_30495_23593# a_30070_23637# 0.460766f
C205 por_dig_0._039_ por_dig_0.cnt_st\[1\] 0.268975f
C206 a_5189_15512# a_5945_15512# 0.296258f
C207 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[2] por_ana_0.rstring_mux_0.vtrip_decoded_b_avdd[2] 0.5727f
C208 por_dig_0._028_ por_dig_0._014_ 0.118155f
C209 a_31814_22885# avdd 0.207177f
C210 por_dig_0.net24 a_32922_30707# 0.167039f
C211 a_32233_33819# dvdd 0.142103f
C212 a_39887_23089# a_39887_21959# 0.170258f
C213 por_ana_0.rstring_mux_0.otrip_decoded_avdd[1] avss 1.63066f
C214 por_ana_0.rstring_mux_0.vtrip0 a_24968_13935# 0.137908f
C215 a_35666_35629# dvdd 0.413326f
C216 a_32906_36179# a_33821_36551# 0.117156f
C217 por_dig_0.net24 a_33256_36551# 0.15503f
C218 a_24159_23593# avdd 0.607971f
C219 por_dig_0.net4 por_dig_0.net19 0.134109f
C220 a_34026_22973# a_34719_21859# 0.264594f
C221 por_dig_0.net23 a_34633_36147# 0.199822f
C222 a_29802_22973# a_30495_21859# 0.264594f
C223 por_dig_0.net19 por_dig_0._037_ 0.372592f
C224 a_31893_33721# a_31932_33595# 0.822296f
C225 por_dig_0._044_ dvdd 0.228467f
C226 a_35130_28673# dvdd 0.20578f
C227 a_35958_31519# dvdd 0.221161f
C228 por_dig_0.net5 por_dig_0.net17 0.248372f
C229 por_dig_0._011_ a_31893_33721# 0.220244f
C230 por_dig_0.osc_ena por_dig_0.otrip_decoded[6] 0.105247f
C231 por_ana_0.rstring_mux_0.vtrip_decoded_b_avdd[0] por_ana_0.rstring_mux_0.vtrip0 0.190544f
C232 por_dig_0.net8 a_31412_31251# 0.278481f
C233 a_35111_28013# a_35217_28013# 0.313533f
C234 a_37442_6535# a_38198_6535# 0.296258f
C235 a_40247_23627# dvdd 0.485404f
C236 por_dig_0.net4 por_dig_0.cnt_por\[10\] 0.120475f
C237 a_36880_33453# a_37396_33453# 0.115353f
C238 por_dig_0.net19 a_31864_30823# 0.119995f
C239 a_22047_21859# avdd 0.607831f
C240 a_5567_22912# avss 0.474081f
C241 a_31776_29864# force_ena_rc_osc 0.200621f
C242 por_dig_0.cnt_por\[10\] por_dig_0._037_ 0.728205f
C243 a_36038_24619# a_36406_23637# 0.138963f
C244 por_dig_0.clknet_1_1__leaf_osc_ck por_dig_0._047_ 0.774094f
C245 a_37584_35389# a_37409_35463# 0.233657f
C246 a_32906_36179# por_dig_0._052_ 0.279146f
C247 a_36831_23593# avdd 0.607928f
C248 a_36038_24619# a_36138_24707# 0.40546f
C249 a_36696_30739# dvdd 0.472893f
C250 por_dig_0.net24 por_dig_0._019_ 0.218781f
C251 a_23466_24707# a_24159_23593# 0.264594f
C252 por_dig_0.net5 por_dig_0.net16 0.110515f
C253 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[3] por_ana_0.rstring_mux_0.vtrip_decoded_b_avdd[3] 0.572316f
C254 avss pwup_filt 0.2207f
C255 a_28897_24371# avdd 0.420074f
C256 a_37820_13935# avss 0.525755f
C257 por_dig_0._004_ dvdd 0.409945f
C258 por_dig_0.net17 por_dig_0.otrip_decoded[6] 0.253355f
C259 a_31413_32339# por_timed_out 0.162074f
C260 por_dig_0.force_pdnb por_dig_0.otrip_decoded[1] 0.125267f
C261 a_17776_27844# avss 0.460203f
C262 a_38136_33213# dvdd 0.35166f
C263 por_dig_0.cnt_st\[4\] por_dig_0.net34 0.114051f
C264 por_dig_0._015_ a_34496_29645# 0.167821f
C265 a_39268_33453# por_dig_0.net33 0.131009f
C266 a_22700_13935# a_23456_13935# 0.296258f
C267 por_dig_0._028_ a_34496_29645# 0.216958f
C268 por_dig_0.cnt_st\[0\] por_dig_0.cnt_st\[2\] 0.190848f
C269 por_dig_0.cnt_por\[1\] a_34672_35451# 0.230285f
C270 por_dig_0.net14 a_37800_28013# 0.178515f
C271 por_dig_0.net25 a_37952_31037# 0.349798f
C272 a_32535_28013# a_32641_28013# 0.313533f
C273 a_36972_30189# dvdd 0.444924f
C274 avss force_ena_rc_osc 0.295693f
C275 por_dig_0._019_ a_33805_32339# 0.169961f
C276 por_dig_0.clknet_1_0__leaf_osc_ck a_36862_30739# 0.133969f
C277 a_33380_35879# dvdd 0.278713f
C278 a_15130_35244# a_15886_35244# 0.296258f
C279 por_dig_0._002_ a_37301_33275# 0.1701f
C280 por_dig_0.net4 por_dig_0._020_ 0.101152f
C281 por_dig_0.clknet_1_1__leaf_osc_ck a_32740_36179# 0.254076f
C282 por_dig_0._039_ por_dig_0._040_ 0.311871f
C283 por_ana_0.rstring_mux_0.otrip_decoded_avdd[0] vin 0.882514f
C284 por_dig_0.net32 a_34116_31821# 0.129568f
C285 a_35224_31277# por_dig_0._015_ 0.158708f
C286 a_32630_32915# a_32980_33287# 0.21907f
C287 a_25578_24707# a_26785_24371# 0.28899f
C288 a_35666_35629# a_36581_35629# 0.125324f
C289 por_dig_0._032_ por_dig_0.net34 0.3312f
C290 por_dig_0.net25 a_38228_30163# 0.292005f
C291 a_32528_13935# avss 0.465978f
C292 a_32630_32915# dvdd 0.578871f
C293 por_ana_0.rstring_mux_0.vtrip_decoded_b_avdd[6] por_ana_0.rstring_mux_0.vtrip6 0.190544f
C294 por_dig_0.net24 a_33821_35463# 0.278253f
C295 por_ana_0.rstring_mux_0.otrip_decoded_avdd[1] por_ana_0.rstring_mux_0.otrip_decoded_avdd[2] 0.101824f
C296 a_20054_6535# dvdd 0.359438f
C297 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[2] avdd 1.66091f
C298 a_32188_30739# a_32704_31111# 0.105995f
C299 a_32354_30739# a_32922_30707# 0.175891f
C300 por_dig_0.net23 por_dig_0._046_ 0.616632f
C301 a_33364_35085# dvdd 0.143483f
C302 por_dig_0.net4 por_dig_0._010_ 0.197042f
C303 por dcomp 1.35556f
C304 a_8213_15512# avss 0.476371f
C305 por_ana_0.dcomp3v3 por_ana_0.ibias_gen_0.vp1 0.543327f
C306 por_dig_0.net24 por_dig_0.net19 0.135015f
C307 a_35293_30189# dvdd 0.27318f
C308 por_ana_0.rstring_mux_0.otrip_decoded_avdd[6] por_ana_0.rstring_mux_0.otrip_decoded_b_avdd[5] 0.155092f
C309 por_dig_0._031_ a_38936_32159# 0.199995f
C310 a_22561_22637# avdd 0.421965f
C311 por_dig_0._033_ por_dig_0._034_ 0.298747f
C312 por_dig_0.osc_ena avdd 0.721152f
C313 a_32150_6535# a_32906_6535# 0.296258f
C314 por_dig_0.clknet_1_0__leaf_osc_ck a_31728_32365# 0.278472f
C315 por_dig_0.net2 a_31413_29619# 0.108726f
C316 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A porb_h 2.45926f
C317 por_ana_0.sky130_fd_sc_hd__inv_4_3.Y dcomp 1.51717f
C318 a_34265_27987# dvdd 0.261335f
C319 a_39457_24371# avdd 0.418585f
C320 por_dig_0.net21 a_38936_32159# 0.110669f
C321 a_34719_21859# dvdd 0.104499f
C322 por_dig_0.net25 a_37396_33453# 0.164981f
C323 por_ana_0.rstring_mux_0.otrip_decoded_b_avdd[0] avss 0.399825f
C324 a_37800_28013# por_dig_0.otrip_decoded[3] 0.187607f
C325 a_31908_32909# dvdd 0.177412f
C326 a_39328_34515# por_dig_0.cnt_st\[0\] 0.338696f
C327 por_dig_0._033_ dvdd 1.67013f
C328 otrip[1] otrip[2] 3.49315f
C329 por_dig_0.clknet_1_0__leaf_osc_ck por_dig_0.cnt_por\[8\] 0.412046f
C330 a_34444_32517# por_dig_0._026_ 0.383836f
C331 avdd porb_h 4.14283f
C332 a_39162_33453# dvdd 0.286534f
C333 a_25724_13935# avss 0.465525f
C334 por_dig_0.net22 a_34357_33427# 0.144025f
C335 por_dig_0.net24 a_32019_33819# 0.160628f
C336 a_39888_24823# a_39888_23693# 0.170258f
C337 a_31413_29619# dvdd 0.247657f
C338 por_dig_0._024_ por_dig_0.cnt_por\[7\] 0.217488f
C339 a_34024_33703# dvdd 0.229385f
C340 por_dig_0.net8 dvdd 0.946233f
C341 por_dig_0.cnt_por\[8\] a_33774_31821# 0.329141f
C342 a_37064_34003# a_38145_34375# 0.102355f
C343 a_2921_15512# avss 0.47306f
C344 a_17408_13935# a_18164_13935# 0.296258f
C345 a_29702_24619# a_30070_23637# 0.138963f
C346 por_dig_0.net4 por_dig_0._035_ 0.243863f
C347 a_21254_24619# dvdd 0.387414f
C348 por_dig_0._016_ por_dig_0.cnt_por\[2\] 0.284689f
C349 por_ana_0.rstring_mux_0.vtrip6 avss 2.27146f
C350 por_dig_0._035_ por_dig_0._037_ 0.564764f
C351 a_36406_21903# dvdd 0.176016f
C352 por_dig_0._014_ a_34378_30189# 0.214165f
C353 por_ana_0.rstring_mux_0.otrip_decoded_b_avdd[7] avss 0.36282f
C354 a_35776_36967# por_dig_0._049_ 0.101385f
C355 por_dig_0.net33 por_dig_0._041_ 0.147233f
C356 por_ana_0.rstring_mux_0.otrip_decoded_avdd[7] por_ana_0.rstring_mux_0.otrip_decoded_b_avdd[6] 0.155152f
C357 a_25595_33708# a_26802_33372# 0.28899f
C358 por_dig_0.net6 a_33155_28640# 0.141579f
C359 por_dig_0.otrip_decoded[0] avdd 0.949356f
C360 a_35174_6535# avss 0.466333f
C361 por_dig_0._007_ dvdd 0.796193f
C362 por_ana_0.rstring_mux_0.vtrip4 por_ana_0.rstring_mux_0.vtrip6 0.859994f
C363 a_31412_31251# dvdd 0.359746f
C364 a_29702_22885# a_29802_22973# 0.40546f
C365 a_34828_29253# por_dig_0.net15 0.142278f
C366 por_ana_0.rstring_mux_0.otrip_decoded_b_avdd[4] avdd 0.903548f
C367 avdd startup_timed_out 0.225449f
C368 a_34294_21903# avdd 0.143952f
C369 avdd osc_ck 1.16667f
C370 a_36862_30739# a_37212_31111# 0.22382f
C371 por_dig_0.net4 por_dig_0.cnt_st\[4\] 0.162271f
C372 por_dig_0.cnt_st\[4\] por_dig_0._042_ 0.509331f
C373 a_20432_13935# avss 0.465068f
C374 a_5567_22912# a_6323_22912# 0.296258f
C375 a_35092_33427# dvdd 0.350227f
C376 a_33121_22637# avdd 0.421965f
C377 por_dig_0.net24 a_33444_31037# 0.276678f
C378 por_dig_0.cnt_por\[7\] dvdd 0.710745f
C379 a_32616_32125# a_32441_32199# 0.233657f
C380 por_dig_0._000_ a_37230_34003# 0.737297f
C381 a_30495_21859# a_30070_21903# 0.460766f
C382 a_36016_35629# dvdd 0.194254f
C383 por_dig_0.net24 a_33821_36551# 0.250567f
C384 por_dig_0.net22 osc_ck 0.178269f
C385 por_dig_0._044_ a_39510_31251# 0.117375f
C386 por_dig_0.net1 a_31592_30965# 0.287535f
C387 por_dig_0._015_ a_35645_31277# 0.15859f
C388 por_ana_0.rstring_mux_0.vtrip_decoded_b_avdd[6] avss 0.363573f
C389 force_short_oneshot otrip[2] 0.239384f
C390 a_31893_33721# a_32019_33819# 0.186387f
C391 a_31932_33595# a_32088_33690# 0.107482f
C392 por_dig_0.net22 por_dig_0.cnt_rsb 0.252439f
C393 a_36480_31251# dvdd 0.364762f
C394 por_ana_0.rstring_mux_0.vtrip_decoded_b_avdd[3] avdd 0.903548f
C395 a_31360_33997# dvdd 0.278577f
C396 por_dig_0.net24 por_dig_0._010_ 0.485912f
C397 a_29882_6535# avss 0.466333f
C398 por_dig_0._051_ por_dig_0._008_ 0.119765f
C399 por_dig_0._033_ por_dig_0.clknet_0_osc_ck 0.209525f
C400 por_ana_0.comparator_0.vnn avss 3.71311f
C401 por_dig_0.net4 por_dig_0._032_ 0.141547f
C402 dvdd otrip[0] 0.541238f
C403 a_23734_23637# dvdd 0.16995f
C404 a_37820_13935# a_38576_13935# 0.296258f
C405 por_dig_0.cnt_por\[0\] a_35450_35124# 0.267756f
C406 por_dig_0._042_ por_dig_0._032_ 0.16328f
C407 a_36880_33453# a_37961_33453# 0.102325f
C408 a_35202_29877# a_35298_29619# 0.419086f
C409 a_17776_27844# a_18532_27844# 0.296258f
C410 por_ana_0.schmitt_trigger_0.in por_ana_0.rstring_mux_0.vtrip_decoded_avdd[2] 0.13771f
C411 por_dig_0._019_ a_35640_32517# 0.112309f
C412 a_31814_24619# dvdd 0.379209f
C413 por_dig_0.net24 por_dig_0._052_ 0.153858f
C414 a_15140_13935# avss 0.465264f
C415 por_dig_0.cnt_por\[5\] por_dig_0.cnt_por\[9\] 0.243535f
C416 a_37138_30189# a_37488_30189# 0.20669f
C417 a_40247_23627# avdd 0.260039f
C418 por_dig_0.cnt_por\[7\] a_34010_31821# 0.101703f
C419 a_36038_22885# a_36406_21903# 0.138963f
C420 a_37430_30707# dvdd 0.208259f
C421 a_36138_24707# a_37345_24371# 0.28899f
C422 por_ana_0.comparator_0.vnn vbg_1v2 0.779817f
C423 por_dig_0._002_ a_37046_32915# 0.74233f
C424 a_29802_24707# avdd 0.863296f
C425 a_32607_21859# dvdd 0.104499f
C426 por_dig_0.net1 por_dig_0.clknet_1_0__leaf_osc_ck 0.548548f
C427 a_38957_32883# dvdd 0.218769f
C428 a_33971_28557# dvdd 0.259587f
C429 a_35500_35629# por_dig_0._005_ 0.160548f
C430 por_dig_0.osc_ena por_dig_0.otrip_decoded[1] 0.115347f
C431 por_dig_0._024_ dvdd 0.515031f
C432 por_dig_0.net7 dvdd 1.97733f
C433 por_dig_0.cnt_por\[1\] por_dig_0._046_ 0.132047f
C434 por_dig_0._001_ a_37301_33453# 0.161376f
C435 a_23078_6535# avss 0.466333f
C436 a_22047_23593# dvdd 0.104499f
C437 a_37706_30431# dvdd 0.204954f
C438 por_ana_0.rstring_mux_0.otrip_decoded_b_avdd[1] vin 0.342078f
C439 por_dig_0._019_ por_dig_0._026_ 0.237245f
C440 por_dig_0.net2 dvdd 0.201708f
C441 por_dig_0._034_ dvdd 2.10474f
C442 por_dig_0.otrip_decoded[5] dvdd 0.634734f
C443 por_ana_0.rstring_mux_0.vtrip4 avss 2.05606f
C444 a_31894_32365# dvdd 0.332984f
C445 por_dig_0._038_ dvdd 0.43689f
C446 por_dig_0._048_ por_dig_0.net4 0.196943f
C447 a_37504_32909# dvdd 0.142116f
C448 a_32630_32915# a_33545_33287# 0.125324f
C449 a_24673_22637# por_ana_0.rstring_mux_0.otrip_decoded_avdd[2] 0.135981f
C450 avss vbg_1v2 16.6753f
C451 a_32980_33287# dvdd 0.206801f
C452 por_dig_0._033_ por_dig_0.net23 1.06931f
C453 por_ana_0.schmitt_trigger_0.in por_dig_0.otrip_decoded[0] 0.368797f
C454 a_25478_22885# dvdd 0.380879f
C455 por_ana_0.rc_osc_0.ena_b por_ana_0.rc_osc_0.in 0.131788f
C456 por_dig_0.cnt_por\[4\] a_34387_32909# 0.278039f
C457 a_37046_33453# dvdd 0.574357f
C458 por_dig_0._052_ por_dig_0._051_ 0.100082f
C459 a_32188_30739# a_33269_31111# 0.102355f
C460 a_32922_30707# a_32704_31111# 0.209641f
C461 a_20054_6535# a_20810_6535# 0.296258f
C462 por_dig_0.otrip_decoded[1] por_dig_0.otrip_decoded[0] 0.8263f
C463 por_dig_0.clknet_1_0__leaf_osc_ck por_dig_0._036_ 0.815716f
C464 por_ana_0.comparator_0.vnn por_ana_0.comparator_0.vm 0.573444f
C465 a_36218_30163# dvdd 0.298248f
C466 a_17786_6535# avss 0.466333f
C467 a_23466_22973# avdd 0.863791f
C468 a_39887_23089# a_40246_23089# 0.249533f
C469 a_32528_13935# a_33284_13935# 0.296258f
C470 a_20054_6535# avdd 0.366615f
C471 por_dig_0.net15 por_dig_0.otrip_decoded[4] 0.100413f
C472 a_33806_33427# por_dig_0._010_ 0.11973f
C473 a_33996_35389# a_33821_35463# 0.233657f
C474 a_32740_36179# a_32906_36179# 0.887568f
C475 a_35100_32339# dvdd 0.356701f
C476 a_33012_33997# dvdd 0.286843f
C477 por_dig_0.cnt_por\[0\] por_dig_0.cnt_por\[2\] 1.01246f
C478 por_dig_0.net21 a_39732_31829# 0.182285f
C479 a_25495_33620# a_25863_32638# 0.138963f
C480 a_21178_35244# avss 0.721623f
C481 por_ana_0.dcomp3v3uv dvdd 1.08827f
C482 por_dig_0.net25 a_37961_33453# 0.267389f
C483 avss ibg_200n 3.46509f
C484 por_dig_0.cnt_por\[3\] por_dig_0._034_ 0.102983f
C485 por_dig_0.net5 por_dig_0.net7 2.0011f
C486 a_8213_15512# a_8969_15512# 0.296258f
C487 a_39718_33605# dvdd 0.179535f
C488 por_dig_0._015_ por_dig_0.net29 0.322f
C489 a_34719_21859# avdd 0.607928f
C490 por_dig_0.net30 dvdd 0.604801f
C491 por_dig_0.otrip_decoded[2] por_dig_0.otrip_decoded[4] 1.8816f
C492 a_34010_31821# dvdd 0.288809f
C493 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[3] dvdd 0.527183f
C494 a_31413_32339# por_dig_0.net19 0.181279f
C495 por_dig_0._028_ por_dig_0.net29 0.315624f
C496 por_dig_0.net4 por_dig_0.cnt_por\[4\] 0.364389f
C497 a_36831_21859# a_36406_21903# 0.460766f
C498 por_dig_0._000_ por_dig_0._039_ 0.146132f
C499 por_ana_0.rstring_mux_0.otrip_decoded_avdd[5] avss 1.34873f
C500 por_dig_0.net21 por_dig_0._030_ 0.219878f
C501 por_dig_0.clknet_1_0__leaf_osc_ck por_dig_0.net27 0.307641f
C502 a_31360_31827# a_31876_32199# 0.112384f
C503 por_ana_0.comparator_0.vm avss 10.399099f
C504 por_dig_0.cnt_por\[3\] dvdd 0.380362f
C505 a_29702_22885# a_30070_21903# 0.138963f
C506 por_ana_0.sky130_fd_sc_hvl__lsbufhv2lv_1_1.X dvdd 0.984529f
C507 por_dig_0.net6 a_36649_28789# 0.154668f
C508 a_39732_31829# startup_timed_out 0.156179f
C509 por_dig_0.cnt_st\[0\] a_38320_34301# 0.103164f
C510 por_dig_0._026_ por_dig_0.cnt_por\[10\] 0.112889f
C511 a_21254_24619# avdd 0.197715f
C512 por_dig_0.net6 a_34290_28557# 0.36041f
C513 a_25578_22973# a_26271_21859# 0.264594f
C514 por_dig_0._033_ por_dig_0.net22 0.163871f
C515 a_34580_34110# dvdd 0.202433f
C516 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[0] dvdd 0.275187f
C517 por_dig_0.net7 por_dig_0.otrip_decoded[6] 0.117452f
C518 por_dig_0.net24 por_dig_0._001_ 0.739404f
C519 a_15886_35244# avss 0.460203f
C520 a_31893_31545# dvdd 0.579842f
C521 a_29802_22973# a_31009_22637# 0.28899f
C522 por_dig_0.cnt_rsb a_34510_31277# 0.298482f
C523 a_41694_3516# a_41694_2760# 0.296258f
C524 por_ana_0.rc_osc_0.in a_19094_1626# 0.516433f
C525 a_36038_22885# dvdd 0.381067f
C526 a_36406_21903# avdd 0.143952f
C527 por_ana_0.rstring_mux_0.otrip_decoded_avdd[2] avss 1.41238f
C528 por_ana_0.sky130_fd_sc_hd__inv_4_1.Y dvdd 1.26215f
C529 por_dig_0.net5 dvdd 2.26522f
C530 a_36862_30739# a_37777_31111# 0.125324f
C531 por_ana_0.rstring_mux_0.otrip_decoded_b_avdd[0] por_ana_0.rstring_mux_0.vtrip0 0.191117f
C532 por_dig_0.clknet_0_osc_ck dvdd 2.16604f
C533 a_31360_33997# force_dis_rc_osc 0.197258f
C534 osc_ck porb 0.282824f
C535 a_34026_22973# avdd 0.863791f
C536 a_35573_33721# dvdd 0.570712f
C537 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[2] por_ana_0.rstring_mux_0.vtrip_decoded_b_avdd[1] 0.155018f
C538 por_ana_0.dcomp3v3uv por_ana_0.sky130_fd_sc_hvl__lsbufhv2lv_1_1.X 2.56892f
C539 por_dig_0.cnt_por\[10\] por_dig_0.cnt_por\[9\] 0.216388f
C540 por_dig_0.otrip_decoded[6] por_dig_0.otrip_decoded[5] 3.92951f
C541 por_ana_0.rstring_mux_0.vtrip0 a_25724_13935# 0.411488f
C542 por_dig_0._000_ por_dig_0.net25 0.141773f
C543 por_dig_0._030_ startup_timed_out 0.439212f
C544 por_dig_0.cnt_por\[9\] por_dig_0.net29 0.330999f
C545 a_36581_35629# dvdd 0.286993f
C546 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[0] por_ana_0.dcomp3v3uv 0.497383f
C547 a_14762_6535# a_15518_6535# 0.296258f
C548 por_dig_0.net24 a_37396_33287# 0.163622f
C549 por_ana_0.rstring_mux_0.vtrip2 avss 2.19733f
C550 por_dig_0.cnt_st\[1\] dvdd 1.20055f
C551 a_32088_33690# a_32019_33819# 0.209641f
C552 por_dig_0.clknet_1_0__leaf_osc_ck a_31932_31419# 0.289403f
C553 a_37392_31251# dvdd 0.168663f
C554 por_ana_0.rstring_mux_0.vtrip2 por_ana_0.rstring_mux_0.vtrip4 0.994518f
C555 a_36381_36691# dvdd 0.254977f
C556 por_dig_0.otrip_decoded[6] dvdd 0.909606f
C557 por_ana_0.rstring_mux_0.otrip_decoded_avdd[7] vin 0.875535f
C558 por_dig_0._001_ por_dig_0._002_ 0.149025f
C559 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[1] por_ana_0.rstring_mux_0.vtrip_decoded_avdd[2] 0.618116f
C560 por_dig_0.otrip_decoded[0] otrip[2] 0.144826f
C561 por_dig_0.net8 a_32088_31514# 0.162429f
C562 a_31413_29075# por_dig_0.force_pdnb 0.168257f
C563 a_27958_23637# dvdd 0.169343f
C564 por_dig_0.net22 por_dig_0.cnt_por\[7\] 0.580397f
C565 por_dig_0._001_ por_dig_0.cnt_st\[2\] 0.12168f
C566 a_35298_29619# a_35556_29619# 0.22264f
C567 a_36328_35091# dvdd 0.442403f
C568 a_6323_22912# avss 0.474704f
C569 a_18154_35244# a_18910_35244# 0.296258f
C570 a_38150_24619# a_38518_23637# 0.138963f
C571 a_37230_34003# a_37580_34375# 0.219633f
C572 por_dig_0.net23 por_dig_0._034_ 0.685534f
C573 avdd otrip[0] 0.225281f
C574 a_2921_15512# a_3677_15512# 0.296258f
C575 a_37138_30189# a_38053_30189# 0.118759f
C576 a_23734_23637# avdd 0.143132f
C577 a_32794_33971# por_dig_0._012_ 0.12144f
C578 por_ana_0.rstring_mux_0.otrip_decoded_avdd[4] vin 0.879587f
C579 a_37952_31037# dvdd 0.347365f
C580 por_dig_0.net31 por_dig_0._039_ 0.137737f
C581 por_dig_0.net24 a_32464_32915# 0.957784f
C582 a_31615_31529# a_31932_31419# 0.102355f
C583 por_dig_0.cnt_st\[1\] a_39718_33605# 0.168023f
C584 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[3] por_ana_0.rstring_mux_0.vtrip_decoded_b_avdd[2] 0.155157f
C585 a_38576_13935# avss 0.82426f
C586 a_31814_24619# avdd 0.206171f
C587 por_dig_0.por_unbuf a_25495_33620# 0.259533f
C588 por_ana_0.comparator_0.vn por_ana_0.comparator_0.n0 1.99139f
C589 por_dig_0._040_ a_38957_32883# 0.184745f
C590 a_18532_27844# avss 0.460203f
C591 osc_ck por_timed_out 0.681172f
C592 a_34467_28557# dvdd 0.21398f
C593 por_dig_0._033_ por_dig_0.cnt_por\[1\] 0.206467f
C594 por_dig_0.net4 por_dig_0.net33 0.349479f
C595 por_ana_0.rstring_mux_0.otrip_decoded_b_avdd[6] por_ana_0.rstring_mux_0.vtrip6 0.190544f
C596 por_dig_0.net23 dvdd 2.01786f
C597 por_ana_0.sky130_fd_sc_hd__inv_4_1.A dvdd 0.677586f
C598 por_dig_0.net24 por_dig_0.cnt_por\[4\] 0.37439f
C599 por_ana_0.rstring_mux_0.otrip_decoded_avdd[3] por_ana_0.rstring_mux_0.otrip_decoded_avdd[4] 0.503487f
C600 a_32607_21859# avdd 0.607928f
C601 a_31894_32365# a_32244_32365# 0.216626f
C602 por_dig_0._012_ a_31728_32365# 0.131264f
C603 dvdd force_dis_rc_osc 0.760658f
C604 por_ana_0.sky130_fd_sc_hvl__inv_1_0.A por_dig_0.por_unbuf 0.166464f
C605 a_39888_24823# a_40247_24823# 0.249533f
C606 a_38228_30163# dvdd 0.389258f
C607 a_35174_6535# a_35930_6535# 0.296258f
C608 por_dig_0._047_ a_33600_34335# 0.155298f
C609 por_dig_0._007_ a_33161_36539# 0.161235f
C610 por_dig_0._035_ por_dig_0._028_ 0.151355f
C611 a_33121_24371# por_ana_0.rstring_mux_0.vtrip_decoded_avdd[3] 0.13699f
C612 por_dig_0.force_pdnb por_dig_0.otrip_decoded[3] 0.147422f
C613 a_38352_32365# dvdd 0.224566f
C614 a_35295_33705# a_35612_33595# 0.102325f
C615 por_dig_0.net4 a_36862_30739# 0.294222f
C616 por_dig_0.net25 a_35224_31277# 0.295232f
C617 a_37156_28013# dvdd 0.297346f
C618 a_22047_23593# avdd 0.607831f
C619 a_32244_32365# dvdd 0.194599f
C620 por_dig_0._024_ por_dig_0.net22 0.908888f
C621 por_ana_0.comparator_0.vn avdd 0.753795f
C622 a_36831_21859# dvdd 0.104499f
C623 a_27590_24619# a_27690_24707# 0.40546f
C624 a_39510_31251# dvdd 0.210633f
C625 a_33284_13935# avss 0.484363f
C626 por_dig_0.otrip_decoded[5] avdd 0.217399f
C627 por_dig_0.net5 por_dig_0.otrip_decoded[6] 0.502126f
C628 a_33545_33287# dvdd 0.297689f
C629 por_dig_0._040_ dvdd 0.344134f
C630 por_dig_0._027_ a_33852_29645# 0.246866f
C631 por_dig_0.clknet_1_1__leaf_osc_ck a_35612_33595# 0.272577f
C632 por_ana_0.dcomp3v3uv por_ana_0.comparator_0.n0 0.388405f
C633 a_38936_32159# dvdd 0.225539f
C634 por_dig_0.cnt_por\[8\] a_33804_31251# 0.12199f
C635 a_37396_33453# dvdd 0.1998f
C636 a_20432_13935# a_21188_13935# 0.296258f
C637 a_8969_15512# avss 0.769579f
C638 a_37046_33453# a_37396_33453# 0.229804f
C639 por_dig_0._048_ por_dig_0._006_ 0.488085f
C640 por_dig_0.otrip_decoded[1] a_21254_24619# 0.249645f
C641 por_ana_0.rstring_mux_0.otrip_decoded_avdd[2] por_ana_0.rstring_mux_0.vtrip2 0.478934f
C642 a_25478_22885# avdd 0.207177f
C643 avdd dvdd 65.8375f
C644 a_33996_36477# a_33821_36551# 0.233657f
C645 por_dig_0.otrip_decoded[4] por_ana_0.rstring_mux_0.otrip_decoded_avdd[2] 0.100242f
C646 por_dig_0._013_ dvdd 0.78665f
C647 por_dig_0.cnt_por\[6\] osc_ck 0.136253f
C648 por_dig_0.net12 a_33172_28165# 0.14168f
C649 a_32740_36179# por_dig_0.net24 0.299864f
C650 por_ana_0.rstring_mux_0.vtrip0 avss 2.36542f
C651 por_dig_0._035_ por_dig_0.cnt_por\[9\] 0.178154f
C652 por_dig_0._016_ por_dig_0.clknet_1_1__leaf_osc_ck 0.598055f
C653 por_dig_0.net6 a_35674_28557# 0.10559f
C654 por_dig_0.net22 dvdd 2.81967f
C655 por_ana_0.rstring_mux_0.vtrip0 por_ana_0.rstring_mux_0.vtrip4 0.655814f
C656 por_ana_0.sky130_fd_sc_hd__inv_4_1.A por_ana_0.sky130_fd_sc_hd__inv_4_1.Y 0.392612f
C657 por_ana_0.rstring_mux_0.otrip_decoded_avdd[1] vin 0.881159f
C658 por_dig_0.net23 por_dig_0.clknet_0_osc_ck 0.621304f
C659 a_39718_33605# por_dig_0._040_ 0.111244f
C660 por_ana_0.sky130_fd_sc_hd__inv_4_0.Y dvdd 1.35239f
C661 por_dig_0._047_ por_dig_0._051_ 0.499693f
C662 por_ana_0.dcomp3v3uv avdd 5.83043f
C663 por_dig_0.cnt_st\[2\] a_38926_33453# 0.290424f
C664 a_40247_23627# a_39888_23693# 0.249269f
C665 por_dig_0.net24 a_36234_35871# 0.166131f
C666 a_35000_31795# dvdd 0.474379f
C667 a_31592_30965# a_31864_30823# 0.13675f
C668 por_dig_0.cnt_por\[8\] por_dig_0._037_ 0.625692f
C669 por_dig_0.net25 por_dig_0._003_ 0.228302f
C670 a_38943_21859# a_38518_21903# 0.460766f
C671 a_3677_15512# avss 0.472978f
C672 a_31814_24619# a_32182_23637# 0.138963f
C673 a_32094_31795# a_31876_32199# 0.209641f
C674 a_31360_31827# a_32441_32199# 0.102355f
C675 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[3] avdd 1.87754f
C676 a_34357_33427# por_dig_0.cnt_por\[5\] 0.122056f
C677 por_dig_0.osc_ena por_ana_0.rc_osc_0.ena_b 0.528234f
C678 por_dig_0._021_ a_34357_33427# 0.101999f
C679 a_29882_6535# a_30638_6535# 0.296258f
C680 por_dig_0.cnt_st\[0\] por_dig_0._039_ 0.25367f
C681 por_dig_0._015_ a_35390_31277# 0.208266f
C682 a_32701_28531# por_dig_0.net12 0.179511f
C683 a_32039_28013# otrip[0] 0.266434f
C684 por_ana_0.rstring_mux_0.otrip_decoded_b_avdd[6] avss 0.36281f
C685 a_36380_33971# dvdd 0.322543f
C686 a_22561_24371# avdd 0.421008f
C687 a_35930_6535# avss 0.466333f
C688 por_dig_0.otrip_decoded[1] otrip[0] 0.575585f
C689 por_dig_0._047_ a_33806_33427# 0.168045f
C690 a_32088_31514# dvdd 0.199628f
C691 a_22561_22637# por_ana_0.rstring_mux_0.otrip_decoded_avdd[0] 0.135767f
C692 por_dig_0.net4 por_dig_0.clknet_1_0__leaf_osc_ck 0.294337f
C693 a_19094_3138# a_19094_2382# 0.296258f
C694 por_ana_0.rstring_mux_0.otrip_decoded_b_avdd[3] avdd 0.903548f
C695 por_ana_0.sky130_fd_sc_hvl__lsbufhv2lv_1_1.X avdd 2.97006f
C696 a_35583_34541# dvdd 1.31595f
C697 a_20800_27844# por_ana_0.schmitt_trigger_0.in 0.303942f
C698 por_dig_0.clknet_1_1__leaf_osc_ck a_32740_35091# 0.271843f
C699 por_dig_0.cnt_st\[1\] a_38352_32365# 0.27322f
C700 por_ana_0.rstring_mux_0.vtop avss 3.611f
C701 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[0] avdd 1.59456f
C702 a_21188_13935# avss 0.465068f
C703 a_35768_33690# dvdd 0.205442f
C704 a_36038_22885# avdd 0.207177f
C705 por_dig_0.clknet_1_0__leaf_osc_ck a_34212_30189# 0.455132f
C706 a_33774_31821# por_dig_0._037_ 0.109537f
C707 a_38320_34301# a_38145_34375# 0.233657f
C708 por_dig_0.cnt_por\[1\] por_dig_0._034_ 0.153524f
C709 a_36124_35995# dvdd 0.140723f
C710 por_dig_0.clknet_1_1__leaf_osc_ck por_dig_0._012_ 0.21602f
C711 por_dig_0.net20 por_dig_0._035_ 0.135015f
C712 por_ana_0.schmitt_trigger_0.m dvdd 2.68035f
C713 a_15140_13935# a_15896_13935# 0.296258f
C714 por_dig_0.net24 a_37961_33287# 0.213015f
C715 por_dig_0.cnt_st\[1\] por_dig_0._040_ 0.262179f
C716 por_dig_0.cnt_st\[0\] por_dig_0.net21 0.113294f
C717 por_ana_0.rstring_mux_0.vtrip_decoded_b_avdd[5] avss 0.363125f
C718 por_dig_0.cnt_st\[0\] por_dig_0.net25 0.605126f
C719 force_pdn pwup_filt 0.754834f
C720 a_35774_28673# dvdd 0.192842f
C721 por_dig_0.cnt_rsb_stg1 a_31566_32909# 0.291561f
C722 por_ana_0.rstring_mux_0.vtrip_decoded_b_avdd[2] avdd 0.903548f
C723 a_31360_28557# dvdd 0.263686f
C724 por_dig_0.cnt_por\[1\] dvdd 1.80403f
C725 por_dig_0.cnt_por\[5\] osc_ck 0.30336f
C726 a_30638_6535# avss 0.466333f
C727 a_37789_31821# por_dig_0._045_ 0.109093f
C728 a_35040_34587# por_dig_0.net4 0.138234f
C729 a_31413_29075# por_dig_0.net9 0.176857f
C730 a_21254_22885# a_21354_22973# 0.40546f
C731 por_dig_0._026_ por_dig_0.net32 0.480494f
C732 por_dig_0._041_ a_39634_32615# 0.131344f
C733 a_32182_23637# dvdd 0.169343f
C734 por_dig_0.otrip_decoded[6] avdd 0.493379f
C735 a_37062_35059# dvdd 0.211024f
C736 a_19666_35244# osc_ck 0.256787f
C737 por_dig_0.net24 a_31728_32365# 0.299648f
C738 a_34026_24707# dvdd 0.238523f
C739 por_dig_0.net25 a_37580_34375# 0.157564f
C740 a_37230_34003# a_38145_34375# 0.124988f
C741 force_ena_rc_osc force_pdn 2.51978f
C742 por_dig_0._044_ por_dig_0._003_ 0.205607f
C743 a_15896_13935# avss 0.466481f
C744 a_38957_32883# a_39094_32909# 0.126609f
C745 a_3299_22912# a_4055_22912# 0.296258f
C746 a_27958_23637# avdd 0.142934f
C747 por_ana_0.comparator_1.vn avss 8.65812f
C748 a_38150_22885# a_38518_21903# 0.138963f
C749 a_38146_31429# a_38242_31251# 0.419086f
C750 a_39497_30849# dvdd 0.173548f
C751 a_38150_24619# a_38250_24707# 0.40546f
C752 por_ana_0.schmitt_trigger_0.in dvdd 2.47753f
C753 por_ana_0.dcomp3v3 por_ana_0.vl 10.0456f
C754 por_dig_0.net24 a_33198_32883# 0.207877f
C755 a_34378_30189# a_34946_30431# 0.182409f
C756 a_31893_31545# a_32088_31514# 0.229804f
C757 a_32039_28013# dvdd 0.227179f
C758 a_33121_24371# avdd 0.420074f
C759 a_33474_36147# dvdd 0.209597f
C760 por_dig_0.cnt_por\[4\] a_35640_32517# 0.170468f
C761 por_dig_0.otrip_decoded[1] dvdd 1.23602f
C762 por_ana_0.rstring_mux_0.vtrip0 por_ana_0.rstring_mux_0.vtrip2 0.847499f
C763 a_23078_6535# a_23834_6535# 0.296258f
C764 por_ana_0.comparator_1.vn vbg_1v2 0.204188f
C765 por_dig_0.clknet_0_osc_ck a_35583_34541# 0.357331f
C766 a_23834_6535# avss 0.466333f
C767 a_31894_32365# a_32809_32365# 0.125324f
C768 por_ana_0.schmitt_trigger_0.in por_ana_0.dcomp3v3uv 0.122613f
C769 por_dig_0._036_ a_33804_31251# 0.109303f
C770 a_35552_13935# a_36308_13935# 0.296258f
C771 a_32906_35091# dvdd 0.573815f
C772 por_dig_0.cnt_por\[0\] a_36756_35603# 0.458658f
C773 por_ana_0.rstring_mux_0.otrip_decoded_b_avdd[0] vin 0.343304f
C774 a_37230_34003# a_37798_33971# 0.175891f
C775 por_dig_0.cnt_por\[1\] por_dig_0.cnt_por\[3\] 0.327055f
C776 a_15508_27844# a_16264_27844# 0.296258f
C777 por_dig_0.cnt_st\[3\] dvdd 0.79651f
C778 a_35573_33721# a_35768_33690# 0.219633f
C779 por_dig_0.net7 a_34934_28013# 0.384846f
C780 por_dig_0.clknet_1_1__leaf_osc_ck a_37064_34003# 0.26365f
C781 avdd force_dis_rc_osc 0.215136f
C782 por_dig_0.osc_ena por_dig_0.otrip_decoded[3] 0.108398f
C783 a_32809_32365# dvdd 0.29816f
C784 por_dig_0._035_ a_36382_31795# 0.162225f
C785 a_39094_32909# dvdd 0.197837f
C786 por_dig_0.net24 por_dig_0.clknet_1_0__leaf_osc_ck 0.379148f
C787 por_dig_0.net5 a_35774_28673# 0.282979f
C788 a_27690_24707# a_28897_24371# 0.28899f
C789 por_ana_0.schmitt_trigger_0.in por_ana_0.rstring_mux_0.vtrip_decoded_avdd[3] 0.14576f
C790 a_40246_21893# dvdd 0.47489f
C791 por_dig_0.cnt_por\[0\] por_dig_0.clknet_1_1__leaf_osc_ck 0.531057f
C792 por_ana_0.comparator_0.n0 avdd 1.07016f
C793 por_dig_0.net23 por_dig_0.net22 0.291169f
C794 por_dig_0._033_ por_dig_0.cnt_por\[6\] 0.128143f
C795 a_36880_32915# dvdd 0.416389f
C796 por_dig_0._003_ a_36972_30189# 0.617494f
C797 a_34510_31277# dvdd 0.262824f
C798 por_ana_0.rc_osc_0.in por_ana_0.rc_osc_0.vr 0.494137f
C799 por_dig_0.otrip_decoded[4] por_dig_0.otrip_decoded[7] 0.106636f
C800 a_39732_31829# dvdd 0.250626f
C801 a_36831_21859# avdd 0.607928f
C802 a_37961_33453# dvdd 0.288491f
C803 a_33444_31037# a_33269_31111# 0.233657f
C804 por_ana_0.rstring_mux_0.vtrip6 vin 2.08469f
C805 por_dig_0.cnt_por\[0\] a_35704_35124# 0.318482f
C806 a_37046_33453# a_37961_33453# 0.125324f
C807 a_36382_31795# por_dig_0.cnt_st\[4\] 0.13586f
C808 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A avdd 3.72269f
C809 por_ana_0.rstring_mux_0.otrip_decoded_b_avdd[7] vin 0.340862f
C810 a_38150_24619# isrc_sel 0.221894f
C811 a_18542_6535# avss 0.466333f
C812 por_dig_0.net4 por_dig_0._036_ 0.508389f
C813 por_ana_0.schmitt_trigger_0.in por_ana_0.rstring_mux_0.vtrip_decoded_avdd[0] 0.128751f
C814 a_26785_22637# avdd 0.421965f
C815 por_dig_0.net28 por_dig_0.net19 0.156259f
C816 a_31615_33705# dvdd 0.299247f
C817 a_37320_30733# dvdd 0.142144f
C818 por_dig_0.cnt_por\[9\] a_35468_30163# 0.114998f
C819 a_34212_33997# dvdd 0.206798f
C820 dvdd porb 2.334f
C821 a_34934_28013# dvdd 0.181122f
C822 por_dig_0._009_ a_36331_33819# 0.170255f
C823 dvdd por 2.0627f
C824 por_dig_0.net20 por_dig_0._048_ 0.865776f
C825 a_37046_32915# a_37614_32883# 0.175891f
C826 por_dig_0.net5 a_32039_28013# 0.159634f
C827 por_dig_0.net23 a_36380_33971# 0.239329f
C828 por_dig_0.net20 por_dig_0.cnt_por\[2\] 0.396402f
C829 por_dig_0._045_ por_dig_0.net34 0.256804f
C830 por_dig_0._030_ dvdd 0.69984f
C831 a_30495_21859# dvdd 0.104499f
C832 por_dig_0.net20 por_dig_0.por_unbuf 0.224859f
C833 por_dig_0._005_ a_35666_35629# 0.206326f
C834 por_dig_0.net25 por_dig_0.cnt_por\[10\] 0.728218f
C835 a_21354_22973# a_22047_21859# 0.264594f
C836 por_dig_0.otrip_decoded[5] a_25478_24619# 0.257733f
C837 por_dig_0.otrip_decoded[3] por_dig_0.otrip_decoded[0] 6.40722f
C838 por_dig_0.net23 a_35583_34541# 0.1487f
C839 por_dig_0.net24 a_35295_33705# 0.247073f
C840 a_37504_33819# dvdd 0.142182f
C841 por_dig_0.otrip_decoded[5] otrip[2] 0.187329f
C842 por_ana_0.sky130_fd_sc_hd__inv_4_3.Y dvdd 1.31104f
C843 por_dig_0.cnt_por\[6\] por_dig_0.cnt_por\[7\] 0.77587f
C844 por_dig_0.cnt_por\[1\] a_36328_35091# 0.609356f
C845 por_dig_0.net24 a_36756_35603# 0.300141f
C846 por_dig_0._042_ a_37789_31821# 0.129217f
C847 a_26271_23593# a_25846_23637# 0.460766f
C848 a_40246_21893# por_ana_0.sky130_fd_sc_hvl__lsbufhv2lv_1_1.X 0.142786f
C849 a_17786_6535# a_18542_6535# 0.296258f
C850 a_36376_28789# a_36649_28789# 0.167615f
C851 por_dig_0._014_ dvdd 0.370755f
C852 a_25478_24619# dvdd 0.38629f
C853 por_dig_0.por_unbuf dcomp 0.47137f
C854 por_dig_0.net8 a_32616_32125# 0.278389f
C855 a_13250_6535# avss 0.732759f
C856 por_dig_0._033_ por_dig_0._011_ 0.661249f
C857 dvdd otrip[2] 0.4752f
C858 por_dig_0.clknet_1_1__leaf_osc_ck por_dig_0.net24 0.524323f
C859 a_31814_22885# a_32182_21903# 0.138963f
C860 a_13894_21948# ibg_200n 0.401026f
C861 a_30260_13935# a_31016_13935# 0.296258f
C862 a_32188_30739# dvdd 0.479501f
C863 por_ana_0.sky130_fd_sc_hvl__inv_4_0.A por_ana_0.sky130_fd_sc_hvl__inv_16_0.A 0.751125f
C864 por_dig_0._000_ dvdd 0.538962f
C865 a_23466_24707# avdd 0.865353f
C866 por_dig_0.net23 por_dig_0.cnt_por\[1\] 0.774112f
C867 a_16642_35244# avss 0.460203f
C868 a_31814_22885# a_31914_22973# 0.40546f
C869 por_ana_0.rc_osc_0.in a_19094_870# 0.770709f
C870 por_ana_0.comparator_1.ena_b avss 1.77799f
C871 a_39070_34515# dvdd 0.283778f
C872 dvdd por_timed_out 0.5288f
C873 por_dig_0.cnt_por\[10\] por_dig_0.cnt_rsb 0.14288f
C874 a_5945_15512# a_6701_15512# 0.296258f
C875 por_ana_0.sky130_fd_sc_hvl__inv_4_0.A avdd 1.01598f
C876 a_37345_22637# avdd 0.421965f
C877 por_dig_0._033_ por_dig_0.cnt_por\[5\] 0.244697f
C878 por_dig_0._014_ por_dig_0.net30 0.131778f
C879 por_dig_0._021_ a_34024_33703# 0.129f
C880 por_ana_0.sky130_fd_sc_hvl__inv_1_0.A avss 2.17417f
C881 por_dig_0.net22 a_36380_33971# 0.166963f
C882 por_ana_0.sky130_fd_sc_hd__inv_4_1.Y porb 1.49255f
C883 a_35233_22637# por_ana_0.rstring_mux_0.vtrip_decoded_avdd[4] 0.135915f
C884 por_dig_0.net7 por_dig_0.net13 0.171866f
C885 por_ana_0.ibias_gen_0.vp1 por_ana_0.dcomp3v3uv 0.195418f
C886 a_33088_32909# dvdd 0.143138f
C887 avss vin 14.4483f
C888 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[4] avss 1.50015f
C889 por_dig_0.cnt_por\[2\] a_34672_35451# 0.125416f
C890 por_ana_0.sky130_fd_sc_hd__inv_4_4.Y dvdd 1.32154f
C891 a_21354_22973# a_22561_22637# 0.28899f
C892 a_38198_6535# a_38954_6535# 0.296258f
C893 a_34496_29645# dvdd 0.16772f
C894 por_ana_0.rstring_mux_0.vtrip4 vin 2.26482f
C895 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[4] por_ana_0.rstring_mux_0.vtrip4 0.497379f
C896 por_dig_0.clknet_1_1__leaf_osc_ck a_31893_33721# 0.173269f
C897 por_dig_0.osc_ena a_19676_13935# 0.318308f
C898 a_37584_35389# dvdd 0.431447f
C899 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[1] dvdd 0.335417f
C900 a_7079_22912# avss 0.471605f
C901 avss force_pdn 0.236529f
C902 por_dig_0.net24 a_32462_32607# 0.166268f
C903 a_36038_24619# dvdd 0.442417f
C904 por_dig_0.net25 a_38145_34375# 0.247703f
C905 por_ana_0.rstring_mux_0.otrip_decoded_avdd[3] avss 1.341f
C906 por_dig_0.cnt_st\[1\] por_dig_0._030_ 0.78139f
C907 vin vbg_1v2 7.770431f
C908 a_32182_23637# avdd 0.142934f
C909 por_ana_0.comparator_1.n0 avss 3.89953f
C910 a_38242_31251# a_38500_31251# 0.22264f
C911 a_38250_24707# a_39457_24371# 0.28899f
C912 a_28897_24371# por_ana_0.rstring_mux_0.otrip_decoded_avdd[7] 0.13699f
C913 por_dig_0._002_ por_dig_0._041_ 0.134256f
C914 por_dig_0.net24 a_33720_33213# 0.337518f
C915 a_34946_30431# a_34728_30189# 0.209641f
C916 a_32535_28013# dvdd 0.206669f
C917 a_34026_24707# avdd 0.863296f
C918 a_19288_27844# avss 0.460203f
C919 por_dig_0.net25 a_36328_29645# 0.176179f
C920 por_dig_0._023_ dvdd 0.302411f
C921 por_dig_0._035_ por_dig_0._031_ 0.106346f
C922 por_dig_0.cnt_por\[6\] dvdd 0.876002f
C923 por_dig_0.net13 dvdd 0.417179f
C924 por_dig_0._033_ por_dig_0._019_ 0.294628f
C925 por_ana_0.rstring_mux_0.otrip_decoded_avdd[6] dvdd 0.256793f
C926 a_35224_31277# dvdd 0.430335f
C927 por_dig_0._042_ por_dig_0.net34 0.789096f
C928 por_ana_0.schmitt_trigger_0.in avdd 4.55897f
C929 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[1] por_ana_0.dcomp3v3uv 0.100293f
C930 por_dig_0.net31 dvdd 0.293837f
C931 a_23456_13935# a_24212_13935# 0.296258f
C932 por_dig_0._042_ por_dig_0._045_ 0.180695f
C933 por_dig_0.net25 a_34946_30431# 0.166154f
C934 por_dig_0.cnt_por\[8\] por_dig_0._028_ 0.125236f
C935 por_dig_0.otrip_decoded[1] avdd 0.633872f
C936 a_40247_24823# a_40247_23627# 0.136815f
C937 a_36880_33453# por_dig_0._001_ 0.172728f
C938 a_33256_35463# dvdd 0.212294f
C939 a_37798_33971# por_dig_0.net25 0.171342f
C940 por_dig_0.otrip_decoded[6] otrip[2] 0.342618f
C941 por_dig_0._031_ por_dig_0.cnt_st\[4\] 0.612203f
C942 a_15886_35244# a_16642_35244# 0.296258f
C943 por_dig_0._033_ a_36100_32517# 0.224537f
C944 por_ana_0.rstring_mux_0.otrip_decoded_avdd[6] por_ana_0.dcomp3v3uv 0.148623f
C945 a_34444_32517# dvdd 0.331713f
C946 por_dig_0.force_pdnb pwup_filt 0.151132f
C947 a_23734_21903# dvdd 0.176016f
C948 a_35592_36286# dvdd 0.244617f
C949 por_dig_0.clknet_1_0__leaf_osc_ck por_dig_0._015_ 0.296199f
C950 a_19676_13935# osc_ck 0.184314f
C951 por_dig_0.net25 por_dig_0.cnt_st\[4\] 0.20778f
C952 por_dig_0.clknet_1_0__leaf_osc_ck por_dig_0._028_ 0.2058f
C953 a_34040_13935# avss 0.525451f
C954 a_35776_36967# dvdd 0.235805f
C955 a_34852_31277# dvdd 0.164259f
C956 por_ana_0.rstring_mux_0.otrip_decoded_avdd[5] vin 0.876971f
C957 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[1] por_ana_0.rstring_mux_0.vtrip_decoded_avdd[0] 1.27051f
C958 por_dig_0.net28 a_31360_31827# 0.468696f
C959 por_ana_0.rc_osc_0.m por_ana_0.rc_osc_0.vr 0.559422f
C960 a_29702_22885# dvdd 0.380879f
C961 por_ana_0.vl a_14752_27844# 0.30641f
C962 a_40246_21893# avdd 0.260659f
C963 por_dig_0._019_ por_dig_0.cnt_por\[7\] 0.520487f
C964 por_dig_0.force_pdnb force_ena_rc_osc 0.15782f
C965 por_dig_0._030_ a_38352_32365# 0.170424f
C966 a_32616_32125# dvdd 0.358725f
C967 a_27690_22973# avdd 0.863791f
C968 por_dig_0.cnt_por\[8\] por_dig_0.cnt_por\[9\] 0.592594f
C969 por_ana_0.vl por_dig_0.osc_ena 0.109357f
C970 por_dig_0._031_ por_dig_0._032_ 0.753976f
C971 a_31932_33595# dvdd 0.466367f
C972 a_34633_36147# por_dig_0.cnt_por\[2\] 0.156245f
C973 a_32906_6535# a_33662_6535# 0.296258f
C974 por_dig_0.net10 por_dig_0.osc_ena 0.138459f
C975 a_31360_31827# a_31526_31827# 0.723725f
C976 a_29802_24707# a_30495_23593# 0.264594f
C977 por_dig_0._030_ a_39510_31251# 0.176794f
C978 por_dig_0._011_ dvdd 0.518808f
C979 por_dig_0.cnt_por\[6\] a_34580_34110# 0.247626f
C980 a_35217_28013# dvdd 0.183789f
C981 por_ana_0.rstring_mux_0.otrip_decoded_avdd[2] vin 0.880848f
C982 a_37614_32883# a_37396_33287# 0.209641f
C983 por_dig_0._003_ dvdd 0.861569f
C984 por_ana_0.comparator_1.vnn avdd 37.0545f
C985 por_dig_0.net5 por_dig_0.net13 0.342073f
C986 por_dig_0.net19 por_dig_0.net8 0.644336f
C987 por_dig_0._042_ por_dig_0._043_ 0.113634f
C988 por_dig_0.net7 por_dig_0.net11 0.120941f
C989 a_38444_28013# por_dig_0.otrip_decoded[0] 0.187607f
C990 por_dig_0.net4 a_33804_31251# 0.135264f
C991 avdd porb 0.341364f
C992 avdd por 0.499894f
C993 por_dig_0.net24 a_35612_33595# 0.299639f
C994 por_ana_0.schmitt_trigger_0.in por_ana_0.schmitt_trigger_0.m 0.95597f
C995 por_dig_0._018_ por_dig_0.cnt_por\[4\] 0.377237f
C996 por_dig_0.net4 a_39417_31795# 0.184301f
C997 por_dig_0._039_ por_dig_0._029_ 0.174782f
C998 por_dig_0.clknet_1_0__leaf_osc_ck por_dig_0.cnt_por\[9\] 0.251464f
C999 por_ana_0.rstring_mux_0.otrip_decoded_avdd[3] por_ana_0.rstring_mux_0.otrip_decoded_avdd[2] 1.42613f
C1000 a_30495_21859# avdd 0.607928f
C1001 por_dig_0._048_ por_dig_0._009_ 0.192166f
C1002 a_34719_23593# dvdd 0.107699f
C1003 por_ana_0.rstring_mux_0.vtrip2 vin 2.09579f
C1004 por_dig_0.clknet_1_1__leaf_osc_ck a_35500_35629# 0.280946f
C1005 por_dig_0.cnt_por\[5\] dvdd 1.2248f
C1006 force_dis_rc_osc por_timed_out 0.813238f
C1007 a_18164_13935# a_18920_13935# 0.296258f
C1008 a_4433_15512# avss 0.472978f
C1009 por_dig_0._021_ dvdd 0.273944f
C1010 por_dig_0.net22 a_34212_33997# 0.166549f
C1011 a_33926_24619# a_34294_23637# 0.138963f
C1012 a_36494_35091# a_36844_35463# 0.206984f
C1013 a_26271_21859# a_25846_21903# 0.460766f
C1014 por_ana_0.rc_osc_0.ena_b dvdd 0.491102f
C1015 por_dig_0.osc_ena por_ana_0.rc_osc_0.vr 1.29552f
C1016 a_32922_30707# dvdd 0.207011f
C1017 por_dig_0.net7 por_dig_0.net14 0.267005f
C1018 por_dig_0._014_ a_34633_30189# 0.161376f
C1019 por_ana_0.comparator_1.vm avdd 0.382522f
C1020 por_dig_0._024_ por_dig_0._019_ 0.157183f
C1021 por_ana_0.vl por_dig_0.otrip_decoded[0] 0.100361f
C1022 dvdd itest 0.232549f
C1023 por_ana_0.rstring_mux_0.otrip_decoded_b_avdd[5] avss 0.36282f
C1024 a_25478_24619# avdd 0.206171f
C1025 a_36686_6535# avss 0.466333f
C1026 a_33256_36551# dvdd 0.211937f
C1027 a_31914_22973# a_33121_22637# 0.28899f
C1028 por_ana_0.rstring_mux_0.otrip_decoded_avdd[0] dvdd 0.197825f
C1029 avdd otrip[2] 0.214638f
C1030 por_dig_0.net11 dvdd 1.76286f
C1031 por_ana_0.vl osc_ck 0.102868f
C1032 a_32004_30189# pwup_filt 0.202985f
C1033 por_ana_0.rstring_mux_0.otrip_decoded_b_avdd[2] avdd 0.903648f
C1034 por_dig_0.net24 a_36494_35091# 0.362828f
C1035 por_dig_0.cnt_rsb_stg1 dvdd 0.715707f
C1036 por_dig_0._013_ a_32188_30739# 0.61726f
C1037 por_dig_0.net21 por_dig_0._029_ 0.123102f
C1038 por_dig_0.cnt_st\[0\] dvdd 1.88636f
C1039 por_dig_0.net4 por_dig_0._042_ 0.288872f
C1040 por_dig_0._010_ a_32630_32915# 0.220826f
C1041 por_dig_0.net4 por_dig_0._037_ 0.370452f
C1042 a_21944_13935# avss 0.465068f
C1043 a_38250_22973# avdd 0.864301f
C1044 a_6323_22912# a_7079_22912# 0.296258f
C1045 por_ana_0.schmitt_trigger_0.in por_dig_0.otrip_decoded[1] 1.76133f
C1046 por_ana_0.ibias_gen_0.vp1 avdd 6.58519f
C1047 por_ana_0.rstring_mux_0.otrip_decoded_avdd[4] por_ana_0.rstring_mux_0.otrip_decoded_b_avdd[4] 0.57199f
C1048 avdd por_timed_out 0.214746f
C1049 a_12598_23626# avdd 0.466408f
C1050 por_ana_0.rstring_mux_0.vtrip_decoded_b_avdd[4] avss 0.36282f
C1051 a_37580_34375# dvdd 0.218678f
C1052 por_dig_0.net14 dvdd 0.695375f
C1053 por_dig_0._019_ dvdd 1.99582f
C1054 por_ana_0.rstring_mux_0.vtrip_decoded_b_avdd[1] avdd 0.903548f
C1055 por_dig_0.cnt_por\[0\] por_dig_0.net4 0.109156f
C1056 por_ana_0.rstring_mux_0.vtrip_decoded_b_avdd[4] por_ana_0.rstring_mux_0.vtrip4 0.190544f
C1057 a_31394_6535# avss 0.466333f
C1058 por_dig_0.cnt_st\[3\] a_39497_30849# 0.178651f
C1059 por_dig_0.cnt_por\[10\] a_36480_31251# 0.132536f
C1060 por_dig_0.net24 a_32740_35091# 0.301193f
C1061 por_dig_0.cnt_st\[0\] a_39718_33605# 0.149125f
C1062 a_31413_29075# dvdd 0.27517f
C1063 a_38518_23637# dvdd 0.172455f
C1064 a_35298_29619# dvdd 0.284002f
C1065 por_dig_0.otrip_decoded[2] otrip[1] 0.213411f
C1066 por_ana_0.rc_osc_0.vr osc_ck 0.678284f
C1067 por_dig_0._000_ a_37485_34363# 0.170092f
C1068 a_18532_27844# a_19288_27844# 0.296258f
C1069 a_20422_35244# osc_ck 0.162386f
C1070 por_dig_0._036_ por_dig_0._028_ 0.165788f
C1071 por_dig_0.net24 a_32984_32339# 0.291345f
C1072 por_dig_0.clknet_0_osc_ck por_dig_0.cnt_por\[5\] 0.140812f
C1073 por_dig_0.cnt_por\[2\] osc_ck 0.421951f
C1074 por_dig_0.net24 por_dig_0._012_ 0.253286f
C1075 por_ana_0.vl a_40247_23627# 0.148644f
C1076 a_16652_13935# avss 0.466465f
C1077 por_ana_0.dcomp3v3 avss 3.77654f
C1078 por_dig_0._005_ dvdd 0.429254f
C1079 por_dig_0.por_unbuf osc_ck 0.141357f
C1080 a_35030_28557# a_35130_28673# 0.167615f
C1081 a_36100_32517# dvdd 0.188641f
C1082 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[1] avdd 1.96911f
C1083 por_dig_0.net24 a_34387_32909# 0.15352f
C1084 a_34357_33427# por_dig_0.cnt_por\[4\] 0.1212f
C1085 por_dig_0.net23 a_35592_36286# 0.247071f
C1086 por_dig_0.force_pdnb por_dig_0.otrip_decoded[2] 0.11543f
C1087 a_33172_28165# dvdd 0.216477f
C1088 a_36038_24619# avdd 0.206171f
C1089 a_35390_31277# a_35958_31519# 0.175891f
C1090 por_ana_0.rc_osc_0.in avss 7.08974f
C1091 por_ana_0.rstring_mux_0.otrip_decoded_avdd[5] por_ana_0.rstring_mux_0.otrip_decoded_b_avdd[5] 0.573322f
C1092 por_ana_0.rstring_mux_0.ena_b avdd 6.38097f
C1093 por_dig_0._026_ por_dig_0._036_ 0.151807f
C1094 por_dig_0.net5 por_dig_0.net11 0.259654f
C1095 por_dig_0.otrip_decoded[5] por_dig_0.otrip_decoded[3] 0.579215f
C1096 por_dig_0.net25 a_35468_30163# 0.330155f
C1097 por_dig_0._034_ por_dig_0.net19 0.112588f
C1098 a_32610_35603# por_dig_0._047_ 0.192552f
C1099 a_24590_6535# avss 0.466333f
C1100 por_dig_0.net24 a_31412_33427# 0.271956f
C1101 por_ana_0.rstring_mux_0.otrip_decoded_avdd[6] avdd 1.62839f
C1102 a_32607_23593# dvdd 0.104499f
C1103 por_ana_0.rstring_mux_0.vtrip0 vin 2.24047f
C1104 por_dig_0.clknet_1_0__leaf_osc_ck a_34378_30189# 0.177451f
C1105 a_33821_35463# dvdd 0.300386f
C1106 por_dig_0.net27 por_dig_0._015_ 0.15533f
C1107 por_dig_0.otrip_decoded[3] dvdd 0.808385f
C1108 por_dig_0._036_ por_dig_0.cnt_por\[9\] 0.184691f
C1109 por_dig_0.cnt_st\[2\] a_38956_32339# 0.139983f
C1110 por_dig_0._019_ a_34580_34110# 0.220646f
C1111 por_dig_0.net22 por_dig_0.cnt_por\[6\] 0.6809f
C1112 por_dig_0.cnt_st\[0\] por_dig_0.cnt_st\[1\] 1.35682f
C1113 por_dig_0.net19 dvdd 1.31161f
C1114 por_dig_0.osc_ena pwup_filt 1.35161f
C1115 a_27958_21903# dvdd 0.176016f
C1116 a_29702_24619# a_29802_24707# 0.40546f
C1117 avss otrip[1] 0.249361f
C1118 avss dcomp 1.20481f
C1119 por_dig_0.net24 por_dig_0.net4 0.34178f
C1120 por_dig_0.net20 por_dig_0.clknet_1_1__leaf_osc_ck 0.763147f
C1121 por_dig_0.net4 a_33600_34335# 0.103511f
C1122 por_dig_0._006_ a_36494_35091# 0.217977f
C1123 a_31566_32909# a_31802_32909# 0.22264f
C1124 a_32701_28531# dvdd 0.266715f
C1125 por_dig_0._137__26.LO dvdd 0.434971f
C1126 a_34444_32517# por_dig_0._013_ 0.150358f
C1127 por_dig_0.cnt_por\[4\] osc_ck 0.414673f
C1128 por_dig_0._038_ a_31651_30341# 0.212464f
C1129 a_23734_21903# avdd 0.145138f
C1130 a_20810_6535# a_21566_6535# 0.296258f
C1131 por_dig_0.cnt_por\[10\] dvdd 1.14051f
C1132 por_dig_0.net23 por_dig_0.cnt_por\[5\] 0.815431f
C1133 por_dig_0.osc_ena force_ena_rc_osc 0.54727f
C1134 a_25595_33708# avdd 0.862939f
C1135 por_dig_0.net29 dvdd 0.338162f
C1136 a_19298_6535# avss 0.466333f
C1137 por_ana_0.rstring_mux_0.otrip_decoded_b_avdd[6] vin 0.340862f
C1138 a_29702_22885# avdd 0.207177f
C1139 a_32019_33819# dvdd 0.204974f
C1140 a_31651_30341# dvdd 0.132989f
C1141 a_33284_13935# a_34040_13935# 0.296258f
C1142 por_dig_0._018_ por_dig_0._017_ 0.557375f
C1143 a_31360_31827# por_dig_0.net8 0.313648f
C1144 a_31526_31827# a_32094_31795# 0.179079f
C1145 por_dig_0._008_ dvdd 0.322562f
C1146 por_dig_0.net6 otrip[1] 0.16727f
C1147 a_35394_28013# dvdd 0.150874f
C1148 por_dig_0.net5 a_33172_28165# 0.132501f
C1149 por_dig_0.cnt_por\[0\] por_dig_0.net24 0.411329f
C1150 a_38146_31429# dvdd 0.163959f
C1151 por_dig_0.net24 a_35699_33819# 0.166861f
C1152 por_dig_0.cnt_por\[1\] a_37584_35389# 0.160237f
C1153 por_dig_0.cnt_rsb_stg1 force_dis_rc_osc 0.23536f
C1154 a_40247_24823# dvdd 0.543199f
C1155 por_ana_0.comparator_1.ena_b por_ana_0.comparator_1.vn 1.12092f
C1156 por porb 0.705431f
C1157 avss force_short_oneshot 0.642954f
C1158 por_dig_0.net22 por_dig_0._011_ 0.270877f
C1159 por_dig_0.net29 por_dig_0.net30 0.128046f
C1160 a_36494_35091# a_37409_35463# 0.125324f
C1161 a_14006_6535# avss 0.466415f
C1162 a_37688_33997# dvdd 0.142441f
C1163 por_dig_0.net25 a_35740_31277# 0.152281f
C1164 a_34719_23593# avdd 0.607928f
C1165 por_dig_0.net10 a_31413_29619# 0.200511f
C1166 a_33926_22885# a_34294_21903# 0.138963f
C1167 por_dig_0.net21 por_dig_0.net33 0.45707f
C1168 a_33444_31037# dvdd 0.347888f
C1169 por_dig_0._020_ dvdd 0.524414f
C1170 por_dig_0.clknet_0_osc_ck por_dig_0.net19 0.208482f
C1171 por_ana_0.comparator_1.vnn por_ana_0.comparator_1.vm 0.563119f
C1172 por_ana_0.schmitt_trigger_0.in por_ana_0.rstring_mux_0.vtrip_decoded_avdd[1] 0.133642f
C1173 a_31009_22637# por_ana_0.rstring_mux_0.vtrip_decoded_avdd[0] 0.135959f
C1174 a_33821_36551# dvdd 0.300009f
C1175 a_26785_24371# avdd 0.420074f
C1176 a_17398_35244# avss 0.460203f
C1177 a_37046_32915# dvdd 0.559204f
C1178 a_41694_2760# a_41694_2004# 0.296258f
C1179 por_dig_0.net24 a_36844_35463# 0.226729f
C1180 por_dig_0.cnt_st\[0\] por_dig_0._040_ 0.218954f
C1181 avdd itest 4.20531f
C1182 por_ana_0.comparator_1.vn vin 0.998331f
C1183 a_30495_23593# dvdd 0.104499f
C1184 por_ana_0.rstring_mux_0.otrip_decoded_avdd[0] avdd 1.34894f
C1185 por_dig_0._017_ por_dig_0._009_ 0.246785f
C1186 por_dig_0._010_ dvdd 0.406243f
C1187 por_ana_0.schmitt_trigger_0.in por_ana_0.rstring_mux_0.otrip_decoded_avdd[6] 0.105908f
C1188 por_dig_0.cnt_por\[0\] por_dig_0._051_ 0.154781f
C1189 por_dig_0.net23 a_36100_32517# 0.11288f
C1190 a_15518_6535# a_16274_6535# 0.296258f
C1191 a_33162_35603# dvdd 0.204284f
C1192 por_dig_0.cnt_por\[1\] a_35592_36286# 0.189554f
C1193 por_dig_0._052_ dvdd 0.855873f
C1194 a_24673_24371# por_ana_0.rstring_mux_0.otrip_decoded_avdd[3] 0.13699f
C1195 por_ana_0.comparator_1.vn por_ana_0.comparator_1.n0 1.97068f
C1196 por_dig_0._033_ por_dig_0.cnt_por\[2\] 0.119988f
C1197 a_38145_34375# dvdd 0.308049f
C1198 a_32464_32915# a_32630_32915# 0.610077f
C1199 a_35666_35629# a_36234_35871# 0.175891f
C1200 a_28383_21859# dvdd 0.104499f
C1201 por_dig_0.net6 por_dig_0.net12 0.154668f
C1202 por_dig_0.net25 a_37138_30189# 0.584861f
C1203 por_dig_0._034_ por_dig_0._035_ 0.59727f
C1204 por_dig_0.net24 a_33474_35059# 0.170223f
C1205 a_23366_22885# a_23466_22973# 0.40546f
C1206 por_dig_0.otrip_decoded[4] otrip[1] 0.234639f
C1207 a_36328_29645# dvdd 0.338518f
C1208 a_19676_13935# dvdd 0.401085f
C1209 a_18910_35244# a_19666_35244# 0.296258f
C1210 a_7835_22912# avss 0.471774f
C1211 a_38250_24707# dvdd 0.241639f
C1212 a_34946_30431# dvdd 0.201345f
C1213 a_3677_15512# a_4433_15512# 0.296258f
C1214 a_38518_23637# avdd 0.143323f
C1215 a_32607_21859# a_32182_21903# 0.460766f
C1216 por_dig_0._036_ a_36382_31795# 0.114183f
C1217 por_dig_0._035_ dvdd 0.748191f
C1218 a_32906_35091# a_33256_35463# 0.229804f
C1219 por_dig_0.net34 a_37751_31251# 0.148464f
C1220 por_dig_0.net24 por_dig_0._002_ 0.137441f
C1221 por_dig_0.force_pdnb por_dig_0.otrip_decoded[4] 0.109883f
C1222 por_ana_0.sky130_fd_sc_hd__inv_4_4.Y por 1.48351f
C1223 a_35958_31519# a_35740_31277# 0.209641f
C1224 a_35468_30163# a_35293_30189# 0.233657f
C1225 por_dig_0._019_ por_dig_0.net22 1.1086f
C1226 a_37345_24371# avdd 0.420074f
C1227 a_31914_22973# a_32607_21859# 0.264594f
C1228 por_dig_0.osc_ena por_dig_0.otrip_decoded[2] 0.116123f
C1229 por_dig_0._045_ a_37751_31251# 0.255891f
C1230 a_37798_33971# dvdd 0.224193f
C1231 a_20044_27844# avss 0.460231f
C1232 a_25863_32638# dvdd 0.175014f
C1233 por_dig_0.clknet_1_1__leaf_osc_ck a_36880_33453# 0.261973f
C1234 por_dig_0._053_ a_33896_35603# 0.13875f
C1235 por_dig_0.cnt_st\[4\] dvdd 1.56926f
C1236 por_dig_0.net16 a_36512_28013# 0.174696f
C1237 a_35930_6535# a_36686_6535# 0.296258f
C1238 a_35450_35124# dvdd 0.151751f
C1239 por_dig_0._033_ por_dig_0.cnt_por\[4\] 1.18984f
C1240 a_31360_31827# dvdd 0.458094f
C1241 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[0] por_ana_0.rstring_mux_0.vtrip_decoded_b_avdd[0] 0.574058f
C1242 a_2543_22912# avss 0.776278f
C1243 a_34026_24707# a_34719_23593# 0.264594f
C1244 por_dig_0._014_ a_34496_29645# 0.133811f
C1245 a_38444_28013# dvdd 0.296904f
C1246 a_32607_23593# avdd 0.607928f
C1247 a_25578_24707# a_26271_23593# 0.264594f
C1248 por_dig_0.net25 por_dig_0.clknet_1_0__leaf_osc_ck 0.242838f
C1249 por_dig_0.clknet_1_0__leaf_osc_ck por_dig_0.net28 0.206366f
C1250 a_32182_21903# dvdd 0.176016f
C1251 a_29802_24707# a_31009_24371# 0.28899f
C1252 a_34796_13935# avss 0.525451f
C1253 por_dig_0.net20 por_dig_0._016_ 0.577487f
C1254 por_dig_0.otrip_decoded[3] avdd 0.512716f
C1255 a_31802_32909# a_31908_32909# 0.419086f
C1256 a_14752_27844# avss 0.4604f
C1257 por_dig_0.cnt_st\[2\] por_dig_0._002_ 0.225497f
C1258 por_dig_0._001_ a_38957_32883# 0.118387f
C1259 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[2] avss 1.41004f
C1260 por_ana_0.rc_osc_0.vr a_19094_3138# 0.301135f
C1261 a_27958_21903# avdd 0.143952f
C1262 a_31984_31821# dvdd 0.134504f
C1263 dvdd isrc_sel 1.41732f
C1264 a_36696_30739# a_36862_30739# 0.701158f
C1265 por_dig_0.cnt_st\[3\] por_dig_0._003_ 0.201306f
C1266 por_dig_0._032_ dvdd 1.69377f
C1267 a_38926_33453# a_39162_33453# 0.22264f
C1268 a_21188_13935# a_21944_13935# 0.296258f
C1269 por_dig_0.clknet_1_0__leaf_osc_ck a_31526_31827# 0.42358f
C1270 por_dig_0.cnt_por\[8\] por_dig_0.cnt_rsb 0.304786f
C1271 por_dig_0._029_ a_38957_32883# 0.132266f
C1272 por_dig_0._004_ a_36862_30739# 0.230258f
C1273 por_dig_0.osc_ena avss 1.09147f
C1274 por_ana_0.rstring_mux_0.otrip_decoded_avdd[7] dvdd 0.291125f
C1275 a_31009_22637# avdd 0.421965f
C1276 por_ana_0.vl dvdd 1.79916f
C1277 por_dig_0.cnt_por\[0\] a_35500_35629# 0.627353f
C1278 a_26288_32594# dvdd 0.103629f
C1279 por_ana_0.schmitt_trigger_0.in por_ana_0.rstring_mux_0.otrip_decoded_avdd[0] 0.260407f
C1280 por_dig_0.net10 dvdd 0.373517f
C1281 a_32094_31795# por_dig_0.net8 0.170638f
C1282 a_33474_36147# a_33256_36551# 0.209641f
C1283 por_dig_0.net4 por_dig_0._026_ 0.132464f
C1284 por_dig_0.clknet_0_osc_ck por_dig_0._035_ 0.118086f
C1285 a_38136_33213# a_37961_33287# 0.233657f
C1286 por_dig_0.cnt_por\[7\] por_dig_0.cnt_por\[4\] 0.166092f
C1287 por_dig_0.net31 por_dig_0._000_ 0.159833f
C1288 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[1] por_ana_0.rstring_mux_0.vtrip_decoded_b_avdd[1] 0.572131f
C1289 a_31615_33705# a_31932_33595# 0.102355f
C1290 a_38500_31251# dvdd 0.289617f
C1291 a_35030_28557# dvdd 0.157993f
C1292 por_dig_0.otrip_decoded[7] a_27590_24619# 0.242839f
C1293 por_ana_0.rstring_mux_0.otrip_decoded_avdd[4] dvdd 0.266045f
C1294 avss porb_h 1.99008f
C1295 a_35390_31277# dvdd 0.578182f
C1296 por_dig_0.clknet_1_0__leaf_osc_ck por_dig_0.cnt_rsb 0.156434f
C1297 a_29504_13935# avss 0.465554f
C1298 por_dig_0._001_ dvdd 0.34437f
C1299 a_38943_23593# dvdd 0.106931f
C1300 por_dig_0._001_ a_37046_33453# 0.224572f
C1301 por_dig_0._046_ a_35040_34587# 0.146591f
C1302 por_dig_0.cnt_por\[9\] por_dig_0._037_ 0.184395f
C1303 a_5189_15512# avss 0.472978f
C1304 por_dig_0.cnt_por\[1\] por_dig_0._005_ 0.339053f
C1305 a_14752_27844# ibg_200n 0.350944f
C1306 a_29702_24619# dvdd 0.379209f
C1307 por_dig_0._029_ dvdd 0.3575f
C1308 por_dig_0.cnt_st\[0\] por_dig_0.cnt_st\[3\] 0.196921f
C1309 a_36972_30189# a_37138_30189# 0.615349f
C1310 por_dig_0.net25 a_36305_31277# 0.220031f
C1311 a_40247_24823# avdd 0.183326f
C1312 por_ana_0.rc_osc_0.vr dvdd 1.39451f
C1313 a_32740_36179# por_dig_0._007_ 0.173269f
C1314 por_dig_0.net32 dvdd 0.346025f
C1315 a_34098_30707# dvdd 1.28208f
C1316 por_dig_0.otrip_decoded[0] avss 0.134228f
C1317 a_30638_6535# a_31394_6535# 0.296258f
C1318 por_ana_0.sky130_fd_sc_hvl__lsbufhv2lv_1_1.X isrc_sel 0.130306f
C1319 por_dig_0._006_ a_36749_35451# 0.157737f
C1320 por_dig_0._048_ dvdd 0.797628f
C1321 por_dig_0.net26 a_31932_31419# 0.247151f
C1322 por_ana_0.rstring_mux_0.otrip_decoded_b_avdd[4] avss 0.36282f
C1323 por_dig_0.cnt_por\[2\] dvdd 1.23045f
C1324 a_27690_24707# avdd 0.863296f
C1325 a_37442_6535# avss 0.466333f
C1326 por_dig_0.net17 a_35960_29101# 0.171361f
C1327 por_dig_0.cnt_por\[0\] por_dig_0._049_ 0.141758f
C1328 avss startup_timed_out 0.266579f
C1329 avss osc_ck 3.89704f
C1330 a_37396_33287# dvdd 0.194667f
C1331 a_33926_22885# a_34026_22973# 0.40546f
C1332 por_dig_0.por_unbuf dvdd 3.21497f
C1333 a_19094_2382# a_19094_1626# 0.296258f
C1334 por_ana_0.vl por_ana_0.sky130_fd_sc_hvl__lsbufhv2lv_1_1.X 0.679849f
C1335 por_dig_0.net24 a_37409_35463# 0.231419f
C1336 por_ana_0.rstring_mux_0.otrip_decoded_avdd[3] vin 0.880782f
C1337 por_ana_0.rstring_mux_0.otrip_decoded_b_avdd[1] avdd 0.904297f
C1338 por_ana_0.rstring_mux_0.otrip_decoded_avdd[7] por_ana_0.rstring_mux_0.vtrip_decoded_avdd[0] 0.333912f
C1339 por_ana_0.rstring_mux_0.otrip_decoded_b_avdd[4] por_ana_0.rstring_mux_0.vtrip4 0.192181f
C1340 por_ana_0.comparator_1.n0 vin 0.567277f
C1341 por_dig_0.net24 a_35500_35629# 0.297288f
C1342 a_22700_13935# avss 0.465068f
C1343 a_32607_23593# a_32182_23637# 0.460766f
C1344 por_dig_0.net25 a_37212_31111# 0.155202f
C1345 por_dig_0.net22 por_dig_0._020_ 0.374976f
C1346 por_dig_0._047_ por_dig_0._024_ 0.307496f
C1347 por_dig_0.net21 por_dig_0._041_ 0.156591f
C1348 por_ana_0.rstring_mux_0.otrip_decoded_avdd[4] por_ana_0.rstring_mux_0.otrip_decoded_b_avdd[3] 0.155509f
C1349 por_dig_0._046_ a_35704_35124# 0.191904f
C1350 por_dig_0.clknet_1_0__leaf_osc_ck a_36696_30739# 0.405188f
C1351 a_15896_13935# a_16652_13935# 0.296258f
C1352 por_dig_0.force_pdnb por_dig_0.otrip_decoded[7] 0.103464f
C1353 a_30495_23593# avdd 0.607928f
C1354 a_21254_24619# a_21622_23637# 0.138963f
C1355 pwup_filt otrip[0] 2.25878f
C1356 por_dig_0._036_ por_dig_0._031_ 0.15031f
C1357 por_ana_0.rstring_mux_0.vtrip_decoded_b_avdd[3] avss 0.362811f
C1358 por_dig_0.net5 a_35030_28557# 0.122572f
C1359 a_32464_32915# a_32980_33287# 0.10241f
C1360 a_32630_32915# a_33198_32883# 0.175891f
C1361 por_dig_0.cnt_st\[0\] por_dig_0._030_ 0.183418f
C1362 a_36234_35871# a_36016_35629# 0.209641f
C1363 a_32464_32915# dvdd 0.437332f
C1364 a_32150_6535# avss 0.466333f
C1365 por_ana_0.rstring_mux_0.vtrip_decoded_b_avdd[0] avdd 0.903548f
C1366 por_dig_0.net25 a_37488_30189# 0.186849f
C1367 a_23466_22973# a_24673_22637# 0.28899f
C1368 por_dig_0.net24 a_33996_35389# 0.310206f
C1369 a_23366_22885# dvdd 0.380879f
C1370 por_dig_0.net20 por_dig_0._037_ 0.208515f
C1371 por_dig_0.clknet_1_0__leaf_osc_ck a_36972_30189# 0.25213f
C1372 a_28383_21859# avdd 0.607928f
C1373 por_dig_0.cnt_por\[2\] por_dig_0.cnt_por\[3\] 0.929531f
C1374 a_21178_35244# osc_ck 0.160246f
C1375 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[2] por_ana_0.rstring_mux_0.vtrip2 0.4803f
C1376 por_ana_0.rstring_mux_0.otrip_decoded_avdd[1] dvdd 0.261341f
C1377 por_dig_0.cnt_por\[4\] dvdd 1.22567f
C1378 a_17408_13935# avss 0.465068f
C1379 a_35612_33595# a_36880_33453# 0.104154f
C1380 a_35468_30163# dvdd 0.34776f
C1381 a_4055_22912# a_4811_22912# 0.296258f
C1382 a_21354_22973# avdd 0.864385f
C1383 a_32352_32731# dvdd 0.132472f
C1384 a_19676_13935# avdd 0.146832f
C1385 a_32812_30733# dvdd 0.142876f
C1386 por_dig_0.net15 a_34265_27987# 0.179572f
C1387 a_32906_35091# a_33821_35463# 0.124988f
C1388 por_dig_0._047_ dvdd 0.606856f
C1389 por_dig_0.clknet_0_osc_ck a_34098_30707# 0.316023f
C1390 a_32701_28531# por_dig_0.otrip_decoded[1] 0.158695f
C1391 a_38250_24707# avdd 0.863819f
C1392 a_33752_28013# dvdd 0.299904f
C1393 por_dig_0.osc_ena por_dig_0.otrip_decoded[4] 0.107181f
C1394 por_dig_0._033_ por_dig_0._017_ 0.209169f
C1395 por_dig_0.cnt_st\[0\] por_dig_0._000_ 0.429422f
C1396 por_dig_0.net6 a_35130_28673# 0.11344f
C1397 por_dig_0.net25 a_37614_33695# 0.170725f
C1398 por_ana_0.rstring_mux_0.otrip_decoded_avdd[5] por_ana_0.rstring_mux_0.otrip_decoded_b_avdd[4] 0.155007f
C1399 por_ana_0.rstring_mux_0.vtrip_decoded_b_avdd[7] avdd 0.839308f
C1400 por_dig_0.net2 pwup_filt 0.145998f
C1401 a_23834_6535# a_24590_6535# 0.296258f
C1402 a_31802_32909# dvdd 0.283022f
C1403 por_dig_0.cnt_st\[1\] por_dig_0._029_ 0.349474f
C1404 a_25346_6535# avss 0.466333f
C1405 a_38926_33453# dvdd 0.322764f
C1406 por_dig_0.net24 a_32088_33690# 0.166183f
C1407 a_25863_32638# avdd 0.138798f
C1408 por_dig_0._038_ pwup_filt 0.160523f
C1409 a_39417_31795# force_short_oneshot 0.180322f
C1410 por_dig_0.net25 por_dig_0.net27 0.390604f
C1411 a_36308_13935# a_37064_13935# 0.296258f
C1412 por_dig_0._023_ por_dig_0._011_ 0.13851f
C1413 a_32094_31795# dvdd 0.204605f
C1414 por_dig_0.cnt_por\[6\] por_dig_0._011_ 1.09895f
C1415 por_dig_0._036_ por_dig_0.cnt_rsb 0.140682f
C1416 a_16264_27844# a_17020_27844# 0.296258f
C1417 por_dig_0.net26 por_dig_0._012_ 0.665859f
C1418 a_34573_28557# a_34750_28557# 0.134298f
C1419 dvdd pwup_filt 2.84251f
C1420 a_22561_24371# por_ana_0.rstring_mux_0.otrip_decoded_avdd[1] 0.13699f
C1421 a_34212_30189# a_34378_30189# 0.830627f
C1422 a_36381_36691# por_dig_0.por_unbuf 0.15489f
C1423 por_dig_0._008_ a_32906_35091# 0.223208f
C1424 por_dig_0._009_ a_35612_33595# 0.61908f
C1425 a_32740_36179# dvdd 0.538291f
C1426 por_dig_0._003_ a_37393_30189# 0.170087f
C1427 por_dig_0._027_ dvdd 0.74648f
C1428 por_dig_0.force_pdnb a_38150_22885# 0.243342f
C1429 a_33926_22885# dvdd 0.382644f
C1430 a_32182_21903# avdd 0.143952f
C1431 por_dig_0.cnt_por\[6\] por_dig_0.cnt_por\[5\] 0.146019f
C1432 a_36696_30739# a_37212_31111# 0.107135f
C1433 a_36862_30739# a_37430_30707# 0.174561f
C1434 a_36952_35085# dvdd 0.140723f
C1435 a_39162_33453# a_39268_33453# 0.419086f
C1436 por_dig_0.clknet_1_0__leaf_osc_ck por_dig_0.net8 0.54455f
C1437 dvdd force_ena_rc_osc 0.457473f
C1438 por_ana_0.sky130_fd_sc_hvl__inv_1_0.A a_26802_33372# 0.141238f
C1439 a_20054_6535# avss 0.466333f
C1440 a_31914_22973# avdd 0.863791f
C1441 por_ana_0.rstring_mux_0.otrip_decoded_b_avdd[5] vin 0.340862f
C1442 por_dig_0.net24 a_32704_31111# 0.156309f
C1443 a_22047_23593# a_21622_23637# 0.460766f
C1444 por_dig_0.clknet_0_osc_ck por_dig_0.cnt_por\[4\] 0.417979f
C1445 por_dig_0._016_ por_dig_0._053_ 0.208828f
C1446 avdd isrc_sel 0.517827f
C1447 a_37064_34003# a_37230_34003# 0.616545f
C1448 a_36234_35871# dvdd 0.213265f
C1449 por_dig_0.net24 a_33996_36477# 0.288614f
C1450 por_dig_0._044_ a_39077_31527# 0.17235f
C1451 por_dig_0.cnt_por\[7\] por_dig_0.cnt_por\[8\] 0.193184f
C1452 por_ana_0.rstring_mux_0.otrip_decoded_avdd[7] avdd 1.81983f
C1453 por_dig_0.net23 por_dig_0._048_ 0.365535f
C1454 por_ana_0.vl avdd 2.52471f
C1455 por_dig_0.net23 por_dig_0.cnt_por\[2\] 0.203161f
C1456 por_dig_0.net20 por_dig_0.net24 0.306376f
C1457 a_26288_32594# avdd 0.602828f
C1458 a_31893_33721# a_32088_33690# 0.229804f
C1459 a_26785_22637# por_ana_0.rstring_mux_0.otrip_decoded_avdd[4] 0.136088f
C1460 por_dig_0.por_unbuf por_ana_0.sky130_fd_sc_hd__inv_4_1.A 0.44008f
C1461 a_21254_24619# a_21354_24707# 0.40546f
C1462 a_35740_31277# dvdd 0.209943f
C1463 por_dig_0._011_ a_31932_33595# 0.271131f
C1464 por_dig_0.otrip_decoded[3] otrip[2] 0.153226f
C1465 por_dig_0.net33 dvdd 0.200906f
C1466 por_dig_0._027_ por_dig_0.net30 0.288915f
C1467 por_dig_0.net8 a_31615_31529# 0.237905f
C1468 a_21622_23637# dvdd 0.169579f
C1469 por_dig_0.cnt_por\[0\] a_34672_35451# 0.213029f
C1470 por_ana_0.rstring_mux_0.otrip_decoded_avdd[4] avdd 1.52955f
C1471 por_dig_0._050_ por_dig_0._006_ 0.153395f
C1472 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[4] por_ana_0.rstring_mux_0.vtrip_decoded_b_avdd[4] 0.572505f
C1473 a_18542_6535# a_19298_6535# 0.296258f
C1474 por_dig_0._029_ por_dig_0._040_ 0.204308f
C1475 a_14762_6535# avss 0.466333f
C1476 a_37138_30189# a_37706_30431# 0.17072f
C1477 a_36972_30189# a_37488_30189# 0.110816f
C1478 a_38943_23593# avdd 0.612302f
C1479 a_36862_30739# dvdd 0.58068f
C1480 a_31016_13935# a_31772_13935# 0.296258f
C1481 por_dig_0._019_ por_dig_0.cnt_por\[6\] 0.45193f
C1482 por_dig_0.otrip_decoded[2] otrip[0] 0.65194f
C1483 a_36880_32915# a_37046_32915# 0.60715f
C1484 a_31412_31251# a_31615_31529# 0.233657f
C1485 a_29702_24619# avdd 0.206171f
C1486 a_34026_22973# a_35233_22637# 0.28899f
C1487 a_18154_35244# avss 0.460203f
C1488 por_dig_0._011_ por_dig_0._021_ 0.100483f
C1489 a_37961_33287# dvdd 0.293626f
C1490 a_33155_28640# dvdd 0.192737f
C1491 por_dig_0.net7 por_dig_0.net15 0.304907f
C1492 a_32794_33971# dvdd 0.237827f
C1493 por_dig_0.net32 por_dig_0._013_ 0.149461f
C1494 a_36512_28013# por_dig_0.otrip_decoded[5] 0.177464f
C1495 a_31728_32365# a_31894_32365# 0.901539f
C1496 por_dig_0.net25 a_37777_31111# 0.241505f
C1497 a_6701_15512# a_7457_15512# 0.296258f
C1498 por_dig_0.por_unbuf avdd 0.300005f
C1499 a_31592_30965# por_dig_0._038_ 0.100645f
C1500 por_dig_0.net23 por_dig_0.cnt_por\[4\] 0.146665f
C1501 a_37138_30189# dvdd 0.280398f
C1502 a_34114_35879# dvdd 0.294002f
C1503 por_dig_0._048_ por_dig_0.net22 0.314042f
C1504 a_35092_33427# a_35295_33705# 0.233657f
C1505 a_36512_28013# dvdd 0.272899f
C1506 por_dig_0.osc_ena por_dig_0.otrip_decoded[7] 0.107303f
C1507 por_dig_0.clknet_1_1__leaf_osc_ck por_dig_0._007_ 0.291644f
C1508 por_ana_0.comparator_1.n0 por_ana_0.dcomp3v3 0.945307f
C1509 a_31728_32365# dvdd 0.4269f
C1510 a_31592_30965# dvdd 0.149647f
C1511 a_21254_22885# a_21622_21903# 0.138963f
C1512 a_32464_32915# a_33545_33287# 0.102355f
C1513 a_33198_32883# a_32980_33287# 0.209641f
C1514 a_27690_22973# a_28383_21859# 0.264594f
C1515 por_dig_0._017_ dvdd 0.304727f
C1516 por_dig_0.net25 a_38053_30189# 0.285741f
C1517 a_33198_32883# dvdd 0.208252f
C1518 por_dig_0.net15 dvdd 0.495811f
C1519 por_dig_0._012_ a_32149_32365# 0.172541f
C1520 a_32354_30739# a_32704_31111# 0.219633f
C1521 a_8591_22912# avss 0.47927f
C1522 avss otrip[0] 0.209734f
C1523 por_dig_0.cnt_por\[8\] dvdd 0.604986f
C1524 por_ana_0.comparator_0.vnn por_ana_0.comparator_0.vn 0.298803f
C1525 por_dig_0._017_ a_35100_32339# 0.194982f
C1526 a_36122_30341# dvdd 0.189224f
C1527 por_dig_0._019_ por_dig_0._011_ 0.139962f
C1528 a_23366_22885# avdd 0.207177f
C1529 por_dig_0.net2 a_31776_29864# 0.139807f
C1530 por_dig_0.cnt_st\[1\] por_dig_0.net33 0.358355f
C1531 a_36480_31251# a_36305_31277# 0.233657f
C1532 a_36122_30341# a_36218_30163# 0.419086f
C1533 por_dig_0.otrip_decoded[2] dvdd 1.04175f
C1534 por_ana_0.rstring_mux_0.otrip_decoded_avdd[1] avdd 1.72246f
C1535 por_dig_0.net4 por_dig_0._039_ 0.170358f
C1536 por_dig_0.net24 por_dig_0.net26 0.820732f
C1537 a_13250_6535# a_14006_6535# 0.296258f
C1538 a_21354_24707# a_22047_23593# 0.264594f
C1539 por_dig_0.cnt_por\[4\] por_dig_0._013_ 0.166132f
C1540 a_20800_27844# avss 0.4604f
C1541 por_ana_0.schmitt_trigger_0.in por_ana_0.rstring_mux_0.otrip_decoded_avdd[7] 0.126209f
C1542 force_dis_rc_osc pwup_filt 0.123157f
C1543 por_dig_0.net25 a_38136_33427# 0.306564f
C1544 por_ana_0.vl por_ana_0.schmitt_trigger_0.in 0.489542f
C1545 por_dig_0.net5 a_33155_28640# 0.178157f
C1546 a_31360_33997# por_dig_0.net1 0.110039f
C1547 a_24212_13935# a_24968_13935# 0.296258f
C1548 por_dig_0.clknet_1_0__leaf_osc_ck dvdd 4.98489f
C1549 a_34828_29253# por_dig_0.net7 0.121927f
C1550 por_dig_0.cnt_por\[9\] por_dig_0._015_ 0.287681f
C1551 por_dig_0.cnt_por\[10\] a_35224_31277# 0.507132f
C1552 por_ana_0.vl por_dig_0.otrip_decoded[1] 0.118122f
C1553 a_39268_33453# dvdd 0.182312f
C1554 por_dig_0.cnt_por\[9\] por_dig_0._028_ 0.180564f
C1555 por_dig_0._019_ por_dig_0.cnt_por\[5\] 0.481699f
C1556 por_dig_0.net22 por_dig_0.cnt_por\[4\] 0.194538f
C1557 a_31776_29864# dvdd 0.221645f
C1558 a_34265_27987# por_dig_0.otrip_decoded[4] 0.184294f
C1559 a_33774_31821# dvdd 0.264292f
C1560 a_28383_23593# dvdd 0.104499f
C1561 por_dig_0.force_pdnb force_pdn 0.61636f
C1562 a_34486_33703# dvdd 0.192605f
C1563 por_dig_0.por_unbuf por_ana_0.schmitt_trigger_0.m 0.13807f
C1564 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[0] por_ana_0.rstring_mux_0.otrip_decoded_b_avdd[7] 0.154952f
C1565 por_dig_0._047_ por_dig_0.net22 0.171048f
C1566 por_ana_0.schmitt_trigger_0.in por_ana_0.rstring_mux_0.otrip_decoded_avdd[4] 0.101976f
C1567 force_ena_rc_osc force_dis_rc_osc 2.4551f
C1568 a_3299_22912# avss 0.484544f
C1569 a_16642_35244# a_17398_35244# 0.296258f
C1570 por_dig_0._031_ por_dig_0._037_ 0.137183f
C1571 a_39887_23089# por_ana_0.dcomp3v3uv 0.223996f
C1572 a_34387_32909# osc_ck 0.383921f
C1573 por_dig_0._049_ por_dig_0._050_ 0.195476f
C1574 por_ana_0.comparator_0.vn avss 8.98681f
C1575 a_33896_35603# dvdd 0.182764f
C1576 por_dig_0.cnt_por\[1\] por_dig_0.cnt_por\[2\] 0.319882f
C1577 por_dig_0.net4 por_dig_0.net21 0.586782f
C1578 por_ana_0.rstring_mux_0.vtop osc_ck 0.109483f
C1579 a_31814_24619# a_31914_24707# 0.40546f
C1580 por_dig_0.net4 por_dig_0.net25 0.297337f
C1581 a_38518_21903# dvdd 0.17571f
C1582 a_34212_30189# a_34728_30189# 0.115353f
C1583 por_dig_0.net25 por_dig_0._042_ 0.293827f
C1584 por_dig_0.clknet_0_osc_ck por_dig_0._017_ 0.23129f
C1585 por_dig_0.cnt_por\[5\] a_36100_32517# 0.247747f
C1586 por_dig_0.net6 a_33971_28557# 0.245434f
C1587 a_35552_13935# avss 0.525451f
C1588 a_26271_21859# dvdd 0.104499f
C1589 a_31615_31529# dvdd 0.296082f
C1590 a_15508_27844# avss 0.460231f
C1591 por_dig_0.net6 por_dig_0.net7 2.14791f
C1592 por_dig_0.net5 por_dig_0.net15 0.166483f
C1593 avdd pwup_filt 0.206066f
C1594 por_dig_0.net25 a_34212_30189# 0.296275f
C1595 a_34828_29253# dvdd 0.23356f
C1596 a_37430_30707# a_37212_31111# 0.209641f
C1597 a_36696_30739# a_37777_31111# 0.102355f
C1598 por_ana_0.comparator_0.vn vbg_1v2 0.728008f
C1599 a_35040_34587# dvdd 0.150022f
C1600 avss dvdd 11.0009f
C1601 por_dig_0.clknet_1_1__leaf_osc_ck por_dig_0._034_ 0.647828f
C1602 a_33926_22885# avdd 0.207177f
C1603 a_35295_33705# dvdd 0.286434f
C1604 a_33774_31821# a_34010_31821# 0.22264f
C1605 por_dig_0.net24 a_33269_31111# 0.227562f
C1606 por_ana_0.rstring_mux_0.vtrip0 a_25346_6535# 0.298434f
C1607 a_33662_6535# a_34418_6535# 0.296258f
C1608 a_37064_34003# por_dig_0.net25 0.307776f
C1609 a_36756_35603# dvdd 0.451645f
C1610 a_22047_21859# a_21622_21903# 0.460766f
C1611 por_ana_0.sky130_fd_sc_hd__inv_4_0.Y pwup_filt 1.47962f
C1612 avdd force_ena_rc_osc 0.215182f
C1613 por_dig_0.net24 a_37614_32883# 0.159851f
C1614 por_dig_0.net5 por_dig_0.otrip_decoded[2] 0.108043f
C1615 por_dig_0.net4 osc_ck 0.105559f
C1616 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[1] por_ana_0.rstring_mux_0.vtrip_decoded_b_avdd[0] 0.155269f
C1617 dvdd vbg_1v2 0.345536f
C1618 a_21354_24707# a_22561_24371# 0.28899f
C1619 a_36305_31277# dvdd 0.293953f
C1620 por_dig_0.clknet_1_1__leaf_osc_ck dvdd 4.20163f
C1621 por_dig_0.net9 por_dig_0.net3 0.165675f
C1622 por_ana_0.dcomp3v3uv avss 7.277201f
C1623 a_35960_29101# dvdd 0.233833f
C1624 por_dig_0.net33 por_dig_0._040_ 0.202586f
C1625 por_dig_0.net1 dvdd 0.518015f
C1626 a_30260_13935# avss 0.465525f
C1627 a_33896_35603# por_dig_0.cnt_por\[3\] 0.186138f
C1628 por_dig_0.net6 dvdd 3.36578f
C1629 por_dig_0.net8 a_31932_31419# 0.321184f
C1630 a_35217_28013# a_35394_28013# 0.134298f
C1631 a_25846_23637# dvdd 0.169343f
C1632 por_dig_0.cnt_por\[0\] por_dig_0._046_ 0.377192f
C1633 por_dig_0.net24 por_dig_0._009_ 0.301503f
C1634 a_5945_15512# avss 0.472978f
C1635 por_ana_0.vl por_ana_0.sky130_fd_sc_hd__inv_4_3.Y 0.396075f
C1636 a_18920_13935# a_19676_13935# 0.296258f
C1637 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[3] avss 1.48249f
C1638 por_ana_0.dcomp3v3uv vbg_1v2 0.3098f
C1639 a_21622_23637# avdd 0.143029f
C1640 a_36972_30189# a_38053_30189# 0.102325f
C1641 a_37706_30431# a_37488_30189# 0.209641f
C1642 a_37212_31111# dvdd 0.204073f
C1643 por_dig_0.otrip_decoded[4] otrip[0] 0.176593f
C1644 a_36880_32915# a_37396_33287# 0.102946f
C1645 dvdd ibg_200n 0.231478f
C1646 a_31615_31529# a_31893_31545# 0.125324f
C1647 a_31009_24371# avdd 0.420074f
C1648 a_36649_28789# dvdd 0.180646f
C1649 a_38198_6535# avss 0.466415f
C1650 por_ana_0.comparator_0.vn por_ana_0.comparator_0.vm 4.66142f
C1651 por_ana_0.rstring_mux_0.otrip_decoded_b_avdd[3] avss 0.362817f
C1652 por_dig_0._034_ por_dig_0._036_ 0.10904f
C1653 por_ana_0.schmitt_trigger_0.in por_ana_0.rstring_mux_0.otrip_decoded_avdd[1] 0.556851f
C1654 por_dig_0.net20 por_dig_0._049_ 0.127006f
C1655 por_dig_0._041_ dvdd 0.449082f
C1656 por_dig_0._033_ por_dig_0._016_ 0.410232f
C1657 por_dig_0._042_ por_dig_0._044_ 0.208006f
C1658 a_34290_28557# dvdd 0.208585f
C1659 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[0] avss 1.37856f
C1660 por_ana_0.rstring_mux_0.otrip_decoded_b_avdd[0] avdd 0.870606f
C1661 a_34828_29253# por_dig_0.net5 0.197275f
C1662 por_dig_0.net23 por_dig_0.cnt_por\[8\] 0.136855f
C1663 a_23456_13935# avss 0.465068f
C1664 a_31728_32365# a_32244_32365# 0.115353f
C1665 a_31894_32365# a_32462_32607# 0.184993f
C1666 a_7079_22912# a_7835_22912# 0.296258f
C1667 a_37488_30189# dvdd 0.210243f
C1668 por_ana_0.rstring_mux_0.otrip_decoded_avdd[5] dvdd 0.416917f
C1669 a_28383_23593# a_27958_23637# 0.460766f
C1670 a_32641_28013# a_32818_28013# 0.134298f
C1671 por_dig_0.cnt_por\[0\] a_35666_35629# 0.616013f
C1672 por_dig_0._036_ dvdd 2.73711f
C1673 por_ana_0.dcomp3v3 a_39888_24823# 0.204909f
C1674 por_dig_0._039_ por_dig_0._002_ 0.41148f
C1675 a_23366_24619# a_23734_23637# 0.138963f
C1676 a_35295_33705# a_35573_33721# 0.123255f
C1677 por_dig_0.net4 a_36696_30739# 0.290738f
C1678 a_32462_32607# dvdd 0.208034f
C1679 por_dig_0.net4 por_dig_0._004_ 0.142903f
C1680 por_ana_0.rstring_mux_0.vtrip_decoded_b_avdd[2] avss 0.362817f
C1681 por_dig_0._039_ por_dig_0.cnt_st\[2\] 0.268582f
C1682 a_40246_23089# dvdd 0.447991f
C1683 por_ana_0.rstring_mux_0.vtrip6 avdd 0.949337f
C1684 a_39077_31527# dvdd 0.25943f
C1685 a_36756_35603# a_36581_35629# 0.234322f
C1686 por_ana_0.rstring_mux_0.otrip_decoded_avdd[2] dvdd 0.255062f
C1687 a_32906_6535# avss 0.466333f
C1688 a_33720_33213# dvdd 0.369059f
C1689 por_dig_0._020_ por_dig_0._021_ 0.135272f
C1690 por_ana_0.rstring_mux_0.otrip_decoded_b_avdd[7] avdd 0.903548f
C1691 por_ana_0.rstring_mux_0.otrip_decoded_avdd[5] por_ana_0.dcomp3v3uv 0.213252f
C1692 a_32233_31643# dvdd 0.142104f
C1693 a_25478_22885# a_25578_22973# 0.40546f
C1694 por_dig_0.net5 por_dig_0.net6 1.84601f
C1695 por_dig_0.otrip_decoded[4] por_dig_0.otrip_decoded[5] 1.62547f
C1696 a_37789_31821# dvdd 0.269995f
C1697 a_37614_33695# dvdd 0.208584f
C1698 a_32354_30739# a_33269_31111# 0.125324f
C1699 a_19288_27844# a_20044_27844# 0.296258f
C1700 a_37046_33453# a_37614_33695# 0.186387f
C1701 por_ana_0.comparator_0.vnn por_ana_0.comparator_0.n0 0.428003f
C1702 por_dig_0.cnt_por\[9\] a_35556_29619# 0.304256f
C1703 a_36476_30163# dvdd 0.271959f
C1704 a_18164_13935# avss 0.465068f
C1705 a_24673_22637# avdd 0.421965f
C1706 por_dig_0.otrip_decoded[1] pwup_filt 1.49992f
C1707 por_dig_0.net24 osc_ck 0.216724f
C1708 a_33934_32615# dvdd 0.200694f
C1709 a_20432_13935# avdd 0.15041f
C1710 por_dig_0.cnt_por\[9\] a_34378_30189# 0.127581f
C1711 por_dig_0._007_ a_32906_36179# 0.282122f
C1712 por_dig_0.net27 dvdd 0.461572f
C1713 por_dig_0.net22 por_dig_0._017_ 0.173149f
C1714 por_dig_0.otrip_decoded[4] a_25478_22885# 0.260032f
C1715 por_ana_0.rstring_mux_0.otrip_decoded_avdd[2] por_ana_0.dcomp3v3uv 0.375655f
C1716 por_dig_0._013_ por_dig_0.cnt_por\[8\] 0.554099f
C1717 por_dig_0.otrip_decoded[4] dvdd 0.74407f
C1718 a_36218_30163# a_36476_30163# 0.22264f
C1719 a_13628_13935# a_14384_13935# 0.296258f
C1720 por_dig_0._008_ a_33161_35451# 0.171386f
C1721 a_37528_31527# dvdd 0.185004f
C1722 a_35960_29101# por_dig_0.otrip_decoded[6] 0.184577f
C1723 por_dig_0.net24 por_dig_0.cnt_rsb 0.18439f
C1724 por_dig_0.net28 a_31781_32187# 0.170162f
C1725 por_ana_0.rstring_mux_0.vtrip_decoded_b_avdd[6] avdd 0.904181f
C1726 por_dig_0.otrip_decoded[2] avdd 0.900195f
C1727 por_dig_0.net23 a_35040_34587# 0.219985f
C1728 por_dig_0.clknet_1_1__leaf_osc_ck a_36328_35091# 0.285795f
C1729 por_ana_0.rstring_mux_0.otrip_decoded_avdd[7] por_ana_0.rstring_mux_0.otrip_decoded_avdd[6] 1.12965f
C1730 a_35100_32339# por_dig_0.net27 0.215457f
C1731 a_39887_23089# avdd 0.538752f
C1732 a_36831_23593# a_36406_23637# 0.460766f
C1733 a_34116_31821# dvdd 0.18439f
C1734 por_ana_0.comparator_0.vnn avdd 37.3292f
C1735 por_dig_0.osc_ena force_pdn 0.339611f
C1736 por_dig_0.clknet_1_0__leaf_osc_ck por_dig_0._013_ 0.388397f
C1737 avss force_dis_rc_osc 0.350678f
C1738 a_40246_21893# a_39887_21959# 0.249269f
C1739 a_36138_24707# a_36831_23593# 0.264594f
C1740 por_dig_0.cnt_st\[1\] por_dig_0._041_ 0.176074f
C1741 por_dig_0._019_ por_dig_0._020_ 0.385183f
C1742 a_23366_24619# dvdd 0.385817f
C1743 a_31526_31827# a_31876_32199# 0.210696f
C1744 por_ana_0.comparator_0.n0 avss 4.20597f
C1745 a_28383_23593# avdd 0.607928f
C1746 a_31914_24707# a_33121_24371# 0.28899f
C1747 a_35224_31277# a_35390_31277# 0.608921f
C1748 a_34212_30189# a_35293_30189# 0.102355f
C1749 por_dig_0.net7 a_35674_28557# 0.178241f
C1750 por_dig_0.net22 por_dig_0.clknet_1_0__leaf_osc_ck 0.316984f
C1751 por_dig_0.net23 por_dig_0.clknet_1_1__leaf_osc_ck 0.251778f
C1752 por_dig_0.cnt_por\[5\] por_dig_0._035_ 0.184651f
C1753 a_21354_24707# avdd 0.865655f
C1754 por_dig_0._022_ dvdd 0.228553f
C1755 por_dig_0.net19 por_dig_0.cnt_por\[10\] 0.113765f
C1756 por_dig_0.por_unbuf por_ana_0.sky130_fd_sc_hd__inv_4_4.Y 0.414643f
C1757 a_31932_31419# dvdd 0.458117f
C1758 por_dig_0._033_ por_dig_0.net4 0.343499f
C1759 a_38518_21903# avdd 0.144336f
C1760 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A avss 4.17343f
C1761 por_ana_0.sky130_fd_sc_hvl__inv_1_0.A osc_ck 0.732369f
C1762 por_dig_0._019_ por_dig_0._010_ 0.243215f
C1763 por_ana_0.comparator_0.n0 vbg_1v2 0.692613f
C1764 a_21566_6535# a_22322_6535# 0.296258f
C1765 por_dig_0.otrip_decoded[6] por_ana_0.rstring_mux_0.otrip_decoded_avdd[5] 0.143657f
C1766 por_dig_0.net1 force_dis_rc_osc 0.17605f
C1767 pwup_filt porb 0.110486f
C1768 a_26271_21859# avdd 0.607928f
C1769 por_dig_0.otrip_decoded[4] por_ana_0.sky130_fd_sc_hvl__lsbufhv2lv_1_1.X 0.766371f
C1770 a_20810_6535# avss 0.466333f
C1771 a_25595_33708# a_26288_32594# 0.264594f
C1772 a_35233_22637# avdd 0.421965f
C1773 a_34010_31821# a_34116_31821# 0.419086f
C1774 a_35612_33595# dvdd 0.421433f
C1775 por_ana_0.rstring_mux_0.otrip_decoded_b_avdd[4] vin 0.340862f
C1776 por_dig_0.cnt_por\[6\] por_dig_0.net32 0.10714f
C1777 a_34040_13935# a_34796_13935# 0.296258f
C1778 por_dig_0.net20 a_36564_32339# 0.242368f
C1779 avdd avss 2.55669p
C1780 por_dig_0.clknet_0_osc_ck por_dig_0.net27 0.261082f
C1781 por_dig_0.net24 a_38136_33213# 0.270076f
C1782 a_34290_28557# a_34467_28557# 0.159555f
C1783 a_35674_28557# dvdd 0.156702f
C1784 por_ana_0.rstring_mux_0.vtrip4 avdd 0.416503f
C1785 por_dig_0.net34 dvdd 0.270051f
C1786 por_dig_0._016_ dvdd 0.491479f
C1787 por_dig_0._033_ por_dig_0.cnt_por\[0\] 0.429718f
C1788 por_dig_0._045_ dvdd 0.464749f
C1789 por_ana_0.rstring_mux_0.vtrip_decoded_b_avdd[2] por_ana_0.rstring_mux_0.vtrip2 0.190544f
C1790 por_dig_0.net8 a_32019_31643# 0.179916f
C1791 avdd vbg_1v2 10.8258f
C1792 a_30070_23637# dvdd 0.169343f
C1793 por_dig_0._025_ por_dig_0.cnt_por\[7\] 0.124044f
C1794 a_36494_35091# dvdd 0.403256f
C1795 a_19288_27844# osc_ck 0.346796f
C1796 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[4] por_ana_0.rstring_mux_0.vtrip_decoded_b_avdd[3] 0.155115f
C1797 por_dig_0.net4 por_dig_0.cnt_por\[7\] 0.519958f
C1798 por_dig_0.net11 a_38444_28013# 0.178319f
C1799 a_33926_24619# dvdd 0.441709f
C1800 a_37798_33971# a_37580_34375# 0.209641f
C1801 a_15518_6535# avss 0.466333f
C1802 por_dig_0.otrip_decoded[6] por_dig_0.otrip_decoded[4] 3.56664f
C1803 a_25846_23637# avdd 0.142934f
C1804 a_34580_34110# por_dig_0._022_ 0.136448f
C1805 a_37777_31111# dvdd 0.289725f
C1806 por_dig_0.net24 a_32630_32915# 0.62121f
C1807 a_36880_32915# a_37961_33287# 0.102355f
C1808 a_31893_31545# a_31932_31419# 0.900887f
C1809 a_31914_24707# avdd 0.863296f
C1810 force_short_oneshot otrip[1] 0.105227f
C1811 por_ana_0.comparator_0.vm por_ana_0.comparator_0.n0 2.61558f
C1812 a_18910_35244# avss 0.460203f
C1813 a_36038_22885# a_36138_22973# 0.40546f
C1814 a_32906_36179# dvdd 0.462191f
C1815 a_41694_2004# a_41694_1248# 0.296258f
C1816 a_34573_28557# dvdd 0.174251f
C1817 a_23466_22973# a_24159_21859# 0.264594f
C1818 avdd ibg_200n 2.33988f
C1819 por_dig_0.otrip_decoded[5] por_dig_0.otrip_decoded[7] 3.81635f
C1820 por_ana_0.sky130_fd_sc_hvl__inv_4_0.A avss 0.98945f
C1821 por_dig_0.cnt_por\[6\] por_dig_0.cnt_por\[4\] 0.140355f
C1822 por_ana_0.schmitt_trigger_0.in por_dig_0.otrip_decoded[2] 0.15479f
C1823 a_32462_32607# a_32244_32365# 0.209641f
C1824 a_31728_32365# a_32809_32365# 0.102355f
C1825 por_dig_0._012_ a_31894_32365# 0.637032f
C1826 a_38053_30189# dvdd 0.296302f
C1827 a_32740_35091# dvdd 0.475531f
C1828 a_39634_32615# dvdd 0.195911f
C1829 por_dig_0._016_ por_dig_0.cnt_por\[3\] 0.110428f
C1830 por_dig_0.otrip_decoded[1] por_dig_0.otrip_decoded[2] 2.20309f
C1831 por_dig_0.net13 a_33752_28013# 0.171599f
C1832 por_ana_0.schmitt_trigger_0.in por_ana_0.comparator_0.vnn 0.268371f
C1833 a_28383_21859# a_27958_21903# 0.460766f
C1834 a_16274_6535# a_17030_6535# 0.296258f
C1835 por_dig_0.net23 por_dig_0.net27 0.325932f
C1836 a_35573_33721# a_35612_33595# 0.616545f
C1837 a_38956_32339# dvdd 0.39818f
C1838 por_dig_0.net7 a_34615_28013# 0.207596f
C1839 por_dig_0.otrip_decoded[7] dvdd 0.65413f
C1840 por_ana_0.rstring_mux_0.otrip_decoded_avdd[5] avdd 1.80973f
C1841 a_32984_32339# dvdd 0.361337f
C1842 por_dig_0._012_ dvdd 1.14892f
C1843 por_dig_0._024_ por_dig_0._025_ 0.277436f
C1844 a_23366_22885# a_23734_21903# 0.138963f
C1845 a_33720_33213# a_33545_33287# 0.233657f
C1846 a_38943_21859# dvdd 0.103731f
C1847 por_ana_0.comparator_0.vm avdd 0.390636f
C1848 por_dig_0._033_ por_dig_0.net24 0.530779f
C1849 por_dig_0._043_ dvdd 0.319006f
C1850 por_dig_0.clknet_1_1__leaf_osc_ck a_35583_34541# 1.71964f
C1851 a_34387_32909# dvdd 1.24967f
C1852 a_33804_31251# dvdd 0.444837f
C1853 a_25578_22973# a_26785_22637# 0.28899f
C1854 a_33162_35603# por_dig_0._008_ 0.116176f
C1855 por_ana_0.rstring_mux_0.vtop dvdd 0.152859f
C1856 por_ana_0.rc_osc_0.ena_b por_ana_0.rc_osc_0.vr 0.746068f
C1857 por_ana_0.rc_osc_0.in por_ana_0.rc_osc_0.m 1.10713f
C1858 a_27590_22885# dvdd 0.380879f
C1859 a_40246_23089# avdd 0.184976f
C1860 a_39417_31795# dvdd 0.228729f
C1861 por_dig_0.net19 por_dig_0._035_ 0.241369f
C1862 a_38136_33427# dvdd 0.358791f
C1863 por_dig_0.net22 por_dig_0._036_ 0.201563f
C1864 a_19666_35244# a_20422_35244# 0.296258f
C1865 a_37614_33695# a_37396_33453# 0.209641f
C1866 por_ana_0.rstring_mux_0.otrip_decoded_avdd[2] avdd 1.52796f
C1867 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[0] por_ana_0.rstring_mux_0.vtrip0 0.485675f
C1868 a_34836_30555# dvdd 0.142103f
C1869 a_4433_15512# a_5189_15512# 0.296258f
C1870 a_25578_22973# avdd 0.863791f
C1871 por_dig_0.cnt_st\[0\] por_dig_0._029_ 0.555235f
C1872 a_39887_23089# a_40246_21893# 0.166612f
C1873 a_31412_33427# dvdd 0.372915f
C1874 por_dig_0._034_ por_dig_0.net4 1.03056f
C1875 por_dig_0._036_ a_35000_31795# 0.160002f
C1876 por_dig_0._034_ por_dig_0._037_ 0.346478f
C1877 a_37392_31251# por_dig_0.net34 0.139322f
C1878 a_34615_28013# dvdd 0.198933f
C1879 por_dig_0._035_ por_dig_0.cnt_por\[10\] 0.414793f
C1880 por_ana_0.schmitt_trigger_0.in avss 9.30104f
C1881 por_dig_0.net6 a_35774_28673# 0.107333f
C1882 por_dig_0.cnt_por\[1\] por_dig_0.clknet_1_1__leaf_osc_ck 0.495024f
C1883 por_ana_0.rstring_mux_0.vtrip2 avdd 0.859231f
C1884 a_35500_35629# a_35666_35629# 0.581111f
C1885 por_dig_0.net25 por_dig_0.cnt_por\[9\] 0.201739f
C1886 por_dig_0._025_ dvdd 0.652364f
C1887 por_dig_0.otrip_decoded[4] avdd 0.435076f
C1888 por_dig_0.otrip_decoded[1] avss 0.513938f
C1889 por_dig_0.net24 a_35092_33427# 0.31903f
C1890 por_dig_0.net4 dvdd 3.47243f
C1891 por_dig_0._042_ dvdd 0.899453f
C1892 por_dig_0.net24 a_36016_35629# 0.153351f
C1893 a_38943_23593# a_38518_23637# 0.460766f
C1894 por_dig_0.otrip_decoded[2] porb 0.140184f
C1895 por_dig_0._037_ dvdd 0.561194f
C1896 a_36686_6535# a_37442_6535# 0.296258f
C1897 por_dig_0.cnt_por\[0\] por_dig_0._034_ 0.296287f
C1898 a_4055_22912# avss 0.472952f
C1899 a_34212_30189# dvdd 0.488174f
C1900 a_36328_35091# a_36494_35091# 0.578782f
C1901 por_dig_0.net8 a_31876_32199# 0.159794f
C1902 a_31526_31827# a_32441_32199# 0.125324f
C1903 por_dig_0.net15 otrip[2] 0.228914f
C1904 a_31009_24371# por_ana_0.rstring_mux_0.vtrip_decoded_avdd[1] 0.13699f
C1905 por_dig_0.cnt_por\[4\] por_dig_0.cnt_por\[5\] 0.567854f
C1906 a_34762_36173# dvdd 0.19092f
C1907 por_dig_0.osc_ena por_ana_0.rc_osc_0.in 0.470443f
C1908 a_36138_22973# a_36831_21859# 0.264594f
C1909 a_35224_31277# a_35740_31277# 0.105995f
C1910 por_dig_0.net7 a_36376_28789# 0.207931f
C1911 por_ana_0.vl por_dig_0.otrip_decoded[3] 0.656143f
C1912 a_37064_34003# dvdd 0.511172f
C1913 a_23366_24619# avdd 0.210108f
C1914 a_36308_13935# avss 0.525451f
C1915 a_32019_31643# dvdd 0.206718f
C1916 a_16264_27844# avss 0.460203f
C1917 por_dig_0.clknet_0_osc_ck a_34387_32909# 1.63966f
C1918 por_dig_0.cnt_por\[7\] a_33805_32339# 0.134881f
C1919 a_38150_22885# dvdd 0.38105f
C1920 por_dig_0.cnt_por\[0\] dvdd 2.64246f
C1921 a_37952_31037# a_37777_31111# 0.233657f
C1922 a_38974_34693# dvdd 0.192026f
C1923 a_21944_13935# a_22700_13935# 0.296258f
C1924 por_dig_0.cnt_st\[1\] a_38956_32339# 0.229237f
C1925 por_ana_0.rstring_mux_0.otrip_decoded_avdd[1] por_ana_0.rstring_mux_0.otrip_decoded_avdd[0] 3.24722f
C1926 a_36138_22973# avdd 0.863791f
C1927 a_35699_33819# dvdd 0.212744f
C1928 por_dig_0.otrip_decoded[6] por_dig_0.otrip_decoded[7] 0.78481f
C1929 por_dig_0.clknet_1_0__leaf_osc_ck a_32188_30739# 0.496475f
C1930 por_ana_0.comparator_1.vnn avss 3.09271f
C1931 por_dig_0.net22 por_dig_0._022_ 0.401276f
C1932 a_34467_28557# a_34573_28557# 0.313533f
C1933 a_33155_28640# por_dig_0.net13 0.141743f
C1934 por_dig_0.net24 por_dig_0._024_ 0.133986f
C1935 por_dig_0.clknet_1_1__leaf_osc_ck a_36880_32915# 0.269673f
C1936 avss porb 0.300604f
C1937 avss por 1.09183f
C1938 a_36376_28789# dvdd 0.216714f
C1939 por_ana_0.schmitt_trigger_0.in por_ana_0.rstring_mux_0.otrip_decoded_avdd[5] 0.101776f
C1940 a_31651_30341# por_dig_0.net10 0.14662f
C1941 a_23366_24619# a_23466_24707# 0.40546f
C1942 por_dig_0.otrip_decoded[6] a_27590_22885# 0.276643f
C1943 por_dig_0._011_ a_32651_33819# 0.155634f
C1944 por_dig_0.net3 dvdd 0.408642f
C1945 a_31016_13935# avss 0.465635f
C1946 por_dig_0.cnt_por\[10\] a_35390_31277# 0.559365f
C1947 por_dig_0.clknet_0_osc_ck por_dig_0.net4 0.172949f
C1948 por_ana_0.comparator_1.vnn vbg_1v2 4.4282f
C1949 a_34294_23637# dvdd 0.176078f
C1950 a_34102_29645# dvdd 0.268994f
C1951 por_dig_0.osc_ena por_dig_0.force_pdnb 0.317991f
C1952 por_dig_0._019_ por_dig_0.cnt_por\[4\] 0.199778f
C1953 por_dig_0.clknet_0_osc_ck por_dig_0._037_ 0.10327f
C1954 a_33852_29645# dvdd 0.308935f
C1955 por_ana_0.rc_osc_0.in osc_ck 1.05907f
C1956 por_ana_0.rstring_mux_0.otrip_decoded_avdd[6] por_ana_0.rstring_mux_0.vtrip6 0.489702f
C1957 a_26271_23593# dvdd 0.104499f
C1958 por_dig_0.osc_ena a_19298_6535# 0.209449f
C1959 a_36844_35463# dvdd 0.196229f
C1960 a_6701_15512# avss 0.472978f
C1961 por_dig_0.net25 a_38320_34301# 0.283723f
C1962 por_dig_0._047_ por_dig_0._019_ 0.472259f
C1963 por_ana_0.schmitt_trigger_0.in por_ana_0.rstring_mux_0.otrip_decoded_avdd[2] 0.10426f
C1964 por_dig_0.cnt_por\[0\] por_dig_0.cnt_por\[3\] 0.437419f
C1965 a_38228_30163# a_38053_30189# 0.233657f
C1966 a_30070_23637# avdd 0.142934f
C1967 por_ana_0.comparator_1.vm avss 10.3298f
C1968 a_32740_36179# a_33256_36551# 0.115353f
C1969 a_31394_6535# a_32150_6535# 0.296258f
C1970 por_dig_0.net24 a_32980_33287# 0.217452f
C1971 por_dig_0.net4 por_dig_0.cnt_st\[1\] 0.198454f
C1972 a_31932_31419# a_32088_31514# 0.115353f
C1973 a_31893_31545# a_32019_31643# 0.186387f
C1974 a_34378_30189# a_34728_30189# 0.228712f
C1975 a_33926_24619# avdd 0.206171f
C1976 a_38954_6535# avss 0.730849f
C1977 avss otrip[2] 0.231167f
C1978 a_32358_28013# dvdd 0.181756f
C1979 por_ana_0.rstring_mux_0.otrip_decoded_b_avdd[2] avss 0.363375f
C1980 por_dig_0.net24 dvdd 4.97092f
C1981 a_36138_22973# a_37345_22637# 0.28899f
C1982 por_ana_0.rstring_mux_0.vtrip0 avdd 0.430845f
C1983 a_19094_1626# a_19094_870# 0.296258f
C1984 a_33600_34335# dvdd 0.225172f
C1985 a_24159_21859# dvdd 0.104499f
C1986 por_dig_0._042_ a_37392_31251# 0.177948f
C1987 por_dig_0.cnt_por\[0\] por_dig_0.clknet_0_osc_ck 0.171016f
C1988 por_dig_0.cnt_por\[6\] por_dig_0.cnt_por\[8\] 0.248085f
C1989 a_37156_28013# por_dig_0.otrip_decoded[7] 0.187726f
C1990 por_ana_0.comparator_1.vm vbg_1v2 0.138741f
C1991 a_24212_13935# avss 0.475109f
C1992 por_ana_0.ibias_gen_0.vp1 avss 2.02475f
C1993 a_39888_24823# a_40247_23627# 0.166612f
C1994 por_dig_0.net24 a_35100_32339# 0.340413f
C1995 avss por_timed_out 0.227948f
C1996 a_33474_35059# dvdd 0.21556f
C1997 a_40246_23089# a_40246_21893# 0.136815f
C1998 por_dig_0._031_ a_36382_31795# 0.140129f
C1999 a_16652_13935# a_17408_13935# 0.296258f
C2000 por_dig_0.otrip_decoded[0] a_21254_22885# 0.235746f
C2001 a_25478_24619# a_25846_23637# 0.138963f
C2002 por_dig_0.force_pdnb por_dig_0.otrip_decoded[0] 2.89793f
C2003 a_35612_33595# a_35768_33690# 0.110816f
C2004 a_35573_33721# a_35699_33819# 0.175891f
C2005 a_37800_28013# dvdd 0.306919f
C2006 por_dig_0._041_ por_dig_0._030_ 0.364258f
C2007 a_33805_32339# dvdd 0.183984f
C2008 por_ana_0.rstring_mux_0.vtrip_decoded_b_avdd[1] avss 0.362828f
C2009 por_dig_0.otrip_decoded[3] por_ana_0.rstring_mux_0.otrip_decoded_avdd[1] 0.190261f
C2010 a_21622_21903# dvdd 0.176029f
C2011 por_dig_0.net21 force_short_oneshot 0.203895f
C2012 por_dig_0.clknet_1_0__leaf_osc_ck a_35224_31277# 0.402314f
C2013 a_19298_6535# osc_ck 0.339112f
C2014 por_dig_0.otrip_decoded[7] avdd 0.231113f
C2015 a_33662_6535# avss 0.466333f
C2016 por_dig_0._002_ dvdd 0.787826f
C2017 por_dig_0._003_ a_37138_30189# 0.732617f
C2018 por_dig_0.net23 por_dig_0.net4 1.06665f
C2019 a_25495_33620# dvdd 0.38154f
C2020 por_ana_0.rstring_mux_0.otrip_decoded_b_avdd[6] avdd 0.903548f
C2021 a_34746_31277# dvdd 0.268347f
C2022 a_14374_35244# a_15130_35244# 0.296258f
C2023 a_38943_21859# avdd 0.61228f
C2024 por_dig_0.cnt_st\[2\] dvdd 0.730893f
C2025 por_dig_0._018_ por_dig_0._009_ 0.150079f
C2026 a_31876_32199# dvdd 0.191061f
C2027 a_18920_13935# avss 0.465068f
C2028 a_4811_22912# a_5567_22912# 0.296258f
C2029 por_ana_0.rstring_mux_0.vtop avdd 10.746201f
C2030 a_27590_22885# avdd 0.207177f
C2031 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[1] avss 1.39274f
C2032 por_ana_0.sky130_fd_sc_hvl__inv_1_0.A dvdd 0.11431f
C2033 a_31893_33721# dvdd 0.589314f
C2034 a_35674_28557# a_35774_28673# 0.167615f
C2035 por_ana_0.rstring_mux_0.otrip_decoded_avdd[0] por_ana_0.rstring_mux_0.otrip_decoded_b_avdd[0] 0.56463f
C2036 por_dig_0._051_ dvdd 1.63412f
C2037 a_35111_28013# dvdd 0.20791f
C2038 por_ana_0.ibias_gen_0.vp1 ibg_200n 0.181982f
C2039 por_ana_0.rstring_mux_0.ena_b avss 1.61845f
C2040 a_37046_32915# a_37396_33287# 0.219633f
C2041 por_dig_0.net5 a_32358_28013# 0.371583f
C2042 force_short_oneshot startup_timed_out 0.206128f
C2043 dvdd vin 0.329013f
C2044 por_dig_0.cnt_por\[1\] por_dig_0._016_ 0.103972f
C2045 por_dig_0.net24 por_dig_0.clknet_0_osc_ck 0.170156f
C2046 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[4] dvdd 0.669746f
C2047 por_dig_0._042_ a_39510_31251# 0.122663f
C2048 a_35500_35629# a_36016_35629# 0.110816f
C2049 por_ana_0.rstring_mux_0.vtrip_decoded_b_avdd[5] avdd 0.90363f
C2050 por_dig_0.net23 por_dig_0.cnt_por\[0\] 1.20897f
C2051 a_24590_6535# a_25346_6535# 0.296258f
C2052 por_ana_0.rstring_mux_0.otrip_decoded_avdd[6] avss 1.36421f
C2053 por_dig_0.cnt_por\[2\] a_34580_35629# 0.112499f
C2054 a_26288_32594# a_25863_32638# 0.460766f
C2055 por_dig_0.cnt_por\[1\] a_36494_35091# 0.589783f
C2056 por_dig_0.net24 a_36581_35629# 0.235709f
C2057 a_37064_13935# a_37820_13935# 0.296258f
C2058 dvdd force_pdn 1.00084f
C2059 por_dig_0.cnt_st\[4\] por_dig_0._032_ 0.514901f
C2060 por_ana_0.rstring_mux_0.otrip_decoded_avdd[3] dvdd 0.375895f
C2061 por_dig_0.cnt_por\[2\] por_dig_0._052_ 0.307908f
C2062 a_17020_27844# a_17776_27844# 0.296258f
C2063 a_33806_33427# dvdd 0.215539f
C2064 a_38250_24707# a_38943_23593# 0.264594f
C2065 a_36494_35091# a_37062_35059# 0.175891f
C2066 a_36328_35091# a_36844_35463# 0.106087f
C2067 por_dig_0.net8 a_32441_32199# 0.237171f
C2068 por_ana_0.rstring_mux_0.otrip_decoded_avdd[2] por_ana_0.rstring_mux_0.otrip_decoded_b_avdd[2] 0.572197f
C2069 por_dig_0.cnt_por\[5\] por_dig_0.cnt_por\[8\] 0.193923f
C2070 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[4] por_ana_0.dcomp3v3uv 0.249577f
C2071 a_13628_13935# avss 0.465267f
C2072 por_dig_0.osc_ena por_ana_0.rc_osc_0.m 0.255672f
C2073 por_dig_0._006_ dvdd 0.449926f
C2074 a_32354_30739# dvdd 0.57524f
C2075 a_33926_24619# a_34026_24707# 0.40546f
C2076 a_35224_31277# a_36305_31277# 0.102355f
C2077 por_ana_0.comparator_1.vn avdd 0.721561f
C2078 a_24673_24371# avdd 0.420074f
C2079 por_dig_0.net25 a_36880_33453# 0.301808f
C2080 por_dig_0.net4 por_dig_0.net22 0.993695f
C2081 por_ana_0.rstring_mux_0.otrip_decoded_avdd[1] por_ana_0.rstring_mux_0.otrip_decoded_b_avdd[1] 0.569059f
C2082 por_dig_0.cnt_st\[4\] a_38500_31251# 0.310614f
C2083 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[3] por_ana_0.rstring_mux_0.vtrip_decoded_avdd[4] 1.04751f
C2084 por_ana_0.rstring_mux_0.otrip_decoded_avdd[3] por_ana_0.dcomp3v3uv 0.156703f
C2085 por_dig_0.net24 a_36328_35091# 0.402642f
C2086 por_ana_0.rstring_mux_0.otrip_decoded_b_avdd[2] por_ana_0.rstring_mux_0.vtrip2 0.190544f
C2087 a_39328_34515# dvdd 0.32722f
C2088 por_dig_0._010_ a_32464_32915# 0.231092f
C2089 por_dig_0.otrip_decoded[4] otrip[2] 0.619319f
C2090 por_dig_0._047_ por_dig_0._020_ 0.405285f
C2091 por_dig_0.net16 por_dig_0.net18 0.167027f
C2092 a_21566_6535# avss 0.466333f
C2093 a_38150_22885# avdd 0.207184f
C2094 por_dig_0._022_ a_34212_33997# 0.100412f
C2095 por_ana_0.vl isrc_sel 1.09217f
C2096 por_ana_0.rstring_mux_0.otrip_decoded_b_avdd[3] vin 0.340862f
C2097 por_dig_0.cnt_por\[7\] por_dig_0.cnt_por\[9\] 0.21587f
C2098 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[0] vin 0.252789f
C2099 a_32906_36179# a_33474_36147# 0.180982f
C2100 por_dig_0.cnt_st\[1\] por_dig_0.cnt_st\[2\] 0.311814f
C2101 por_dig_0.net23 por_dig_0.net24 0.133472f
C2102 a_23466_24707# a_24673_24371# 0.28899f
C2103 por_ana_0.rstring_mux_0.otrip_decoded_avdd[3] por_ana_0.rstring_mux_0.otrip_decoded_b_avdd[3] 0.571961f
C2104 por_ana_0.rstring_mux_0.otrip_decoded_avdd[3] por_ana_0.sky130_fd_sc_hvl__lsbufhv2lv_1_1.X 1.37931f
C2105 por_dig_0._033_ por_dig_0.net20 0.477793f
C2106 por_ana_0.rstring_mux_0.otrip_decoded_avdd[5] por_ana_0.rstring_mux_0.otrip_decoded_avdd[6] 0.340239f
C2107 por_dig_0._047_ a_33162_35603# 0.194921f
C2108 a_34746_29645# dvdd 0.253454f
C2109 a_36406_23637# dvdd 0.172761f
C2110 a_35202_29877# dvdd 0.178763f
C2111 por_dig_0._052_ por_dig_0._047_ 0.163106f
C2112 por_ana_0.rc_osc_0.m osc_ck 1.09311f
C2113 por_dig_0.clknet_1_1__leaf_osc_ck a_31932_33595# 0.444807f
C2114 a_37409_35463# dvdd 0.299783f
C2115 por_dig_0._043_ a_39497_30849# 0.107389f
C2116 a_19298_6535# a_20054_6535# 0.296258f
C2117 por_dig_0._039_ por_dig_0.net21 0.183141f
C2118 por_dig_0.net24 a_32244_32365# 0.153457f
C2119 a_36138_24707# dvdd 0.243001f
C2120 a_16274_6535# avss 0.466333f
C2121 a_34294_23637# avdd 0.142934f
C2122 a_35500_35629# dvdd 0.442291f
C2123 a_32740_36179# a_33821_36551# 0.102325f
C2124 a_31772_13935# a_32528_13935# 0.296258f
C2125 a_35640_32517# dvdd 0.178477f
C2126 a_26271_23593# avdd 0.607928f
C2127 a_32740_35091# a_32906_35091# 0.906454f
C2128 por_dig_0.net24 a_33545_33287# 0.271215f
C2129 a_32088_31514# a_32019_31643# 0.209641f
C2130 a_34378_30189# a_35293_30189# 0.118759f
C2131 a_35233_24371# avdd 0.420074f
C2132 a_32641_28013# dvdd 0.178716f
C2133 a_19666_35244# avss 0.460203f
C2134 por_dig_0.cnt_por\[4\] por_dig_0._035_ 0.167587f
C2135 avss itest 3.62448f
C2136 por_dig_0._015_ dvdd 0.479362f
C2137 por_dig_0._013_ a_32609_31099# 0.170087f
C2138 por_dig_0._028_ dvdd 0.495212f
C2139 por_dig_0.net25 a_34728_30189# 0.153286f
C2140 por_ana_0.rstring_mux_0.otrip_decoded_avdd[0] avss 1.64125f
C2141 a_32984_32339# a_32809_32365# 0.233657f
C2142 por_ana_0.vl por_dig_0.por_unbuf 0.129633f
C2143 a_7457_15512# a_8213_15512# 0.296258f
C2144 por_dig_0.net24 por_dig_0._013_ 0.113983f
C2145 a_24159_21859# avdd 0.607928f
C2146 por_dig_0.net19 a_31728_32365# 0.222506f
C2147 por_dig_0.net19 a_31592_30965# 0.135905f
C2148 a_37596_30555# dvdd 0.132556f
C2149 por_dig_0.net30 a_35202_29877# 0.135907f
C2150 a_33996_35389# dvdd 0.371682f
C2151 por_dig_0._017_ por_dig_0.net19 0.113322f
C2152 por_dig_0.net27 a_35224_31277# 0.296022f
C2153 vbg_1v2 itest 0.152663f
C2154 a_35768_33690# a_35699_33819# 0.209641f
C2155 por_dig_0.net4 a_39497_30849# 0.135147f
C2156 por_dig_0.net7 a_35776_28013# 0.168145f
C2157 por_dig_0.osc_ena por_dig_0.otrip_decoded[0] 3.95147f
C2158 por_dig_0.cnt_st\[2\] a_38352_32365# 0.200444f
C2159 por_dig_0._026_ dvdd 0.360588f
C2160 por_dig_0.net24 por_dig_0.net22 0.203362f
C2161 por_dig_0.net22 a_33600_34335# 0.191752f
C2162 a_31413_32339# dvdd 0.255122f
C2163 a_25478_22885# a_25846_21903# 0.138963f
C2164 a_33121_22637# por_ana_0.rstring_mux_0.vtrip_decoded_avdd[2] 0.135857f
C2165 por_dig_0._050_ dvdd 0.594161f
C2166 a_25846_21903# dvdd 0.176016f
C2167 por_dig_0.osc_ena osc_ck 4.63024f
C2168 por_dig_0.net11 a_35960_29101# 0.125932f
C2169 por_dig_0._006_ a_36328_35091# 0.216312f
C2170 por_dig_0.cnt_por\[0\] por_dig_0.cnt_por\[1\] 1.95704f
C2171 por_dig_0.net1 por_dig_0.cnt_rsb_stg1 0.629951f
C2172 por_dig_0.net6 por_dig_0.net11 0.252295f
C2173 por_dig_0._049_ dvdd 0.239638f
C2174 a_27590_22885# a_27690_22973# 0.40546f
C2175 por_dig_0._015_ por_dig_0.net30 0.240262f
C2176 por_dig_0.net28 a_31526_31827# 0.54292f
C2177 por_dig_0.otrip_decoded[2] por_dig_0.otrip_decoded[3] 0.316118f
C2178 a_21622_21903# avdd 0.143941f
C2179 a_38136_33427# a_37961_33453# 0.233657f
C2180 por_dig_0.cnt_por\[9\] dvdd 1.93742f
C2181 por_ana_0.comparator_1.ena_b avdd 0.998725f
C2182 a_32441_32199# dvdd 0.29735f
C2183 a_25495_33620# avdd 0.191575f
C2184 a_28897_22637# avdd 0.421965f
C2185 force_dis_rc_osc force_pdn 0.319714f
C2186 por_dig_0.cnt_por\[10\] por_dig_0.cnt_por\[8\] 0.119476f
C2187 a_39077_31527# por_dig_0._003_ 0.106913f
C2188 a_32088_33690# dvdd 0.196979f
C2189 por_dig_0.net27 a_34852_31277# 0.130538f
C2190 por_dig_0.net4 por_dig_0.cnt_st\[3\] 0.847277f
C2191 por_dig_0._022_ por_dig_0._023_ 0.244938f
C2192 por_dig_0.clknet_1_0__leaf_osc_ck por_dig_0.net19 0.325148f
C2193 a_32828_35879# dvdd 0.194001f
C2194 por_dig_0.cnt_por\[6\] por_dig_0._022_ 0.379825f
C2195 por_dig_0.cnt_st\[3\] por_dig_0._042_ 0.463837f
C2196 a_35776_28013# dvdd 0.252579f
C2197 a_36122_30341# por_dig_0.net29 0.131599f
C2198 a_14006_6535# a_14762_6535# 0.296258f
C2199 otrip[1] otrip[0] 3.57166f
C2200 a_26785_24371# por_ana_0.rstring_mux_0.otrip_decoded_avdd[5] 0.13699f
C2201 a_37046_32915# a_37961_33287# 0.125324f
C2202 por_dig_0.net6 por_dig_0.net14 0.103373f
C2203 a_31360_28557# por_dig_0.net3 0.134646f
C2204 por_ana_0.sky130_fd_sc_hvl__inv_1_0.A avdd 0.728126f
C2205 a_31412_33427# a_31615_33705# 0.233657f
C2206 a_37751_31251# dvdd 0.193476f
C2207 a_35500_35629# a_36581_35629# 0.102325f
C2208 a_24968_13935# a_25724_13935# 0.296258f
C2209 a_13844_23626# ibg_200n 0.398549f
C2210 por_dig_0.net24 a_35768_33690# 0.153794f
C2211 por_dig_0.otrip_decoded[7] otrip[2] 0.162044f
C2212 por_dig_0.force_pdnb otrip[0] 0.174496f
C2213 avdd vin 8.665781f
C2214 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[4] avdd 1.61396f
C2215 a_39888_24823# dvdd 0.13819f
C2216 a_35913_33819# dvdd 0.142103f
C2217 por_dig_0.clknet_1_1__leaf_osc_ck por_dig_0._005_ 0.29702f
C2218 a_4811_22912# avss 0.471605f
C2219 a_17398_35244# a_18154_35244# 0.296258f
C2220 por_ana_0.dcomp3v3 dvdd 1.17353f
C2221 a_33971_28557# otrip[1] 0.261941f
C2222 a_27590_24619# dvdd 0.387197f
C2223 por_dig_0.net20 por_dig_0._034_ 0.503575f
C2224 a_36328_35091# a_37409_35463# 0.102355f
C2225 a_37062_35059# a_36844_35463# 0.209641f
C2226 a_2165_15512# a_2921_15512# 0.296258f
C2227 por_dig_0.net25 a_35958_31519# 0.159426f
C2228 avdd force_pdn 0.222115f
C2229 por_ana_0.rc_osc_0.in dvdd 5.41497f
C2230 a_38250_22973# a_38943_21859# 0.264594f
C2231 a_34026_24707# a_35233_24371# 0.28899f
C2232 por_ana_0.rstring_mux_0.otrip_decoded_avdd[3] avdd 1.72013f
C2233 por_dig_0.net6 a_33172_28165# 0.165328f
C2234 a_32704_31111# dvdd 0.198277f
C2235 por_dig_0.net8 a_32004_30189# 0.123008f
C2236 por_dig_0.cnt_por\[1\] por_dig_0.net24 1.56558f
C2237 por_dig_0._005_ a_35704_35124# 0.124183f
C2238 por_ana_0.comparator_1.n0 avdd 0.966571f
C2239 por_ana_0.comparator_1.vnn por_ana_0.comparator_1.vn 0.290508f
C2240 por_dig_0._033_ por_dig_0._018_ 0.144204f
C2241 a_25578_24707# avdd 0.863296f
C2242 a_35848_31643# dvdd 0.142416f
C2243 a_33996_36477# dvdd 0.415564f
C2244 a_37064_13935# avss 0.525451f
C2245 por_dig_0.net4 por_dig_0._030_ 0.145576f
C2246 a_17020_27844# avss 0.460203f
C2247 por_dig_0.cnt_por\[4\] por_dig_0.net32 0.148219f
C2248 por_dig_0._030_ por_dig_0._042_ 0.189781f
C2249 por_dig_0.net24 a_37062_35059# 0.176368f
C2250 por_dig_0._013_ a_32354_30739# 0.737247f
C2251 por_dig_0.net20 dvdd 2.13581f
C2252 a_34615_28013# otrip[2] 0.259384f
C2253 por_dig_0.net25 a_36696_30739# 0.342123f
C2254 a_39457_22637# avdd 0.420442f
C2255 por_ana_0.sky130_fd_sc_hvl__inv_1_0.A por_ana_0.sky130_fd_sc_hvl__inv_4_0.A 0.166308f
C2256 a_34418_6535# a_35174_6535# 0.296258f
C2257 a_14374_35244# avss 0.743991f
C2258 por_dig_0.net23 a_35640_32517# 0.249334f
C2259 a_31914_24707# a_32607_23593# 0.264594f
C2260 a_33474_36147# por_dig_0.net24 0.170427f
C2261 por_dig_0.net1 por_dig_0.net19 0.231828f
C2262 por_dig_0.force_pdnb por_dig_0.otrip_decoded[5] 0.103672f
C2263 por_dig_0.net5 a_35776_28013# 0.249451f
C2264 a_27690_24707# a_28383_23593# 0.264594f
C2265 dvdd otrip[1] 0.790889f
C2266 dvdd dcomp 2.40097f
C2267 por_ana_0.comparator_1.vn por_ana_0.comparator_1.vm 4.6608f
C2268 a_33364_36173# dvdd 0.137085f
C2269 a_38320_34301# dvdd 0.360195f
C2270 a_34212_30189# por_dig_0._014_ 0.166346f
C2271 por_dig_0.net25 a_36972_30189# 0.386941f
C2272 a_31772_13935# avss 0.465592f
C2273 por_dig_0.force_pdnb dvdd 1.15218f
C2274 a_21254_22885# dvdd 0.382499f
C2275 a_35556_29619# dvdd 0.326413f
C2276 a_7457_15512# avss 0.472978f
C2277 a_19676_13935# a_20432_13935# 0.296258f
C2278 por_ana_0.rstring_mux_0.vtrip6 a_29126_6535# 0.298448f
C2279 a_24159_23593# a_23734_23637# 0.460766f
C2280 a_38150_24619# dvdd 0.441504f
C2281 por_dig_0.net24 a_32809_32365# 0.258141f
C2282 a_34378_30189# dvdd 0.536464f
C2283 por_ana_0.rstring_mux_0.otrip_decoded_avdd[6] por_ana_0.rstring_mux_0.otrip_decoded_b_avdd[6] 0.573474f
C2284 a_36406_23637# avdd 0.142934f
C2285 por_dig_0.cnt_por\[1\] por_dig_0._051_ 0.23013f
C2286 a_37064_34003# por_dig_0._000_ 0.617523f
C2287 por_ana_0.rstring_mux_0.ena_b por_ana_0.rstring_mux_0.vtop 2.52783f
C2288 por_dig_0.net20 por_dig_0.cnt_por\[3\] 0.147803f
C2289 a_36564_32339# dvdd 0.237515f
C2290 a_32740_35091# a_33256_35463# 0.115353f
C2291 a_32906_35091# a_33474_35059# 0.186387f
C2292 a_37392_31251# a_37751_31251# 0.141213f
C2293 por_dig_0._034_ a_36382_31795# 0.141269f
C2294 por_dig_0.net24 a_36880_32915# 0.662434f
C2295 a_35390_31277# a_35740_31277# 0.219633f
C2296 a_36138_24707# avdd 0.863296f
C2297 por_dig_0._035_ por_dig_0.cnt_por\[8\] 0.267127f
C2298 a_37230_34003# dvdd 0.600481f
C2299 a_38150_22885# a_38250_22973# 0.40546f
C2300 por_ana_0.rstring_mux_0.otrip_decoded_b_avdd[1] avss 0.365652f
C2301 por_dig_0.force_pdnb por_ana_0.dcomp3v3uv 0.103342f
C2302 por_dig_0.net23 por_dig_0._049_ 0.107472f
C2303 a_14374_35244# ibg_200n 0.253354f
C2304 por_dig_0.net25 a_35293_30189# 0.242247f
C2305 a_31360_28557# force_pdn 0.20079f
C2306 a_38974_34693# a_39070_34515# 0.419086f
C2307 a_24968_13935# avss 0.482553f
C2308 a_7835_22912# a_8591_22912# 0.296258f
C2309 por_dig_0.net24 a_31615_33705# 0.22274f
C2310 a_36382_31795# dvdd 0.607023f
C2311 dvdd force_short_oneshot 0.700383f
C2312 por_dig_0.cnt_por\[6\] a_31412_33427# 0.128929f
C2313 a_31413_29619# por_dig_0.osc_ena 0.156202f
C2314 a_34672_35451# dvdd 0.394835f
C2315 por_ana_0.rstring_mux_0.vtop a_13628_13935# 0.348335f
C2316 por_ana_0.schmitt_trigger_0.in por_ana_0.rstring_mux_0.vtrip_decoded_avdd[4] 0.158489f
C2317 por_dig_0._013_ por_dig_0._028_ 0.203345f
C2318 a_2165_15512# avss 0.761384f
C2319 a_27590_24619# a_27958_23637# 0.138963f
C2320 por_dig_0._014_ a_33852_29645# 0.173603f
C2321 isrc_sel dvss 3.56289f
C2322 otrip[2] dvss 3.80763f
C2323 otrip[0] dvss 3.465244f
C2324 otrip[1] dvss 3.349186f
C2325 porb dvss 6.254727f
C2326 pwup_filt dvss 9.044774f
C2327 dcomp dvss 4.621289f
C2328 por dvss 3.872764f
C2329 ibg_200n dvss 5.74584f
C2330 startup_timed_out dvss 1.99626f
C2331 force_short_oneshot dvss 4.52209f
C2332 por_timed_out dvss 3.41504f
C2333 osc_ck dvss 19.978914f
C2334 force_pdn dvss 4.168776f
C2335 force_dis_rc_osc dvss 4.305812f
C2336 force_ena_rc_osc dvss 4.143809f
C2337 itest dvss 7.16946f
C2338 vbg_1v2 dvss 51.201763f
C2339 porb_h dvss -0.231006f
C2340 vin dvss 26.508797f
C2341 dvdd dvss 1.468185p
C2342 avss dvss 0.293557p
C2343 avdd dvss 3.758295p
C2344 a_41694_492# dvss 1.27808f
C2345 a_19094_870# dvss 1.12408f
C2346 a_41694_1248# dvss 0.990226f
C2347 a_19094_1626# dvss 1.1316f
C2348 a_41694_2004# dvss 0.990193f
C2349 a_19094_2382# dvss 1.30717f
C2350 a_41694_2760# dvss 0.996823f
C2351 a_19094_3138# dvss 1.18151f
C2352 a_41694_3516# dvss 1.30652f
C2353 por_ana_0.rc_osc_0.vr dvss 3.37131f
C2354 por_ana_0.rc_osc_0.m dvss 3.35105f
C2355 por_ana_0.rc_osc_0.in dvss 0.433849p
C2356 por_ana_0.rc_osc_0.ena_b dvss 1.37315f
C2357 a_38954_6535# dvss 0.612822f
C2358 a_38576_13935# dvss 0.659772f
C2359 a_38198_6535# dvss 0.61321f
C2360 a_37820_13935# dvss 0.659772f
C2361 a_37442_6535# dvss 0.61321f
C2362 a_37064_13935# dvss 0.659772f
C2363 a_36686_6535# dvss 0.61321f
C2364 a_36308_13935# dvss 0.659772f
C2365 a_35930_6535# dvss 0.61321f
C2366 a_35552_13935# dvss 0.659772f
C2367 a_35174_6535# dvss 0.61321f
C2368 a_34796_13935# dvss 0.659772f
C2369 a_34418_6535# dvss 0.618291f
C2370 a_34040_13935# dvss 0.659772f
C2371 a_33662_6535# dvss 0.61321f
C2372 a_33284_13935# dvss 0.647659f
C2373 a_32906_6535# dvss 0.61321f
C2374 a_32528_13935# dvss 0.653638f
C2375 a_32150_6535# dvss 0.61321f
C2376 a_31772_13935# dvss 0.656775f
C2377 a_31394_6535# dvss 0.61321f
C2378 a_31016_13935# dvss 0.656775f
C2379 a_30638_6535# dvss 0.61321f
C2380 a_30260_13935# dvss 0.656775f
C2381 a_29882_6535# dvss 0.61321f
C2382 a_29504_13935# dvss 0.642157f
C2383 a_29126_6535# dvss 0.61321f
C2384 a_25724_13935# dvss 0.635008f
C2385 a_25346_6535# dvss 0.61321f
C2386 a_24968_13935# dvss 0.640419f
C2387 a_24590_6535# dvss 0.61321f
C2388 a_24212_13935# dvss 0.643911f
C2389 a_23834_6535# dvss 0.61321f
C2390 a_23456_13935# dvss 0.643911f
C2391 a_23078_6535# dvss 0.61321f
C2392 a_22700_13935# dvss 0.643911f
C2393 a_22322_6535# dvss 0.61321f
C2394 a_21944_13935# dvss 0.645008f
C2395 a_21566_6535# dvss 0.621617f
C2396 a_21188_13935# dvss 0.651324f
C2397 a_20810_6535# dvss 0.644889f
C2398 a_20432_13935# dvss 1.03302f
C2399 a_20054_6535# dvss 0.908892f
C2400 a_19676_13935# dvss 0.592431f
C2401 a_19298_6535# dvss 0.594185f
C2402 a_18920_13935# dvss 0.642912f
C2403 a_18542_6535# dvss 0.61321f
C2404 a_18164_13935# dvss 0.643911f
C2405 a_17786_6535# dvss 0.61321f
C2406 a_17408_13935# dvss 0.643911f
C2407 a_17030_6535# dvss 0.61321f
C2408 a_16652_13935# dvss 0.643911f
C2409 a_16274_6535# dvss 0.61321f
C2410 a_15896_13935# dvss 0.643911f
C2411 a_15518_6535# dvss 0.612139f
C2412 a_15140_13935# dvss 0.643911f
C2413 a_14762_6535# dvss 0.615216f
C2414 a_14384_13935# dvss 0.643911f
C2415 a_14006_6535# dvss 0.61321f
C2416 a_13628_13935# dvss 0.628722f
C2417 a_13250_6535# dvss 0.612803f
C2418 por_ana_0.comparator_0.n0 dvss 5.074068f
C2419 por_ana_0.comparator_0.vm dvss 9.48255f
C2420 por_ana_0.comparator_0.vn dvss 5.932258f
C2421 por_ana_0.comparator_0.vnn dvss 47.770573f
C2422 por_ana_0.rstring_mux_0.vtrip6 dvss 6.67504f
C2423 por_ana_0.rstring_mux_0.vtrip4 dvss 5.681643f
C2424 por_ana_0.rstring_mux_0.vtrip2 dvss 5.372343f
C2425 por_ana_0.rstring_mux_0.vtrip0 dvss 6.512494f
C2426 por_ana_0.rstring_mux_0.vtop dvss 16.1712f
C2427 por_ana_0.rstring_mux_0.ena_b dvss 2.14242f
C2428 por_ana_0.rstring_mux_0.vtrip_decoded_b_avdd[7] dvss 0.214336f
C2429 por_ana_0.rstring_mux_0.vtrip_decoded_b_avdd[6] dvss 0.191802f
C2430 por_ana_0.rstring_mux_0.vtrip_decoded_b_avdd[5] dvss 0.191802f
C2431 por_ana_0.rstring_mux_0.vtrip_decoded_b_avdd[4] dvss 0.191802f
C2432 por_ana_0.rstring_mux_0.vtrip_decoded_b_avdd[3] dvss 0.191802f
C2433 por_ana_0.rstring_mux_0.vtrip_decoded_b_avdd[2] dvss 0.191802f
C2434 por_ana_0.rstring_mux_0.vtrip_decoded_b_avdd[1] dvss 0.191801f
C2435 por_ana_0.rstring_mux_0.vtrip_decoded_b_avdd[0] dvss 0.193218f
C2436 por_ana_0.rstring_mux_0.otrip_decoded_b_avdd[7] dvss 0.191802f
C2437 por_ana_0.rstring_mux_0.otrip_decoded_b_avdd[6] dvss 0.191802f
C2438 por_ana_0.rstring_mux_0.otrip_decoded_b_avdd[5] dvss 0.191802f
C2439 por_ana_0.rstring_mux_0.otrip_decoded_b_avdd[4] dvss 0.191802f
C2440 por_ana_0.rstring_mux_0.otrip_decoded_b_avdd[3] dvss 0.181122f
C2441 por_ana_0.rstring_mux_0.otrip_decoded_b_avdd[2] dvss 0.191802f
C2442 por_ana_0.rstring_mux_0.otrip_decoded_b_avdd[1] dvss 0.191802f
C2443 por_ana_0.rstring_mux_0.otrip_decoded_b_avdd[0] dvss 0.195093f
C2444 por_ana_0.sky130_fd_sc_hvl__lsbufhv2lv_1_1.X dvss 2.76911f
C2445 a_38518_21903# dvss 1.70784f
C2446 a_36406_21903# dvss 1.72434f
C2447 a_39887_21959# dvss 0.901636f
C2448 a_34294_21903# dvss 1.72666f
C2449 a_32182_21903# dvss 1.72672f
C2450 a_30070_21903# dvss 1.72474f
C2451 a_27958_21903# dvss 1.71031f
C2452 a_25846_21903# dvss 1.70837f
C2453 a_23734_21903# dvss 1.70837f
C2454 a_21622_21903# dvss 1.70965f
C2455 a_40246_21893# dvss 1.01257f
C2456 a_38943_21859# dvss 0.849946f
C2457 a_36831_21859# dvss 0.870955f
C2458 a_40246_23089# dvss 0.860748f
C2459 por_ana_0.dcomp3v3uv dvss 7.57486f
C2460 a_39887_23089# dvss 1.27483f
C2461 a_34719_21859# dvss 0.876718f
C2462 a_32607_21859# dvss 0.876774f
C2463 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[4] dvss 2.471994f
C2464 a_30495_21859# dvss 0.875757f
C2465 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[2] dvss 1.71779f
C2466 a_28383_21859# dvss 0.873335f
C2467 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[0] dvss 1.50396f
C2468 a_26271_21859# dvss 0.867563f
C2469 por_ana_0.rstring_mux_0.otrip_decoded_avdd[6] dvss 1.21873f
C2470 a_24159_21859# dvss 0.867563f
C2471 por_ana_0.rstring_mux_0.otrip_decoded_avdd[4] dvss 1.03707f
C2472 a_22047_21859# dvss 0.867659f
C2473 por_ana_0.rstring_mux_0.otrip_decoded_avdd[2] dvss 1.39669f
C2474 por_ana_0.rstring_mux_0.otrip_decoded_avdd[0] dvss 1.07955f
C2475 a_39457_22637# dvss 0.492237f
C2476 a_38250_22973# dvss 1.52132f
C2477 a_38150_22885# dvss 1.97869f
C2478 a_37345_22637# dvss 0.503164f
C2479 a_36138_22973# dvss 1.52795f
C2480 a_36038_22885# dvss 2.199f
C2481 a_35233_22637# dvss 0.503164f
C2482 a_34026_22973# dvss 1.52792f
C2483 a_33926_22885# dvss 2.19988f
C2484 a_33121_22637# dvss 0.503164f
C2485 a_31914_22973# dvss 1.52796f
C2486 a_31814_22885# dvss 2.19989f
C2487 a_31009_22637# dvss 0.503164f
C2488 a_29802_22973# dvss 1.52795f
C2489 a_29702_22885# dvss 2.19989f
C2490 a_28897_22637# dvss 0.503164f
C2491 a_27690_22973# dvss 1.52227f
C2492 a_27590_22885# dvss 1.97975f
C2493 a_26785_22637# dvss 0.503164f
C2494 a_25578_22973# dvss 1.52226f
C2495 a_25478_22885# dvss 1.97975f
C2496 a_24673_22637# dvss 0.503164f
C2497 a_23466_22973# dvss 1.52226f
C2498 a_23366_22885# dvss 1.97975f
C2499 a_22561_22637# dvss 0.503164f
C2500 a_21354_22973# dvss 1.52865f
C2501 a_21254_22885# dvss 2.03022f
C2502 a_38518_23637# dvss 1.69131f
C2503 a_36406_23637# dvss 1.70825f
C2504 a_39888_23693# dvss 0.891927f
C2505 a_34294_23637# dvss 1.71064f
C2506 a_32182_23637# dvss 1.70983f
C2507 a_30070_23637# dvss 1.70983f
C2508 a_27958_23637# dvss 1.69341f
C2509 a_25846_23637# dvss 1.69148f
C2510 a_23734_23637# dvss 1.69215f
C2511 a_21622_23637# dvss 1.69266f
C2512 a_40247_23627# dvss 1.00552f
C2513 a_38943_23593# dvss 0.85f
C2514 a_36831_23593# dvss 0.871007f
C2515 a_40247_24823# dvss 0.865908f
C2516 a_39888_24823# dvss 1.28707f
C2517 a_34719_23593# dvss 0.87832f
C2518 a_32607_23593# dvss 0.876774f
C2519 a_30495_23593# dvss 0.876774f
C2520 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[3] dvss 2.08084f
C2521 a_28383_23593# dvss 0.873329f
C2522 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[1] dvss 2.16902f
C2523 a_26271_23593# dvss 0.867563f
C2524 por_ana_0.rstring_mux_0.otrip_decoded_avdd[7] dvss 1.87055f
C2525 a_24159_23593# dvss 0.867974f
C2526 por_ana_0.rstring_mux_0.otrip_decoded_avdd[5] dvss 1.73534f
C2527 a_22047_23593# dvss 0.867659f
C2528 por_ana_0.rstring_mux_0.otrip_decoded_avdd[3] dvss 1.52516f
C2529 por_ana_0.rstring_mux_0.otrip_decoded_avdd[1] dvss 1.64366f
C2530 a_39457_24371# dvss 0.495673f
C2531 a_38250_24707# dvss 1.53892f
C2532 a_38150_24619# dvss 1.99086f
C2533 a_37345_24371# dvss 0.506586f
C2534 a_36138_24707# dvss 1.543f
C2535 a_36038_24619# dvss 2.2054f
C2536 a_35233_24371# dvss 0.506586f
C2537 a_34026_24707# dvss 1.5398f
C2538 a_33926_24619# dvss 2.18683f
C2539 a_33121_24371# dvss 0.501383f
C2540 a_31914_24707# dvss 1.53264f
C2541 a_31814_24619# dvss 2.18683f
C2542 a_31009_24371# dvss 0.501383f
C2543 a_29802_24707# dvss 1.53264f
C2544 a_29702_24619# dvss 2.18683f
C2545 a_28897_24371# dvss 0.501383f
C2546 a_27690_24707# dvss 1.52954f
C2547 a_27590_24619# dvss 1.96643f
C2548 a_26785_24371# dvss 0.500163f
C2549 a_25578_24707# dvss 1.52683f
C2550 a_25478_24619# dvss 1.96734f
C2551 a_24673_24371# dvss 0.512534f
C2552 a_23466_24707# dvss 1.53695f
C2553 a_23366_24619# dvss 1.97338f
C2554 a_22561_24371# dvss 0.501043f
C2555 a_21354_24707# dvss 1.53541f
C2556 a_21254_24619# dvss 2.02178f
C2557 por_dig_0.otrip_decoded[0] dvss 4.302717f
C2558 a_38444_28013# dvss 0.3838f
C2559 por_dig_0.otrip_decoded[3] dvss 3.291277f
C2560 a_37800_28013# dvss 0.37203f
C2561 por_dig_0.otrip_decoded[7] dvss 2.997841f
C2562 a_37156_28013# dvss 0.387358f
C2563 por_dig_0.otrip_decoded[5] dvss 3.351318f
C2564 a_36512_28013# dvss 0.343397f
C2565 por_dig_0.net18 dvss 0.621031f
C2566 a_35394_28013# dvss 0.164915f
C2567 a_35776_28013# dvss 0.274615f
C2568 a_35217_28013# dvss 0.24219f
C2569 a_35111_28013# dvss 0.232859f
C2570 a_34934_28013# dvss 0.268731f
C2571 a_34615_28013# dvss 0.241123f
C2572 por_dig_0.otrip_decoded[4] dvss 3.56096f
C2573 por_dig_0.otrip_decoded[2] dvss 4.793302f
C2574 a_34265_27987# dvss 0.30886f
C2575 a_33752_28013# dvss 0.34545f
C2576 a_33172_28165# dvss 0.231975f
C2577 a_32641_28013# dvss 0.23192f
C2578 a_32535_28013# dvss 0.222239f
C2579 a_32358_28013# dvss 0.22677f
C2580 a_32039_28013# dvss 0.296078f
C2581 a_36649_28789# dvss 0.201035f
C2582 por_dig_0.net16 dvss 0.337342f
C2583 por_dig_0.net14 dvss 1.59787f
C2584 a_36376_28789# dvss 0.228014f
C2585 a_35774_28673# dvss 0.230016f
C2586 a_35674_28557# dvss 0.19951f
C2587 a_35130_28673# dvss 0.244253f
C2588 a_35030_28557# dvss 0.231636f
C2589 a_34750_28557# dvss 0.100256f
C2590 por_dig_0.net13 dvss 0.534295f
C2591 por_dig_0.otrip_decoded[1] dvss 2.63538f
C2592 a_34573_28557# dvss 0.230498f
C2593 a_34467_28557# dvss 0.212635f
C2594 a_34290_28557# dvss 0.218905f
C2595 a_33971_28557# dvss 0.277531f
C2596 a_33155_28640# dvss 0.22912f
C2597 por_dig_0.net12 dvss 0.474535f
C2598 a_32701_28531# dvss 0.334929f
C2599 por_dig_0.net3 dvss 0.427479f
C2600 a_31360_28557# dvss 0.273019f
C2601 por_dig_0.otrip_decoded[6] dvss 3.869673f
C2602 a_35960_29101# dvss 0.327517f
C2603 por_dig_0.net17 dvss 0.614123f
C2604 por_dig_0.net11 dvss 1.32322f
C2605 por_dig_0.net15 dvss 0.731015f
C2606 por_dig_0.net7 dvss 3.990962f
C2607 por_dig_0.net6 dvss 2.43654f
C2608 por_dig_0.net5 dvss 3.124185f
C2609 a_34828_29253# dvss 0.310914f
C2610 por_dig_0.net9 dvss 0.728411f
C2611 por_dig_0.force_pdnb dvss 5.16598f
C2612 a_31413_29075# dvss 0.353378f
C2613 por_dig_0.osc_ena dvss 26.099129f
C2614 a_36328_29645# dvss 0.395978f
C2615 a_35556_29619# dvss 0.411875f
C2616 a_35298_29619# dvss 0.394245f
C2617 a_35202_29877# dvss 0.238278f
C2618 a_34496_29645# dvss 0.378687f
C2619 a_33852_29645# dvss 0.367043f
C2620 por_dig_0.net30 dvss 0.455623f
C2621 a_31776_29864# dvss 0.262061f
C2622 a_31413_29619# dvss 0.314853f
C2623 a_38053_30189# dvss 0.268968f
C2624 a_38228_30163# dvss 0.497809f
C2625 a_37488_30189# dvss 0.256733f
C2626 a_37706_30431# dvss 0.187359f
C2627 a_37138_30189# dvss 0.29158f
C2628 a_36972_30189# dvss 0.649262f
C2629 por_dig_0.net29 dvss 0.88173f
C2630 a_36476_30163# dvss 0.411157f
C2631 a_36218_30163# dvss 0.388736f
C2632 a_36122_30341# dvss 0.232288f
C2633 a_35293_30189# dvss 0.269083f
C2634 a_35468_30163# dvss 0.508445f
C2635 a_34728_30189# dvss 0.290694f
C2636 a_34946_30431# dvss 0.203018f
C2637 a_34378_30189# dvss 0.323539f
C2638 por_dig_0._014_ dvss 0.574137f
C2639 a_34212_30189# dvss 0.683184f
C2640 por_dig_0.net2 dvss 0.485956f
C2641 por_dig_0.net10 dvss 0.493712f
C2642 a_32004_30189# dvss 0.239736f
C2643 a_31651_30341# dvss 0.211356f
C2644 a_39497_30849# dvss 0.248151f
C2645 a_37777_31111# dvss 0.271498f
C2646 a_37952_31037# dvss 0.487788f
C2647 a_37212_31111# dvss 0.257257f
C2648 a_37430_30707# dvss 0.185656f
C2649 a_36862_30739# dvss 0.30057f
C2650 a_36696_30739# dvss 0.607855f
C2651 a_34098_30707# dvss 2.06157f
C2652 a_33269_31111# dvss 0.27467f
C2653 a_33444_31037# dvss 0.525342f
C2654 a_32704_31111# dvss 0.279218f
C2655 a_32922_30707# dvss 0.19942f
C2656 a_32354_30739# dvss 0.318008f
C2657 a_32188_30739# dvss 0.566937f
C2658 a_31864_30823# dvss 0.219358f
C2659 por_dig_0._038_ dvss 0.240102f
C2660 a_31592_30965# dvss 0.35305f
C2661 a_38904_31277# dvss 0.17078f
C2662 por_dig_0._003_ dvss 0.739811f
C2663 por_dig_0._004_ dvss 0.59653f
C2664 por_dig_0._043_ dvss 0.631373f
C2665 a_39510_31251# dvss 0.265957f
C2666 a_39077_31527# dvss 0.249618f
C2667 por_dig_0._044_ dvss 0.159151f
C2668 a_38500_31251# dvss 0.430824f
C2669 a_38242_31251# dvss 0.398572f
C2670 a_38146_31429# dvss 0.213359f
C2671 a_37751_31251# dvss 0.207257f
C2672 por_dig_0.net34 dvss 0.329308f
C2673 a_37392_31251# dvss 0.389154f
C2674 a_36305_31277# dvss 0.262583f
C2675 a_36480_31251# dvss 0.484427f
C2676 a_35740_31277# dvss 0.264561f
C2677 a_35958_31519# dvss 0.176508f
C2678 a_35390_31277# dvss 0.301357f
C2679 por_dig_0._015_ dvss 0.619478f
C2680 a_35224_31277# dvss 0.507709f
C2681 a_33940_31277# dvss 0.231785f
C2682 a_33374_31277# dvss 0.194529f
C2683 por_dig_0._027_ dvss 0.874481f
C2684 a_34852_31277# dvss 0.267339f
C2685 a_34746_31277# dvss 0.396914f
C2686 a_34510_31277# dvss 0.373061f
C2687 a_33804_31251# dvss 0.254674f
C2688 por_ana_0.sky130_fd_sc_hd__inv_4_1.Y dvss 2.05013f
C2689 por_ana_0.sky130_fd_sc_hd__inv_4_1.A dvss 0.775852f
C2690 por_ana_0.sky130_fd_sc_hd__inv_4_0.Y dvss 1.95044f
C2691 por_ana_0.schmitt_trigger_0.m dvss 2.177533f
C2692 por_ana_0.sky130_fd_sc_hd__inv_4_3.Y dvss 1.97752f
C2693 por_ana_0.sky130_fd_sc_hd__inv_4_4.Y dvss 1.98989f
C2694 a_8969_15512# dvss 0.639031f
C2695 a_8591_22912# dvss 0.502711f
C2696 a_8213_15512# dvss 0.639742f
C2697 a_7835_22912# dvss 0.502711f
C2698 a_7457_15512# dvss 0.646835f
C2699 a_7079_22912# dvss 0.502711f
C2700 a_6701_15512# dvss 0.639742f
C2701 a_6323_22912# dvss 0.502711f
C2702 a_5945_15512# dvss 0.639742f
C2703 a_5567_22912# dvss 0.502711f
C2704 a_5189_15512# dvss 0.639742f
C2705 a_4811_22912# dvss 0.502711f
C2706 a_4433_15512# dvss 0.639742f
C2707 a_4055_22912# dvss 0.502711f
C2708 a_3677_15512# dvss 0.639742f
C2709 a_3299_22912# dvss 0.502711f
C2710 a_2921_15512# dvss 0.639742f
C2711 a_2543_22912# dvss 0.502711f
C2712 a_2165_15512# dvss 0.614478f
C2713 a_32019_31643# dvss 0.185646f
C2714 a_32088_31514# dvss 0.264918f
C2715 a_31932_31419# dvss 0.62897f
C2716 a_31893_31545# dvss 0.301254f
C2717 a_31615_31529# dvss 0.274805f
C2718 a_31412_31251# dvss 0.50174f
C2719 por_dig_0._045_ dvss 0.413083f
C2720 a_37616_32141# dvss 0.181183f
C2721 a_36567_32141# dvss 0.202045f
C2722 a_35433_32141# dvss 0.177715f
C2723 por_dig_0._028_ dvss 0.762773f
C2724 por_dig_0.cnt_rsb dvss 0.511383f
C2725 a_39732_31829# dvss 0.317485f
C2726 a_39417_31795# dvss 0.2949f
C2727 a_38936_32159# dvss 0.261117f
C2728 a_37789_31821# dvss 0.25658f
C2729 por_dig_0._032_ dvss 0.484905f
C2730 por_dig_0._042_ dvss 2.47467f
C2731 por_dig_0.cnt_st\[4\] dvss 1.064f
C2732 a_36382_31795# dvss 0.301798f
C2733 por_dig_0._037_ dvss 1.40386f
C2734 a_35000_31795# dvss 0.268709f
C2735 a_34116_31821# dvss 0.209869f
C2736 a_34010_31821# dvss 0.355541f
C2737 a_33774_31821# dvss 0.351466f
C2738 por_dig_0.cnt_por\[9\] dvss 0.817876f
C2739 por_dig_0.cnt_por\[8\] dvss 1.37275f
C2740 por_dig_0.cnt_por\[10\] dvss 0.83742f
C2741 a_32441_32199# dvss 0.272411f
C2742 a_32616_32125# dvss 0.504085f
C2743 a_31876_32199# dvss 0.260641f
C2744 por_dig_0.net8 dvss 1.55159f
C2745 a_32094_31795# dvss 0.181538f
C2746 a_31526_31827# dvss 0.304913f
C2747 a_31360_31827# dvss 0.699432f
C2748 por_dig_0._031_ dvss 1.95506f
C2749 por_dig_0._036_ dvss 1.432947f
C2750 a_34486_32365# dvss 0.213359f
C2751 por_dig_0._013_ dvss 0.748917f
C2752 por_dig_0.cnt_st\[3\] dvss 1.04416f
C2753 a_38956_32339# dvss 0.256662f
C2754 a_38352_32365# dvss 0.249873f
C2755 por_dig_0._035_ dvss 0.93037f
C2756 a_36564_32339# dvss 0.340524f
C2757 a_36100_32517# dvss 0.247446f
C2758 a_35640_32517# dvss 0.235159f
C2759 por_dig_0.net27 dvss 1.66642f
C2760 a_35100_32339# dvss 0.548573f
C2761 por_dig_0.net32 dvss 0.535324f
C2762 por_dig_0._026_ dvss 0.928339f
C2763 a_34444_32517# dvss 0.254412f
C2764 a_33805_32339# dvss 0.314329f
C2765 a_32809_32365# dvss 0.273158f
C2766 a_32984_32339# dvss 0.4887f
C2767 a_32244_32365# dvss 0.265952f
C2768 a_32462_32607# dvss 0.184641f
C2769 a_31894_32365# dvss 0.296168f
C2770 a_31728_32365# dvss 0.600767f
C2771 por_dig_0.net19 dvss 1.79011f
C2772 a_31413_32339# dvss 0.314835f
C2773 a_39630_33229# dvss 0.164227f
C2774 por_dig_0.net28 dvss 0.418359f
C2775 a_25863_32638# dvss 1.69345f
C2776 por_dig_0._030_ dvss 0.771854f
C2777 por_dig_0._041_ dvss 0.1877f
C2778 a_38957_32883# dvss 0.400143f
C2779 a_37961_33287# dvss 0.258338f
C2780 a_38136_33213# dvss 0.475257f
C2781 a_37396_33287# dvss 0.274149f
C2782 a_37614_32883# dvss 0.189998f
C2783 a_37046_32915# dvss 0.31817f
C2784 por_dig_0._002_ dvss 0.260394f
C2785 a_36880_32915# dvss 0.543472f
C2786 a_34387_32909# dvss 2.01048f
C2787 a_33545_33287# dvss 0.262397f
C2788 a_33720_33213# dvss 0.492859f
C2789 a_32980_33287# dvss 0.254696f
C2790 a_33198_32883# dvss 0.180058f
C2791 a_32630_32915# dvss 0.295885f
C2792 a_32464_32915# dvss 0.57102f
C2793 por_dig_0.clknet_1_0__leaf_osc_ck dvss 4.863647f
C2794 a_31908_32909# dvss 0.233198f
C2795 a_31802_32909# dvss 0.373978f
C2796 a_31566_32909# dvss 0.389637f
C2797 por_dig_0.cnt_rsb_stg1 dvss 0.427499f
C2798 por_dig_0._040_ dvss 0.429313f
C2799 por_dig_0.net33 dvss 0.325385f
C2800 a_39718_33605# dvss 0.231325f
C2801 a_39268_33453# dvss 0.220833f
C2802 a_39162_33453# dvss 0.36477f
C2803 a_38926_33453# dvss 0.398955f
C2804 por_dig_0.cnt_st\[2\] dvss 0.809782f
C2805 a_37961_33453# dvss 0.264811f
C2806 a_38136_33427# dvss 0.49602f
C2807 a_37396_33453# dvss 0.260195f
C2808 a_37614_33695# dvss 0.180187f
C2809 a_37046_33453# dvss 0.293799f
C2810 por_dig_0._001_ dvss 1.38534f
C2811 a_36880_33453# dvss 0.632453f
C2812 por_dig_0._010_ dvss 0.944998f
C2813 a_35699_33819# dvss 0.18811f
C2814 a_35768_33690# dvss 0.265945f
C2815 a_35612_33595# dvss 0.66609f
C2816 a_35573_33721# dvss 0.306155f
C2817 a_35295_33705# dvss 0.269636f
C2818 a_35092_33427# dvss 0.494098f
C2819 por_dig_0.cnt_por\[5\] dvss 0.843921f
C2820 por_dig_0.cnt_por\[4\] dvss 1.20545f
C2821 a_34357_33427# dvss 0.319182f
C2822 por_dig_0._021_ dvss 0.243403f
C2823 a_33806_33427# dvss 0.268235f
C2824 por_dig_0.cnt_por\[7\] dvss 0.622451f
C2825 a_26288_32594# dvss 0.891608f
C2826 a_32019_33819# dvss 0.194554f
C2827 a_32088_33690# dvss 0.278465f
C2828 a_31932_33595# dvss 0.551605f
C2829 a_31893_33721# dvss 0.30233f
C2830 a_31615_33705# dvss 0.259832f
C2831 a_31412_33427# dvss 0.4827f
C2832 por_dig_0._029_ dvss 0.387779f
C2833 a_35582_34317# dvss 0.196128f
C2834 por_dig_0._009_ dvss 0.314556f
C2835 por_dig_0._011_ dvss 0.447596f
C2836 a_35040_34317# dvss 0.162559f
C2837 por_dig_0._020_ dvss 0.323506f
C2838 por_dig_0._012_ dvss 0.380846f
C2839 por_dig_0.net21 dvss 1.40053f
C2840 por_dig_0.cnt_st\[1\] dvss 1.39054f
C2841 por_dig_0._039_ dvss 0.909561f
C2842 a_38145_34375# dvss 0.267047f
C2843 a_38320_34301# dvss 0.498337f
C2844 a_37580_34375# dvss 0.25679f
C2845 por_dig_0.net25 dvss 4.37773f
C2846 a_37798_33971# dvss 0.179609f
C2847 a_37230_34003# dvss 0.291264f
C2848 por_dig_0._000_ dvss 0.388445f
C2849 a_37064_34003# dvss 0.685006f
C2850 a_36380_33971# dvss 0.393557f
C2851 por_dig_0._017_ dvss 0.323377f
C2852 por_dig_0._018_ dvss 0.230693f
C2853 por_dig_0._023_ dvss 0.31248f
C2854 por_dig_0._022_ dvss 0.196188f
C2855 a_34580_34110# dvss 0.253752f
C2856 por_dig_0.cnt_por\[6\] dvss 3.06436f
C2857 a_33600_34335# dvss 0.216171f
C2858 por_dig_0.net22 dvss 2.465436f
C2859 por_dig_0._019_ dvss 1.41516f
C2860 por_dig_0._025_ dvss 0.299053f
C2861 por_dig_0._024_ dvss 0.397571f
C2862 a_32794_33971# dvss 0.274178f
C2863 por_dig_0.net26 dvss 1.14393f
C2864 por_dig_0._137__26.LO dvss 0.109179f
C2865 a_26802_33372# dvss 0.506452f
C2866 a_25595_33708# dvss 1.5407f
C2867 a_25495_33620# dvss 2.02903f
C2868 por_dig_0.net1 dvss 0.594622f
C2869 a_31360_33997# dvss 0.266867f
C2870 por_dig_0.net31 dvss 0.489147f
C2871 por_dig_0.net4 dvss 3.41785f
C2872 por_dig_0.cnt_st\[0\] dvss 1.85298f
C2873 a_39328_34515# dvss 0.420633f
C2874 a_39070_34515# dvss 0.429148f
C2875 a_38974_34693# dvss 0.254547f
C2876 a_35583_34541# dvss 1.98572f
C2877 por_dig_0.clknet_0_osc_ck dvss 2.961383f
C2878 a_35040_34587# dvss 0.240476f
C2879 a_37409_35463# dvss 0.283602f
C2880 a_37584_35389# dvss 0.64359f
C2881 a_36844_35463# dvss 0.257515f
C2882 a_37062_35059# dvss 0.187382f
C2883 a_36494_35091# dvss 0.316105f
C2884 a_36328_35091# dvss 0.658569f
C2885 a_35704_35124# dvss 0.252068f
C2886 por_dig_0._046_ dvss 0.36484f
C2887 a_35450_35124# dvss 0.28937f
C2888 a_34672_35451# dvss 0.272753f
C2889 a_33821_35463# dvss 0.269524f
C2890 a_33996_35389# dvss 0.491531f
C2891 a_33256_35463# dvss 0.27368f
C2892 a_33474_35059# dvss 0.187573f
C2893 a_32906_35091# dvss 0.339645f
C2894 a_32740_35091# dvss 0.700583f
C2895 a_35024_35629# dvss 0.262738f
C2896 a_34580_35629# dvss 0.326744f
C2897 a_36581_35629# dvss 0.287456f
C2898 a_36756_35603# dvss 0.864129f
C2899 a_36016_35629# dvss 0.265707f
C2900 a_36234_35871# dvss 0.190162f
C2901 a_35666_35629# dvss 0.306105f
C2902 por_dig_0._005_ dvss 0.619131f
C2903 a_35500_35629# dvss 0.578178f
C2904 por_dig_0._034_ dvss 1.813131f
C2905 por_dig_0._008_ dvss 0.523559f
C2906 por_dig_0.cnt_por\[3\] dvss 1.15782f
C2907 a_33896_35603# dvss 0.252949f
C2908 por_dig_0._053_ dvss 0.536011f
C2909 a_33162_35603# dvss 0.278554f
C2910 por_dig_0._051_ dvss 0.644875f
C2911 por_dig_0._047_ dvss 1.66549f
C2912 a_32610_35603# dvss 0.299079f
C2913 por_dig_0._006_ dvss 0.434393f
C2914 a_36328_36493# dvss 0.198276f
C2915 por_dig_0._052_ dvss 0.336732f
C2916 por_dig_0._048_ dvss 1.30139f
C2917 por_dig_0._050_ dvss 0.216649f
C2918 a_35592_36286# dvss 0.256178f
C2919 por_dig_0.cnt_por\[2\] dvss 1.42661f
C2920 a_34633_36147# dvss 0.389318f
C2921 a_33821_36551# dvss 0.271886f
C2922 a_33996_36477# dvss 0.494284f
C2923 a_33256_36551# dvss 0.271821f
C2924 por_dig_0.net24 dvss 6.35507f
C2925 a_33474_36147# dvss 0.188733f
C2926 a_32906_36179# dvss 0.297354f
C2927 por_dig_0._007_ dvss 0.343057f
C2928 a_32740_36179# dvss 0.68436f
C2929 por_dig_0.clknet_1_1__leaf_osc_ck dvss 4.445326f
C2930 por_dig_0.por_unbuf dvss 10.65833f
C2931 por_dig_0._049_ dvss 0.504484f
C2932 por_dig_0._016_ dvss 0.927091f
C2933 a_36381_36691# dvss 0.371116f
C2934 por_dig_0.cnt_por\[1\] dvss 2.19138f
C2935 por_dig_0.cnt_por\[0\] dvss 3.317825f
C2936 por_dig_0.net23 dvss 4.048819f
C2937 por_dig_0.net20 dvss 2.61139f
C2938 por_dig_0._033_ dvss 2.1776f
C2939 por_ana_0.ibias_gen_0.vp1 dvss 4.776463f
C2940 por_ana_0.schmitt_trigger_0.in dvss 0.407856p
C2941 a_21178_35244# dvss 0.502711f
C2942 a_20800_27844# dvss 0.502711f
C2943 a_20422_35244# dvss 0.502711f
C2944 a_20044_27844# dvss 0.502711f
C2945 a_19666_35244# dvss 0.502711f
C2946 a_19288_27844# dvss 0.502711f
C2947 a_18910_35244# dvss 0.502711f
C2948 a_18532_27844# dvss 0.502711f
C2949 a_18154_35244# dvss 0.502711f
C2950 a_17776_27844# dvss 0.502711f
C2951 a_17398_35244# dvss 0.502711f
C2952 a_17020_27844# dvss 0.502711f
C2953 a_16642_35244# dvss 0.502711f
C2954 a_16264_27844# dvss 0.502711f
C2955 a_15886_35244# dvss 0.502711f
C2956 a_15508_27844# dvss 0.502711f
C2957 a_15130_35244# dvss 0.502711f
C2958 a_14752_27844# dvss 0.502711f
C2959 por_ana_0.vl dvss 6.05527f
C2960 a_14374_35244# dvss 0.502711f
C2961 por_ana_0.dcomp3v3 dvss 1.18668f
C2962 por_ana_0.comparator_1.n0 dvss 4.818092f
C2963 por_ana_0.comparator_1.vm dvss 9.239901f
C2964 por_ana_0.comparator_1.vn dvss 5.471683f
C2965 por_ana_0.comparator_1.ena_b dvss 0.625987f
C2966 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A dvss 0.460997f
C2967 por_ana_0.sky130_fd_sc_hvl__inv_4_0.A dvss 0.477453f
C2968 por_ana_0.sky130_fd_sc_hvl__inv_1_0.A dvss 2.32373f
C2969 por_ana_0.comparator_1.vnn dvss 33.55585f
C2970 itest.n0 dvss 1.68127f
C2971 por_ana_0.rstring_mux_0.vtrip1.t7 dvss 0.216167f
C2972 por_ana_0.rstring_mux_0.vtrip1.n0 dvss 0.234604f
C2973 por_ana_0.rstring_mux_0.vtrip1.n1 dvss 0.15382f
C2974 por_ana_0.rstring_mux_0.vtrip1.n2 dvss 0.961398f
C2975 por_ana_0.rstring_mux_0.vtrip1.n3 dvss 0.234604f
C2976 por_ana_0.rstring_mux_0.vtrip1.n4 dvss 0.15382f
C2977 por_ana_0.rstring_mux_0.vtrip1.n5 dvss 1.52407f
C2978 por_ana_0.rstring_mux_0.vtrip1.n6 dvss 1.30427f
C2979 por_ana_0.rstring_mux_0.vtrip1.n7 dvss 3.51872f
C2980 por_ana_0.rstring_mux_0.vtrip1.t4 dvss 0.21619f
C2981 por_ana_0.comparator_1.vn.n0 dvss 3.53898f
C2982 por_ana_0.comparator_1.vn.n1 dvss 0.64177f
C2983 por_ana_0.comparator_1.vn.n2 dvss 1.13914f
C2984 por_ana_0.comparator_1.vn.t7 dvss 1.97015f
C2985 por_ana_0.comparator_1.vn.t8 dvss 1.70312f
C2986 por_ana_0.comparator_1.vn.t5 dvss 1.70312f
C2987 por_ana_0.comparator_1.vn.t3 dvss 1.84324f
C2988 por_ana_0.comparator_0.ibias.t1 dvss 0.101238f
C2989 por_ana_0.comparator_0.ibias.n0 dvss 9.838731f
C2990 por_ana_0.comparator_0.ibias.n1 dvss 4.99964f
C2991 por_ana_0.comparator_0.ibias.t2 dvss 0.101238f
C2992 por_ana_0.ibias_gen_0.vr.n0 dvss 0.183081f
C2993 por_ana_0.ibias_gen_0.vr.n1 dvss 0.161866f
C2994 por_ana_0.ibias_gen_0.vr.n2 dvss 1.54735f
C2995 por_ana_0.ibias_gen_0.vr.t4 dvss 0.540543f
C2996 por_ana_0.comparator_0.n0.n0 dvss 1.17312f
C2997 por_ana_0.comparator_0.n0.t7 dvss 0.173496f
C2998 por_ana_0.comparator_0.n0.t5 dvss 0.173312f
C2999 por_ana_0.comparator_0.n0.n2 dvss 0.364558f
C3000 por_ana_0.comparator_0.n0.t8 dvss 0.168852f
C3001 por_ana_0.comparator_0.n0.t6 dvss 0.168669f
C3002 por_ana_0.comparator_0.n0.t4 dvss 0.158872f
C3003 force_pdn.n3 dvss 1.11667f
C3004 force_pdn.n4 dvss 0.792682f
C3005 force_dis_rc_osc.n3 dvss 0.946473f
C3006 force_dis_rc_osc.n4 dvss 0.614422f
C3007 por_ana_0.sky130_fd_sc_hvl__lsbuflv2hv_1_0[1|6].X dvss 0.153815f
C3008 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[5].t5 dvss 0.402957f
C3009 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[5].t4 dvss 0.402805f
C3010 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[5].n2 dvss 0.388303f
C3011 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[5].n5 dvss 1.87247f
C3012 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[5].n6 dvss 1.02015f
C3013 otrip[0].n4 dvss 3.10696f
C3014 otrip[0].n5 dvss 1.75839f
C3015 ibg_200n.t1 dvss 0.222198f
C3016 ibg_200n.t0 dvss 0.270728f
C3017 ibg_200n.n0 dvss 2.74902f
C3018 por_dig_0.otrip_decoded[0].n0 dvss 8.50069f
C3019 por_dig_0.otrip_decoded[0].n4 dvss 0.100675f
C3020 por_dig_0.otrip_decoded[0].n6 dvss 3.84731f
C3021 por_ana_0.rstring_mux_0.vtrip4.t7 dvss 0.171176f
C3022 por_ana_0.rstring_mux_0.vtrip4.n0 dvss 0.18541f
C3023 por_ana_0.rstring_mux_0.vtrip4.n1 dvss 0.121565f
C3024 por_ana_0.rstring_mux_0.vtrip4.n2 dvss 1.18871f
C3025 por_ana_0.rstring_mux_0.vtrip4.n3 dvss 0.18541f
C3026 por_ana_0.rstring_mux_0.vtrip4.n4 dvss 0.121565f
C3027 por_ana_0.rstring_mux_0.vtrip4.n5 dvss 0.749847f
C3028 por_ana_0.rstring_mux_0.vtrip4.n6 dvss 1.88677f
C3029 por_ana_0.rstring_mux_0.vtrip4.n7 dvss 2.28683f
C3030 por_ana_0.rstring_mux_0.vtrip4.t0 dvss 0.726836f
C3031 por_ana_0.ibias_gen_0.ve.n0 dvss -12.936501f
C3032 por_ana_0.ibias_gen_0.ve.t1 dvss 13.1014f
C3033 por_ana_0.ibias_gen_0.ve.t2 dvss 0.129205f
C3034 por_ana_0.ibias_gen_0.ve.t4 dvss 0.129205f
C3035 por_ana_0.ibias_gen_0.ve.n2 dvss 0.510582f
C3036 por_ana_0.ibias_gen_0.ve.t3 dvss 0.129205f
C3037 por_ana_0.ibias_gen_0.ve.t0 dvss 0.129205f
C3038 por_ana_0.ibias_gen_0.ve.n3 dvss 0.54803f
C3039 por_ana_0.ibias_gen_0.ve.n4 dvss 10.5378f
C3040 por_ana_0.ibias_gen_0.ve.n5 dvss 11.8523f
C3041 force_ena_rc_osc.n3 dvss 2.26949f
C3042 force_ena_rc_osc.n4 dvss 1.51058f
C3043 por_ana_0.ibias_gen_0.ena_b.n0 dvss 0.149893f
C3044 por_ana_0.ibias_gen_0.ena_b.t5 dvss 0.511691f
C3045 por_ana_0.ibias_gen_0.ena_b.t6 dvss 0.504751f
C3046 por_ana_0.ibias_gen_0.ena_b.n1 dvss 0.96914f
C3047 por_ana_0.ibias_gen_0.ena_b.t4 dvss 1.60711f
C3048 por_ana_0.ibias_gen_0.ena_b.t7 dvss 1.60105f
C3049 por_ana_0.ibias_gen_0.ena_b.n2 dvss 1.06345f
C3050 por_ana_0.ibias_gen_0.ena_b.n3 dvss 0.862249f
C3051 por_ana_0.ibias_gen_0.ena_b.n4 dvss 0.88086f
C3052 por_ana_0.ibias_gen_0.ena_b.n5 dvss 0.206991f
C3053 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[4].t3 dvss 0.218655f
C3054 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[4].t4 dvss 0.218573f
C3055 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[4].n2 dvss 0.210813f
C3056 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[4].n5 dvss 0.442354f
C3057 por_dig_0._036_.n5 dvss 0.598338f
C3058 por_dig_0._036_.n7 dvss 0.406869f
C3059 por_dig_0._036_.n8 dvss 0.200218f
C3060 por_ana_0.ibias_gen_0.isrc_sel_b.n0 dvss 0.450144f
C3061 por_ana_0.ibias_gen_0.isrc_sel_b.n1 dvss 1.93854f
C3062 por_ana_0.ibias_gen_0.isrc_sel_b.n2 dvss 0.153124f
C3063 por_ana_0.ibias_gen_0.isrc_sel_b.t7 dvss 0.501892f
C3064 por_ana_0.ibias_gen_0.isrc_sel_b.t4 dvss 0.511128f
C3065 por_ana_0.ibias_gen_0.isrc_sel_b.t6 dvss 0.507022f
C3066 por_ana_0.ibias_gen_0.isrc_sel_b.n3 dvss 0.523179f
C3067 por_ana_0.ibias_gen_0.isrc_sel_b.t5 dvss 1.64159f
C3068 por_ana_0.ibias_gen_0.isrc_sel_b.t8 dvss 1.66569f
C3069 por_ana_0.ibias_gen_0.isrc_sel_b.n4 dvss 0.860441f
C3070 por_ana_0.ibias_gen_0.isrc_sel_b.n5 dvss 0.203349f
C3071 por_ana_0.sky130_fd_sc_hvl__lsbuflv2hv_1_0[1|8].X dvss 0.239136f
C3072 por_ana_0.ibias_gen_0.isrc_sel.n0 dvss 9.46205f
C3073 por_ana_0.ibias_gen_0.isrc_sel.t8 dvss 0.708102f
C3074 por_ana_0.ibias_gen_0.isrc_sel.t5 dvss 0.702792f
C3075 por_ana_0.ibias_gen_0.isrc_sel.n3 dvss 0.871189f
C3076 por_ana_0.ibias_gen_0.isrc_sel.t7 dvss 0.712847f
C3077 por_ana_0.ibias_gen_0.isrc_sel.n4 dvss 0.595984f
C3078 por_ana_0.ibias_gen_0.isrc_sel.t3 dvss 0.591134f
C3079 por_ana_0.ibias_gen_0.isrc_sel.n5 dvss 0.878681f
C3080 por_ana_0.ibias_gen_0.isrc_sel.t9 dvss 2.34029f
C3081 por_ana_0.ibias_gen_0.isrc_sel.t6 dvss 2.36007f
C3082 por_ana_0.ibias_gen_0.isrc_sel.t4 dvss 1.15565f
C3083 por_ana_0.ibias_gen_0.isrc_sel.t2 dvss 1.17014f
C3084 por_ana_0.ibias_gen_0.isrc_sel.n6 dvss 1.18897f
C3085 por_ana_0.ibias_gen_0.isrc_sel.n7 dvss 3.58505f
C3086 por_ana_0.comparator_0.ena_b.n0 dvss 1.46363f
C3087 por_ana_0.comparator_0.ena_b.t5 dvss 0.213702f
C3088 por_ana_0.comparator_0.ena_b.t4 dvss 0.207774f
C3089 por_ana_0.comparator_0.ena_b.t3 dvss 0.207146f
C3090 por_ana_0.comparator_0.ena_b.t2 dvss 0.207146f
C3091 por_ana_0.comparator_1.vm.n0 dvss 2.33715f
C3092 por_ana_0.comparator_1.vm.t6 dvss 0.17369f
C3093 por_ana_0.comparator_1.vm.t7 dvss 2.77148f
C3094 por_ana_0.comparator_1.vm.t8 dvss 2.39583f
C3095 por_ana_0.comparator_1.vm.t4 dvss 2.39583f
C3096 por_ana_0.comparator_1.vm.t2 dvss 2.59294f
C3097 por_ana_0.comparator_0.vm.n0 dvss 2.35043f
C3098 por_ana_0.comparator_0.vm.t6 dvss 0.174677f
C3099 por_ana_0.comparator_0.vm.t7 dvss 2.78722f
C3100 por_ana_0.comparator_0.vm.t8 dvss 2.40944f
C3101 por_ana_0.comparator_0.vm.t0 dvss 2.40944f
C3102 por_ana_0.comparator_0.vm.t2 dvss 2.60767f
C3103 por_ana_0.rc_osc_0.n.t11 dvss 0.143388f
C3104 por_ana_0.rc_osc_0.n.t9 dvss 0.143249f
C3105 por_ana_0.rc_osc_0.n.n2 dvss 0.164777f
C3106 por_ana_0.rc_osc_0.n.t8 dvss 0.143249f
C3107 por_ana_0.rc_osc_0.n.n3 dvss 0.156263f
C3108 por_ana_0.rc_osc_0.n.t10 dvss 0.14446f
C3109 por_ana_0.rc_osc_0.n.n4 dvss 0.529644f
C3110 por_ana_0.rc_osc_0.n.t12 dvss 0.287357f
C3111 por_ana_0.rc_osc_0.n.t13 dvss 0.286497f
C3112 por_ana_0.rc_osc_0.n.n5 dvss 0.277287f
C3113 por_ana_0.rc_osc_0.n.t7 dvss 0.287213f
C3114 por_ana_0.rc_osc_0.n.n6 dvss 0.196012f
C3115 por_ana_0.rc_osc_0.n.t6 dvss 0.283047f
C3116 por_ana_0.rc_osc_0.n.n7 dvss 0.360416f
C3117 por_ana_0.rc_osc_0.n.n8 dvss 0.222174f
C3118 por_ana_0.rc_osc_0.n.n9 dvss 0.477653f
C3119 por_ana_0.rc_osc_0.n.n10 dvss 0.555032f
C3120 por_ana_0.sky130_fd_sc_hvl__lsbuflv2hv_1_0[0|8].X dvss 0.226888f
C3121 por_ana_0.rstring_mux_0.ena.n0 dvss 1.32231f
C3122 por_ana_0.rstring_mux_0.ena.n1 dvss 5.11834f
C3123 por_ana_0.rstring_mux_0.ena.n2 dvss 0.727712f
C3124 por_ana_0.rstring_mux_0.ena.n3 dvss 4.36283f
C3125 por_ana_0.rstring_mux_0.ena.t13 dvss 0.942417f
C3126 por_ana_0.rstring_mux_0.ena.t3 dvss 0.93785f
C3127 por_ana_0.rstring_mux_0.ena.t8 dvss 1.85232f
C3128 por_ana_0.rstring_mux_0.ena.t5 dvss 0.226724f
C3129 por_ana_0.rstring_mux_0.ena.t7 dvss 0.22603f
C3130 por_ana_0.rstring_mux_0.ena.t6 dvss 0.22603f
C3131 por_ana_0.rstring_mux_0.ena.t2 dvss 0.222066f
C3132 por_ana_0.rstring_mux_0.ena.t10 dvss 0.220765f
C3133 por_ana_0.rstring_mux_0.ena.t4 dvss 0.569038f
C3134 por_ana_0.rstring_mux_0.ena.t11 dvss 2.03175f
C3135 por_ana_0.rstring_mux_0.ena.t1 dvss 2.03868f
C3136 por_ana_0.rstring_mux_0.ena.n6 dvss 0.254369f
C3137 por_ana_0.rstring_mux_0.ena.n7 dvss 3.59107f
C3138 por_ana_0.rstring_mux_0.sky130_fd_sc_hvl__inv_1_1.A dvss 0.129333f
C3139 por_ana_0.rstring_mux_0.ena.t12 dvss 0.115978f
C3140 por_ana_0.rstring_mux_0.ena.n8 dvss 0.101063f
C3141 por_ana_0.rstring_mux_0.ena.n10 dvss 11.322f
C3142 por_ana_0.rstring_mux_0.ena.n11 dvss 1.8749f
C3143 por_dig_0.otrip_decoded[2].n5 dvss 0.586277f
C3144 por_dig_0.osc_ena.t7 dvss 0.147442f
C3145 por_dig_0.osc_ena.n0 dvss 0.414577f
C3146 por_dig_0.osc_ena.t4 dvss 0.151346f
C3147 por_dig_0.osc_ena.n1 dvss 0.178359f
C3148 por_ana_0.comparator_0.vn.n0 dvss 3.61821f
C3149 por_ana_0.comparator_0.vn.n1 dvss 0.656138f
C3150 por_ana_0.comparator_0.vn.n2 dvss 1.16465f
C3151 por_ana_0.comparator_0.vn.t7 dvss 2.01426f
C3152 por_ana_0.comparator_0.vn.t8 dvss 1.74125f
C3153 por_ana_0.comparator_0.vn.t1 dvss 1.74125f
C3154 por_ana_0.comparator_0.vn.t3 dvss 1.88451f
C3155 otrip[1].n1 dvss 0.117098f
C3156 otrip[1].n3 dvss 3.63341f
C3157 otrip[1].n4 dvss 2.06762f
C3158 por_dig_0.otrip_decoded[7].n0 dvss 5.30962f
C3159 por_dig_0.otrip_decoded[7].n4 dvss 0.103821f
C3160 por_dig_0.otrip_decoded[7].n6 dvss 2.10778f
C3161 por_ana_0.rstring_mux_0.vtrip7.t7 dvss 0.16069f
C3162 por_ana_0.rstring_mux_0.vtrip7.n0 dvss 0.174395f
C3163 por_ana_0.rstring_mux_0.vtrip7.n1 dvss 0.114343f
C3164 por_ana_0.rstring_mux_0.vtrip7.n2 dvss 0.752155f
C3165 por_ana_0.rstring_mux_0.vtrip7.n3 dvss 0.174395f
C3166 por_ana_0.rstring_mux_0.vtrip7.n4 dvss 0.114343f
C3167 por_ana_0.rstring_mux_0.vtrip7.n5 dvss 1.19247f
C3168 por_ana_0.rstring_mux_0.vtrip7.n6 dvss 0.918289f
C3169 por_ana_0.rstring_mux_0.vtrip7.n7 dvss 2.50533f
C3170 por_ana_0.rstring_mux_0.vtrip7.t6 dvss 0.160707f
C3171 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[7].t2 dvss 0.257237f
C3172 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[7].t3 dvss 0.25714f
C3173 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[7].n2 dvss 0.25938f
C3174 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[7].n5 dvss 1.25258f
C3175 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[7].n6 dvss 0.745985f
C3176 por_dig_0.net20.n4 dvss 0.131616f
C3177 por_dig_0.net20.n5 dvss 0.415396f
C3178 por_dig_0.net20.n8 dvss 0.414104f
C3179 por_dig_0.net20.n11 dvss 0.461008f
C3180 por_ana_0.rstring_mux_0.vtrip0.t7 dvss 0.17627f
C3181 por_ana_0.rstring_mux_0.vtrip0.n0 dvss 0.190942f
C3182 por_ana_0.rstring_mux_0.vtrip0.n1 dvss 0.125183f
C3183 por_ana_0.rstring_mux_0.vtrip0.n2 dvss 0.776085f
C3184 por_ana_0.rstring_mux_0.vtrip0.n3 dvss 0.190927f
C3185 por_ana_0.rstring_mux_0.vtrip0.n4 dvss 0.125183f
C3186 por_ana_0.rstring_mux_0.vtrip0.n5 dvss 1.22742f
C3187 por_ana_0.rstring_mux_0.vtrip0.n6 dvss 2.02058f
C3188 por_ana_0.rstring_mux_0.vtrip0.n7 dvss 2.41105f
C3189 por_ana_0.rstring_mux_0.vtrip0.t0 dvss 0.748466f
C3190 por_ana_0.ibias_gen_0.vp1.n0 dvss 2.2551f
C3191 por_ana_0.ibias_gen_0.vp1.t12 dvss 2.72493f
C3192 por_ana_0.ibias_gen_0.vp1.n1 dvss 0.130918f
C3193 por_ana_0.ibias_gen_0.vp1.n2 dvss 0.257085f
C3194 por_ana_0.ibias_gen_0.vp1.n3 dvss 2.14115f
C3195 por_ana_0.ibias_gen_0.vp1.t10 dvss 2.72114f
C3196 por_ana_0.ibias_gen_0.vp1.n4 dvss 0.225585f
C3197 por_ana_0.ibias_gen_0.vp1.n5 dvss 0.978301f
C3198 por_ana_0.ibias_gen_0.vp1.n6 dvss 0.154917f
C3199 por_ana_0.ibias_gen_0.vp1.n7 dvss 0.213443f
C3200 por_ana_0.ibias_gen_0.vp1.n8 dvss 0.168888f
C3201 por_ana_0.ibias_gen_0.vp1.n9 dvss 0.998605f
C3202 por_ana_0.ibias_gen_0.vp1.n10 dvss 0.168888f
C3203 por_ana_0.ibias_gen_0.vp1.n11 dvss 0.677866f
C3204 por_ana_0.ibias_gen_0.vp1.n12 dvss 0.163248f
C3205 por_ana_0.ibias_gen_0.vp1.n13 dvss 0.666034f
C3206 por_ana_0.ibias_gen_0.vp1.n14 dvss 0.19773f
C3207 por_ana_0.ibias_gen_0.vp1.n15 dvss 0.829697f
C3208 por_ana_0.ibias_gen_0.vn1.n0 dvss 0.745323f
C3209 por_ana_0.ibias_gen_0.vn1.t2 dvss 2.11164f
C3210 por_ana_0.ibias_gen_0.vn1.t16 dvss 2.11164f
C3211 por_ana_0.ibias_gen_0.vn1.t11 dvss 2.19722f
C3212 por_ana_0.ibias_gen_0.vn1.n2 dvss 1.40052f
C3213 por_ana_0.ibias_gen_0.vn1.t10 dvss 2.11164f
C3214 por_ana_0.ibias_gen_0.vn1.t12 dvss 2.19722f
C3215 por_ana_0.ibias_gen_0.vn1.n3 dvss 1.3685f
C3216 por_ana_0.ibias_gen_0.vn1.n4 dvss 0.140807f
C3217 por_ana_0.ibias_gen_0.vn1.t13 dvss 2.11164f
C3218 por_ana_0.ibias_gen_0.vn1.t15 dvss 2.19722f
C3219 por_ana_0.ibias_gen_0.vn1.n5 dvss 1.40052f
C3220 por_ana_0.ibias_gen_0.vn1.t14 dvss 2.11164f
C3221 por_ana_0.ibias_gen_0.vn1.t17 dvss 2.19722f
C3222 por_ana_0.ibias_gen_0.vn1.n6 dvss 1.3685f
C3223 por_ana_0.ibias_gen_0.vn1.n7 dvss 0.140807f
C3224 por_ana_0.ibias_gen_0.vn1.n8 dvss 0.110984f
C3225 por_ana_0.ibias_gen_0.vn1.n9 dvss 0.705651f
C3226 por_ana_0.ibias_gen_0.vn1.t4 dvss 2.15704f
C3227 por_ana_0.ibias_gen_0.vn1.n10 dvss 0.71883f
C3228 por_ana_0.ibias_gen_0.vn1.n12 dvss 0.218051f
C3229 por_ana_0.ibias_gen_0.vn1.n13 dvss 0.120433f
C3230 por_dig_0.otrip_decoded[6].n5 dvss 1.91813f
C3231 por_dig_0.otrip_decoded[6].n6 dvss 4.41497f
C3232 por_ana_0.comparator_0.vt.n0 dvss 0.523395f
C3233 por_ana_0.comparator_0.vt.n1 dvss 0.801271f
C3234 por_ana_0.comparator_0.vt.n2 dvss 0.685785f
C3235 por_ana_0.comparator_0.vt.n3 dvss 0.496385f
C3236 por_ana_0.comparator_0.vt.n4 dvss 0.441765f
C3237 por_ana_0.comparator_0.vt.n5 dvss 0.797975f
C3238 por_ana_0.comparator_0.vt.n6 dvss 0.409965f
C3239 por_ana_0.comparator_0.vt.n7 dvss 0.797975f
C3240 por_ana_0.comparator_0.vt.n8 dvss 0.351948f
C3241 por_ana_0.comparator_0.vt.n9 dvss 0.514339f
C3242 por_ana_0.comparator_0.vt.n10 dvss 0.441765f
C3243 por_ana_0.comparator_0.vt.n11 dvss 0.409965f
C3244 por_ana_0.comparator_0.vt.n12 dvss 1.5498f
C3245 por_ana_0.comparator_0.vt.n13 dvss 1.49274f
C3246 por_ana_0.comparator_0.vt.n14 dvss 1.5498f
C3247 por_ana_0.comparator_0.vt.n15 dvss 1.49274f
C3248 por_ana_0.comparator_0.vt.n19 dvss 15.0811f
C3249 por_ana_0.comparator_0.vt.n20 dvss 1.80115f
C3250 por_ana_0.comparator_0.vt.n21 dvss 1.80115f
C3251 por_ana_0.comparator_0.vt.t21 dvss 24.817999f
C3252 por_ana_0.comparator_0.vt.t3 dvss 31.202501f
C3253 por_ana_0.comparator_0.vt.t36 dvss 23.401901f
C3254 por_ana_0.comparator_0.vt.n22 dvss 15.6012f
C3255 por_ana_0.comparator_0.vt.t40 dvss 23.401901f
C3256 por_ana_0.comparator_0.vt.t0 dvss 31.202501f
C3257 por_ana_0.comparator_0.vt.t18 dvss 24.817999f
C3258 por_ana_0.comparator_0.vt.n23 dvss 15.0811f
C3259 por_ana_0.comparator_0.vt.n31 dvss 0.657642f
C3260 por_ana_0.comparator_0.vt.n32 dvss 0.691554f
C3261 por_ana_0.comparator_0.vt.n33 dvss 0.695733f
C3262 por_ana_0.comparator_0.vt.n34 dvss 0.653967f
C3263 por_ana_0.comparator_0.vt.n36 dvss 0.653967f
C3264 por_ana_0.comparator_0.vt.n37 dvss 0.695733f
C3265 por_ana_0.comparator_0.vt.n38 dvss 0.691554f
C3266 por_ana_0.comparator_0.vt.n39 dvss 0.657642f
C3267 por_dig_0.otrip_decoded[3].n0 dvss 7.16931f
C3268 por_dig_0.otrip_decoded[3].n6 dvss 3.04427f
C3269 por_dig_0.otrip_decoded[5].n5 dvss 1.94776f
C3270 por_dig_0.otrip_decoded[5].n6 dvss 4.65989f
C3271 porb_h.n2 dvss 0.242179f
C3272 porb_h.n8 dvss 0.242179f
C3273 porb_h.n11 dvss 0.14665f
C3274 porb_h.n14 dvss 0.242179f
C3275 porb_h.n16 dvss 0.125734f
C3276 porb_h.n17 dvss 0.201073f
C3277 porb_h.n20 dvss 0.242179f
C3278 porb_h.n22 dvss 0.165959f
C3279 porb_h.n23 dvss 0.255495f
C3280 porb_h.n26 dvss 0.242179f
C3281 porb_h.n28 dvss 0.206184f
C3282 porb_h.n29 dvss 0.309917f
C3283 porb_h.n32 dvss 0.242179f
C3284 porb_h.n34 dvss 0.246409f
C3285 porb_h.n35 dvss 0.364339f
C3286 porb_h.n38 dvss 0.242179f
C3287 porb_h.n40 dvss 0.261752f
C3288 porb_h.n43 dvss 0.243049f
C3289 porb_h.n44 dvss 0.988928f
C3290 porb_h.n45 dvss 0.522358f
C3291 por_ana_0.comparator_0.n1.n0 dvss 0.765455f
C3292 por_ana_0.comparator_0.n1.n1 dvss 1.18081f
C3293 por_ana_0.comparator_0.n1.n2 dvss 0.795794f
C3294 por_ana_0.comparator_0.n1.t8 dvss 0.177538f
C3295 por_ana_0.comparator_0.n1.t19 dvss 0.177346f
C3296 por_ana_0.comparator_0.n1.t14 dvss 0.177346f
C3297 por_ana_0.comparator_0.n1.t13 dvss 0.177346f
C3298 por_ana_0.comparator_0.n1.t4 dvss 0.177346f
C3299 por_ana_0.comparator_0.n1.t15 dvss 0.177346f
C3300 por_ana_0.comparator_0.n1.t9 dvss 0.177346f
C3301 por_ana_0.comparator_0.n1.t5 dvss 0.177346f
C3302 por_ana_0.comparator_0.n1.t16 dvss 0.172786f
C3303 por_ana_0.comparator_0.n1.t10 dvss 0.172595f
C3304 por_ana_0.comparator_0.n1.t6 dvss 0.172595f
C3305 por_ana_0.comparator_0.n1.t17 dvss 0.172595f
C3306 por_ana_0.comparator_0.n1.t12 dvss 0.172595f
C3307 por_ana_0.comparator_0.n1.t7 dvss 0.172595f
C3308 por_ana_0.comparator_0.n1.t18 dvss 0.172595f
C3309 por_ana_0.comparator_0.n1.t11 dvss 0.172595f
C3310 por_ana_0.comparator_1.vt.n0 dvss 0.50117f
C3311 por_ana_0.comparator_1.vt.n1 dvss 0.692396f
C3312 por_ana_0.comparator_1.vt.n2 dvss 0.808996f
C3313 por_ana_0.comparator_1.vt.n3 dvss 0.692396f
C3314 por_ana_0.comparator_1.vt.n4 dvss 0.413917f
C3315 por_ana_0.comparator_1.vt.n5 dvss 0.805668f
C3316 por_ana_0.comparator_1.vt.n6 dvss 0.446024f
C3317 por_ana_0.comparator_1.vt.n7 dvss 0.805668f
C3318 por_ana_0.comparator_1.vt.n8 dvss 0.355341f
C3319 por_ana_0.comparator_1.vt.n9 dvss 0.355341f
C3320 por_ana_0.comparator_1.vt.n10 dvss 0.660272f
C3321 por_ana_0.comparator_1.vt.n11 dvss 0.70244f
C3322 por_ana_0.comparator_1.vt.n12 dvss 0.413917f
C3323 por_ana_0.comparator_1.vt.n13 dvss 0.446024f
C3324 por_ana_0.comparator_1.vt.n14 dvss 1.56474f
C3325 por_ana_0.comparator_1.vt.n15 dvss 0.70244f
C3326 por_ana_0.comparator_1.vt.n16 dvss 1.56474f
C3327 por_ana_0.comparator_1.vt.n17 dvss 1.50713f
C3328 por_ana_0.comparator_1.vt.n18 dvss 1.50713f
C3329 por_ana_0.comparator_1.vt.n20 dvss 1.81851f
C3330 por_ana_0.comparator_1.vt.n21 dvss 15.2265f
C3331 por_ana_0.comparator_1.vt.n22 dvss 15.2265f
C3332 por_ana_0.comparator_1.vt.t3 dvss 25.0573f
C3333 por_ana_0.comparator_1.vt.t36 dvss 31.5033f
C3334 por_ana_0.comparator_1.vt.t20 dvss 23.627499f
C3335 por_ana_0.comparator_1.vt.t0 dvss 25.0573f
C3336 por_ana_0.comparator_1.vt.t41 dvss 31.5033f
C3337 por_ana_0.comparator_1.vt.t18 dvss 23.627499f
C3338 por_ana_0.comparator_1.vt.n23 dvss 15.7517f
C3339 por_ana_0.comparator_1.vt.n24 dvss 1.81851f
C3340 por_ana_0.comparator_1.vt.n33 dvss 0.663982f
C3341 por_ana_0.comparator_1.vt.n34 dvss 0.698221f
C3342 por_ana_0.comparator_1.vt.n35 dvss 0.660272f
C3343 por_ana_0.comparator_1.vt.n44 dvss 0.663982f
C3344 por_ana_0.comparator_1.vt.n45 dvss 0.698221f
C3345 por_ana_0.comparator_1.vnn.n0 dvss 1.1742f
C3346 por_ana_0.comparator_1.vnn.n1 dvss 5.21987f
C3347 por_ana_0.comparator_1.vnn.n2 dvss 1.04141f
C3348 por_ana_0.comparator_1.vnn.n3 dvss 1.04141f
C3349 por_ana_0.comparator_1.vnn.n4 dvss 1.04141f
C3350 por_ana_0.comparator_1.vnn.n5 dvss 1.04141f
C3351 por_ana_0.comparator_1.vnn.n6 dvss 5.59691f
C3352 por_ana_0.comparator_1.vnn.n7 dvss 3.18503f
C3353 por_ana_0.comparator_1.vnn.t0 dvss 1.40931f
C3354 por_ana_0.comparator_1.vnn.t12 dvss 1.40931f
C3355 por_ana_0.comparator_1.vnn.t10 dvss 1.40931f
C3356 por_ana_0.comparator_1.vnn.t6 dvss 1.40931f
C3357 por_ana_0.comparator_1.vnn.t2 dvss 1.40931f
C3358 por_ana_0.comparator_1.vnn.t14 dvss 1.40931f
C3359 por_ana_0.comparator_1.vnn.t8 dvss 1.40931f
C3360 por_ana_0.comparator_1.vnn.t4 dvss 1.40931f
C3361 por_ana_0.comparator_1.vnn.t56 dvss 1.50501f
C3362 por_ana_0.comparator_1.vnn.t54 dvss 1.30362f
C3363 por_ana_0.comparator_1.vnn.t47 dvss 1.50501f
C3364 por_ana_0.comparator_1.vnn.t58 dvss 1.30362f
C3365 por_ana_0.comparator_1.vnn.t48 dvss 1.50501f
C3366 por_ana_0.comparator_1.vnn.t59 dvss 1.30362f
C3367 por_ana_0.comparator_1.vnn.t49 dvss 1.50501f
C3368 por_ana_0.comparator_1.vnn.t60 dvss 1.30362f
C3369 por_ana_0.comparator_1.vnn.t50 dvss 1.50501f
C3370 por_ana_0.comparator_1.vnn.t61 dvss 1.30362f
C3371 por_ana_0.comparator_1.vnn.t53 dvss 1.50501f
C3372 por_ana_0.comparator_1.vnn.t52 dvss 1.30362f
C3373 por_ana_0.comparator_1.vnn.t51 dvss 1.50501f
C3374 por_ana_0.comparator_1.vnn.t62 dvss 1.30362f
C3375 por_ana_0.comparator_1.vnn.t57 dvss 1.50501f
C3376 por_ana_0.comparator_1.vnn.t55 dvss 1.30362f
C3377 otrip[2].n4 dvss 1.84271f
C3378 otrip[2].n5 dvss 0.896023f
C3379 por_ana_0.ibias_gen_0.vstart.n0 dvss 1.41043f
C3380 por_ana_0.ibias_gen_0.vstart.n1 dvss 0.258324f
C3381 por_ana_0.ibias_gen_0.vstart.t10 dvss 0.344828f
C3382 por_ana_0.ibias_gen_0.vstart.n2 dvss 0.255572f
C3383 por_ana_0.ibias_gen_0.vstart.n3 dvss 0.255572f
C3384 por_ana_0.ibias_gen_0.vstart.n4 dvss 0.398642f
C3385 por_ana_0.ibias_gen_0.vstart.n5 dvss 0.260069f
C3386 por_ana_0.ibias_gen_0.vstart.n6 dvss 0.750761f
C3387 por_ana_0.ibias_gen_0.vstart.n7 dvss 0.255572f
C3388 vin.n0 dvss 0.138413f
C3389 vin.t22 dvss 0.220728f
C3390 vin.t35 dvss 0.236822f
C3391 vin.n1 dvss 0.638413f
C3392 vin.n2 dvss 0.155091f
C3393 vin.t16 dvss 0.104118f
C3394 vin.n3 dvss 0.167086f
C3395 vin.n4 dvss 0.604032f
C3396 vin.n5 dvss 0.3334f
C3397 vin.n6 dvss 0.138413f
C3398 vin.n7 dvss 0.122475f
C3399 vin.t3 dvss 0.104118f
C3400 vin.n8 dvss 0.135924f
C3401 vin.n9 dvss 0.155091f
C3402 vin.t18 dvss 0.104118f
C3403 vin.n10 dvss 0.167086f
C3404 vin.n11 dvss 0.604032f
C3405 vin.n12 dvss 0.155091f
C3406 vin.t15 dvss 0.104118f
C3407 vin.n13 dvss 0.167086f
C3408 vin.n14 dvss 0.604032f
C3409 vin.n15 dvss 0.155091f
C3410 vin.t19 dvss 0.104118f
C3411 vin.n16 dvss 0.167086f
C3412 vin.n17 dvss 0.604032f
C3413 vin.n18 dvss 0.3334f
C3414 vin.n19 dvss 0.296494f
C3415 vin.n20 dvss 0.122475f
C3416 vin.t5 dvss 0.104118f
C3417 vin.n21 dvss 0.135924f
C3418 vin.n22 dvss 0.155091f
C3419 vin.t21 dvss 0.104118f
C3420 vin.n23 dvss 0.167086f
C3421 vin.n24 dvss 0.604032f
C3422 vin.n25 dvss 0.155091f
C3423 vin.t17 dvss 0.104118f
C3424 vin.n26 dvss 0.167086f
C3425 vin.n27 dvss 0.122475f
C3426 vin.n28 dvss 0.3334f
C3427 vin.n29 dvss 0.155091f
C3428 vin.n30 dvss 0.604032f
C3429 vin.n31 dvss 0.167086f
C3430 vin.t20 dvss 0.104118f
C3431 vin.n32 dvss 0.155091f
C3432 vin.n33 dvss 0.604032f
C3433 vin.n34 dvss 0.135924f
C3434 vin.t8 dvss 0.104118f
C3435 vin.n35 dvss 0.122475f
C3436 vin.n36 dvss 0.3334f
C3437 vin.n37 dvss 0.287503f
C3438 vin.n38 dvss 0.218289f
C3439 vin.n39 dvss 0.138413f
C3440 vin.n40 dvss 0.287503f
C3441 vin.n41 dvss 0.135924f
C3442 vin.t9 dvss 0.104118f
C3443 vin.n42 dvss 0.122475f
C3444 vin.n43 dvss 0.3334f
C3445 vin.n44 dvss 0.287503f
C3446 vin.n45 dvss 0.135924f
C3447 vin.t7 dvss 0.104118f
C3448 vin.n46 dvss 0.122475f
C3449 vin.n47 dvss 0.3334f
C3450 vin.n48 dvss 0.287503f
C3451 vin.n49 dvss 0.138413f
C3452 vin.n50 dvss 0.138413f
C3453 vin.n51 dvss 0.287503f
C3454 vin.n52 dvss 0.135924f
C3455 vin.t6 dvss 0.104118f
C3456 vin.n53 dvss 0.122475f
C3457 vin.n54 dvss 0.3334f
C3458 vin.n55 dvss 0.287503f
C3459 vin.n56 dvss 0.135924f
C3460 vin.t4 dvss 0.104118f
C3461 vin.n57 dvss 0.122475f
C3462 vin.n58 dvss 0.3334f
C3463 vin.n59 dvss 0.306818f
C3464 vin.n60 dvss 3.86107f
C3465 vin.n61 dvss 1.22167f
C3466 vin.t64 dvss 1.955f
C3467 vin.t52 dvss 1.7889f
C3468 vin.n62 dvss 1.21671f
C3469 vin.t56 dvss 1.955f
C3470 vin.n65 dvss 1.21671f
C3471 vin.t61 dvss 1.7889f
C3472 vin.n66 dvss 1.21671f
C3473 vin.t63 dvss 1.955f
C3474 vin.n69 dvss 1.21671f
C3475 vin.t51 dvss 1.7889f
C3476 vin.n70 dvss 1.21671f
C3477 vin.t55 dvss 1.955f
C3478 vin.n73 dvss 1.21671f
C3479 vin.t60 dvss 1.7889f
C3480 vin.n74 dvss 1.21671f
C3481 vin.t57 dvss 1.955f
C3482 vin.n77 dvss 1.21671f
C3483 vin.t65 dvss 1.7889f
C3484 vin.n78 dvss 1.21671f
C3485 vin.t54 dvss 1.955f
C3486 vin.n81 dvss 1.21671f
C3487 vin.t59 dvss 1.7889f
C3488 vin.n82 dvss 1.21671f
C3489 vin.t62 dvss 1.955f
C3490 vin.n85 dvss 1.21671f
C3491 vin.t50 dvss 1.7889f
C3492 vin.n86 dvss 1.21671f
C3493 vin.t53 dvss 1.955f
C3494 vin.n89 dvss 1.21671f
C3495 vin.t58 dvss 1.7889f
C3496 vin.n90 dvss 1.21671f
C3497 vin.n91 dvss 0.200089f
C3498 vin.n92 dvss 4.33737f
C3499 vin.n94 dvss 1.03025f
C3500 por_dig_0.net5.n13 dvss 0.195529f
C3501 por_dig_0.net5.n14 dvss 0.307202f
C3502 por_dig_0.net5.n15 dvss 0.225418f
C3503 por_dig_0.net5.n18 dvss 0.379091f
C3504 por_dig_0.net5.n19 dvss 0.398344f
C3505 por_dig_0.net5.n21 dvss 0.215812f
C3506 por_dig_0.net5.n24 dvss 0.336755f
C3507 por_dig_0.clknet_0_osc_ck.n25 dvss 0.228312f
C3508 por_ana_0.rstring_mux_0.vtop.n0 dvss 0.188061f
C3509 por_ana_0.rstring_mux_0.vtop.n1 dvss 0.186982f
C3510 por_ana_0.rstring_mux_0.vtop.n2 dvss 1.02937f
C3511 por_ana_0.rstring_mux_0.vtop.n3 dvss 0.163921f
C3512 por_ana_0.rstring_mux_0.vtop.n4 dvss 0.697228f
C3513 por_ana_0.rstring_mux_0.vtop.n5 dvss 0.262825f
C3514 por_ana_0.rstring_mux_0.vtop.n6 dvss 0.186982f
C3515 por_ana_0.rstring_mux_0.vtop.n7 dvss 0.567273f
C3516 por_ana_0.rstring_mux_0.vtop.n8 dvss 0.186982f
C3517 por_ana_0.rstring_mux_0.vtop.n9 dvss 0.567273f
C3518 por_ana_0.rstring_mux_0.vtop.n10 dvss 0.186982f
C3519 por_ana_0.rstring_mux_0.vtop.n11 dvss 0.567273f
C3520 por_ana_0.rstring_mux_0.vtop.n12 dvss 0.188542f
C3521 por_ana_0.rstring_mux_0.vtop.n13 dvss 0.741617f
C3522 por_ana_0.rstring_mux_0.vtop.n14 dvss 0.163921f
C3523 por_ana_0.rstring_mux_0.vtop.n15 dvss 0.694974f
C3524 por_ana_0.rstring_mux_0.vtop.t17 dvss 2.67225f
C3525 por_dig_0.por_unbuf.n10 dvss 0.104846f
C3526 por_dig_0.por_unbuf.n22 dvss 0.616589f
C3527 por_dig_0.por_unbuf.n27 dvss 0.876778f
C3528 por_dig_0.por_unbuf.n28 dvss 0.989697f
C3529 por_ana_0.schmitt_trigger_0.out.n5 dvss 0.689226f
C3530 por_ana_0.schmitt_trigger_0.out.t12 dvss 0.155689f
C3531 por_ana_0.schmitt_trigger_0.out.t5 dvss 0.155538f
C3532 por_ana_0.schmitt_trigger_0.out.n6 dvss 0.163942f
C3533 por_ana_0.schmitt_trigger_0.out.t4 dvss 0.155622f
C3534 por_ana_0.schmitt_trigger_0.out.n7 dvss 0.113412f
C3535 por_ana_0.schmitt_trigger_0.out.t10 dvss 0.162392f
C3536 por_ana_0.schmitt_trigger_0.out.n8 dvss 0.688643f
C3537 por_ana_0.schmitt_trigger_0.out.n9 dvss 0.41845f
C3538 por_ana_0.schmitt_trigger_0.out.n10 dvss 0.606738f
C3539 por_ana_0.schmitt_trigger_0.out.n11 dvss 0.342028f
C3540 por_dig_0.clknet_1_0__leaf_osc_ck.n18 dvss 0.135513f
C3541 por_dig_0.clknet_1_0__leaf_osc_ck.n30 dvss 0.106117f
C3542 por_dig_0.clknet_1_0__leaf_osc_ck.n40 dvss 0.257698f
C3543 por_dig_0.clknet_1_0__leaf_osc_ck.n41 dvss 0.231497f
C3544 por_dig_0.clknet_1_0__leaf_osc_ck.n42 dvss 0.263956f
C3545 por_dig_0.clknet_1_0__leaf_osc_ck.n46 dvss 0.249567f
C3546 por_dig_0.clknet_1_0__leaf_osc_ck.n50 dvss 0.261802f
C3547 por_dig_0.clknet_1_0__leaf_osc_ck.n51 dvss 0.21642f
C3548 por_dig_0.clknet_1_0__leaf_osc_ck.n54 dvss 0.207182f
C3549 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n0 dvss 1.20316f
C3550 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n1 dvss 0.160523f
C3551 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n2 dvss 0.178108f
C3552 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n3 dvss 0.211986f
C3553 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n5 dvss 0.211924f
C3554 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n6 dvss 0.211986f
C3555 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n7 dvss 0.211924f
C3556 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n8 dvss 0.211986f
C3557 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n10 dvss 0.211924f
C3558 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n11 dvss 0.211986f
C3559 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n12 dvss 0.211924f
C3560 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n13 dvss 0.211986f
C3561 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n15 dvss 0.211924f
C3562 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n16 dvss 0.194362f
C3563 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n17 dvss 0.211979f
C3564 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n18 dvss 0.400799f
C3565 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n20 dvss 0.600313f
C3566 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n21 dvss 0.500556f
C3567 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n26 dvss 0.250062f
C3568 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.t20 dvss 0.175854f
C3569 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.t16 dvss 0.175854f
C3570 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.t24 dvss 0.175854f
C3571 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.t11 dvss 0.175854f
C3572 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.t14 dvss 0.175854f
C3573 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.t13 dvss 0.175854f
C3574 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.t8 dvss 0.175854f
C3575 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.t37 dvss 0.175854f
C3576 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.t28 dvss 0.175854f
C3577 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.t39 dvss 0.184266f
C3578 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n27 dvss 0.196778f
C3579 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.t18 dvss 0.175854f
C3580 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.t19 dvss 0.175854f
C3581 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.t12 dvss 0.175854f
C3582 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.t15 dvss 0.175854f
C3583 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.t21 dvss 0.175854f
C3584 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.t22 dvss 0.19333f
C3585 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n30 dvss 0.188483f
C3586 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n35 dvss 0.166326f
C3587 por_ana_0.sky130_fd_sc_hvl__inv_16_0.A.n37 dvss 0.288952f
C3588 pwup_filt.n17 dvss 0.455046f
C3589 pwup_filt.n18 dvss 1.93487f
C3590 por_dig_0.cnt_por\[0\].n9 dvss 0.154942f
C3591 por_dig_0.cnt_por\[0\].n14 dvss 0.191777f
C3592 por_dig_0.cnt_por\[0\].n19 dvss 0.136753f
C3593 por_dig_0.cnt_por\[0\].n21 dvss 0.109641f
C3594 por_dig_0.cnt_por\[0\].n27 dvss 0.134021f
C3595 por_dig_0.cnt_por\[0\].n28 dvss 0.122413f
C3596 por_dig_0.cnt_por\[0\].n29 dvss 0.19557f
C3597 por_ana_0.comparator_0.vinn.n0 dvss 0.589592f
C3598 por_ana_0.comparator_0.vinn.n1 dvss 0.589592f
C3599 por_ana_0.comparator_0.vinn.n2 dvss 0.589592f
C3600 por_ana_0.comparator_0.vinn.n3 dvss 0.589592f
C3601 por_ana_0.comparator_0.vinn.n4 dvss 0.589592f
C3602 por_ana_0.comparator_0.vinn.n5 dvss 0.59813f
C3603 por_ana_0.comparator_0.vinn.n6 dvss 0.61612f
C3604 por_ana_0.comparator_0.vinn.n7 dvss 0.589592f
C3605 por_ana_0.comparator_0.vinn.n8 dvss 0.15866f
C3606 por_ana_0.comparator_0.vinn.n9 dvss 0.12907f
C3607 por_ana_0.comparator_0.vinn.n10 dvss 0.116299f
C3608 por_ana_0.comparator_0.vinn.n11 dvss 0.12907f
C3609 por_ana_0.comparator_0.vinn.t46 dvss 0.214071f
C3610 por_ana_0.comparator_0.vinn.n12 dvss 0.605638f
C3611 por_ana_0.comparator_0.vinn.t27 dvss 0.197177f
C3612 por_ana_0.comparator_0.vinn.n13 dvss 0.116299f
C3613 por_ana_0.comparator_0.vinn.n14 dvss 0.12907f
C3614 por_ana_0.comparator_0.vinn.n15 dvss 0.207281f
C3615 por_ana_0.comparator_0.vinn.n16 dvss 0.116299f
C3616 por_ana_0.comparator_0.vinn.n17 dvss 0.12907f
C3617 por_ana_0.comparator_0.vinn.n18 dvss 0.131433f
C3618 por_ana_0.comparator_0.vinn.n19 dvss 0.116299f
C3619 por_ana_0.comparator_0.vinn.n20 dvss 0.12907f
C3620 por_ana_0.comparator_0.vinn.n21 dvss 0.131433f
C3621 por_ana_0.comparator_0.vinn.n22 dvss 0.116299f
C3622 por_ana_0.comparator_0.vinn.n23 dvss 0.12907f
C3623 por_ana_0.comparator_0.vinn.n24 dvss 0.131433f
C3624 por_ana_0.comparator_0.vinn.n25 dvss 0.116299f
C3625 por_ana_0.comparator_0.vinn.n26 dvss 0.12907f
C3626 por_ana_0.comparator_0.vinn.n27 dvss 0.131433f
C3627 por_ana_0.comparator_0.vinn.n28 dvss 0.207281f
C3628 por_ana_0.comparator_0.vinn.n29 dvss 0.12907f
C3629 por_ana_0.comparator_0.vinn.n30 dvss 0.116299f
C3630 por_ana_0.comparator_0.vinn.n31 dvss 0.15754f
C3631 por_ana_0.comparator_0.vinn.t49 dvss 2.07788f
C3632 por_ana_0.comparator_0.vinn.t55 dvss 1.98852f
C3633 por_ana_0.comparator_0.vinn.n32 dvss 1.65591f
C3634 por_ana_0.comparator_0.vinn.t63 dvss 1.98852f
C3635 por_ana_0.comparator_0.vinn.n33 dvss 0.874582f
C3636 por_ana_0.comparator_0.vinn.t54 dvss 1.98852f
C3637 por_ana_0.comparator_0.vinn.n34 dvss 0.874582f
C3638 por_ana_0.comparator_0.vinn.t62 dvss 1.98852f
C3639 por_ana_0.comparator_0.vinn.n35 dvss 0.874582f
C3640 por_ana_0.comparator_0.vinn.t48 dvss 1.98852f
C3641 por_ana_0.comparator_0.vinn.n36 dvss 0.874582f
C3642 por_ana_0.comparator_0.vinn.t53 dvss 1.98852f
C3643 por_ana_0.comparator_0.vinn.n37 dvss 0.874582f
C3644 por_ana_0.comparator_0.vinn.t59 dvss 1.98852f
C3645 por_ana_0.comparator_0.vinn.n38 dvss 1.03441f
C3646 por_ana_0.comparator_0.vinn.t57 dvss 2.09565f
C3647 por_ana_0.comparator_0.vinn.t61 dvss 2.00504f
C3648 por_ana_0.comparator_0.vinn.n39 dvss 1.69313f
C3649 por_ana_0.comparator_0.vinn.t52 dvss 2.00504f
C3650 por_ana_0.comparator_0.vinn.n40 dvss 0.893824f
C3651 por_ana_0.comparator_0.vinn.t60 dvss 2.00504f
C3652 por_ana_0.comparator_0.vinn.n41 dvss 0.893824f
C3653 por_ana_0.comparator_0.vinn.t51 dvss 2.00504f
C3654 por_ana_0.comparator_0.vinn.n42 dvss 0.893824f
C3655 por_ana_0.comparator_0.vinn.t56 dvss 2.00504f
C3656 por_ana_0.comparator_0.vinn.n43 dvss 0.893824f
C3657 por_ana_0.comparator_0.vinn.t58 dvss 2.00504f
C3658 por_ana_0.comparator_0.vinn.n44 dvss 0.893824f
C3659 por_ana_0.comparator_0.vinn.t50 dvss 2.00504f
C3660 por_ana_0.comparator_0.vinn.n45 dvss 0.98848f
C3661 por_ana_0.comparator_0.vinn.n46 dvss 3.52107f
C3662 por_ana_0.comparator_0.vinn.n47 dvss 3.48273f
C3663 por_ana_0.comparator_0.vinn.n48 dvss 0.29169f
C3664 por_ana_0.comparator_0.vinn.n49 dvss 0.14727f
C3665 por_ana_0.comparator_0.vinn.n50 dvss 0.15866f
C3666 por_ana_0.comparator_0.vinn.n51 dvss 0.573572f
C3667 por_ana_0.comparator_0.vinn.n52 dvss 0.14727f
C3668 por_ana_0.comparator_0.vinn.n53 dvss 0.15866f
C3669 por_ana_0.comparator_0.vinn.n54 dvss 0.573572f
C3670 por_ana_0.comparator_0.vinn.n55 dvss 0.14727f
C3671 por_ana_0.comparator_0.vinn.n56 dvss 0.15866f
C3672 por_ana_0.comparator_0.vinn.n57 dvss 0.573572f
C3673 por_ana_0.comparator_0.vinn.n58 dvss 0.14727f
C3674 por_ana_0.comparator_0.vinn.n59 dvss 0.15866f
C3675 por_ana_0.comparator_0.vinn.n60 dvss 0.573572f
C3676 por_ana_0.comparator_0.vinn.n61 dvss 0.14727f
C3677 por_ana_0.comparator_0.vinn.n62 dvss 0.15866f
C3678 por_ana_0.comparator_0.vinn.n63 dvss 0.573572f
C3679 por_ana_0.comparator_0.vinn.n64 dvss 0.14727f
C3680 por_ana_0.comparator_0.vinn.n65 dvss 0.15866f
C3681 por_ana_0.comparator_0.vinn.n66 dvss 0.573572f
C3682 por_ana_0.comparator_0.vinn.n67 dvss 0.14727f
C3683 por_ana_0.comparator_0.vnn.n0 dvss 1.16602f
C3684 por_ana_0.comparator_0.vnn.n1 dvss 5.1835f
C3685 por_ana_0.comparator_0.vnn.n2 dvss 1.03415f
C3686 por_ana_0.comparator_0.vnn.n3 dvss 1.03415f
C3687 por_ana_0.comparator_0.vnn.n4 dvss 1.03415f
C3688 por_ana_0.comparator_0.vnn.n5 dvss 1.03415f
C3689 por_ana_0.comparator_0.vnn.n6 dvss 5.5579f
C3690 por_ana_0.comparator_0.vnn.n7 dvss 3.16283f
C3691 por_ana_0.comparator_0.vnn.t35 dvss 1.39949f
C3692 por_ana_0.comparator_0.vnn.t39 dvss 1.39949f
C3693 por_ana_0.comparator_0.vnn.t37 dvss 1.39949f
C3694 por_ana_0.comparator_0.vnn.t41 dvss 1.39949f
C3695 por_ana_0.comparator_0.vnn.t43 dvss 1.39949f
C3696 por_ana_0.comparator_0.vnn.t45 dvss 1.39949f
C3697 por_ana_0.comparator_0.vnn.t31 dvss 1.39949f
C3698 por_ana_0.comparator_0.vnn.t33 dvss 1.39949f
C3699 por_ana_0.comparator_0.vnn.t54 dvss 1.49452f
C3700 por_ana_0.comparator_0.vnn.t48 dvss 1.29454f
C3701 por_ana_0.comparator_0.vnn.t56 dvss 1.49452f
C3702 por_ana_0.comparator_0.vnn.t50 dvss 1.29454f
C3703 por_ana_0.comparator_0.vnn.t55 dvss 1.49452f
C3704 por_ana_0.comparator_0.vnn.t49 dvss 1.29454f
C3705 por_ana_0.comparator_0.vnn.t62 dvss 1.49452f
C3706 por_ana_0.comparator_0.vnn.t58 dvss 1.29454f
C3707 por_ana_0.comparator_0.vnn.t57 dvss 1.49452f
C3708 por_ana_0.comparator_0.vnn.t53 dvss 1.29454f
C3709 por_ana_0.comparator_0.vnn.t51 dvss 1.49452f
C3710 por_ana_0.comparator_0.vnn.t59 dvss 1.29454f
C3711 por_ana_0.comparator_0.vnn.t52 dvss 1.49452f
C3712 por_ana_0.comparator_0.vnn.t60 dvss 1.29454f
C3713 por_ana_0.comparator_0.vnn.t61 dvss 1.49452f
C3714 por_ana_0.comparator_0.vnn.t47 dvss 1.29454f
C3715 por_ana_0.schmitt_trigger_0.m.n2 dvss 0.65613f
C3716 por_ana_0.schmitt_trigger_0.m.n4 dvss 0.195435f
C3717 por_ana_0.schmitt_trigger_0.m.t15 dvss 0.161114f
C3718 por_ana_0.schmitt_trigger_0.m.t17 dvss 0.164304f
C3719 por_ana_0.schmitt_trigger_0.m.t16 dvss 0.16415f
C3720 por_ana_0.schmitt_trigger_0.m.n5 dvss 0.16975f
C3721 por_ana_0.schmitt_trigger_0.m.t14 dvss 0.16428f
C3722 por_ana_0.schmitt_trigger_0.m.n6 dvss 0.3748f
C3723 por_ana_0.schmitt_trigger_0.m.n7 dvss 0.537335f
C3724 por_ana_0.schmitt_trigger_0.m.n10 dvss 0.732652f
C3725 por_ana_0.schmitt_trigger_0.m.n11 dvss 0.312554f
C3726 por_ana_0.schmitt_trigger_0.m.n13 dvss 0.192206f
C3727 por_ana_0.schmitt_trigger_0.m.n15 dvss 0.222965f
C3728 por_ana_0.schmitt_trigger_0.in.t6 dvss 2.51822f
C3729 por_ana_0.schmitt_trigger_0.in.t14 dvss 1.35606f
C3730 por_ana_0.schmitt_trigger_0.in.n5 dvss 1.52632f
C3731 por_ana_0.schmitt_trigger_0.in.t8 dvss 1.35606f
C3732 por_ana_0.schmitt_trigger_0.in.n6 dvss 1.34684f
C3733 por_ana_0.schmitt_trigger_0.in.t7 dvss 1.35606f
C3734 por_ana_0.schmitt_trigger_0.in.n7 dvss 1.34684f
C3735 por_ana_0.schmitt_trigger_0.in.t13 dvss 1.35606f
C3736 por_ana_0.schmitt_trigger_0.in.n8 dvss 1.34684f
C3737 por_ana_0.schmitt_trigger_0.in.t10 dvss 1.35606f
C3738 por_ana_0.schmitt_trigger_0.in.n9 dvss 1.43721f
C3739 por_ana_0.rstring_mux_0.vtrip6.t0 dvss 0.775728f
C3740 por_ana_0.rstring_mux_0.vtrip6.n0 dvss 0.187027f
C3741 por_ana_0.rstring_mux_0.vtrip6.n1 dvss 0.122626f
C3742 por_ana_0.rstring_mux_0.vtrip6.n2 dvss 0.800766f
C3743 por_ana_0.rstring_mux_0.vtrip6.n3 dvss 0.187027f
C3744 por_ana_0.rstring_mux_0.vtrip6.n4 dvss 0.122626f
C3745 por_ana_0.rstring_mux_0.vtrip6.n5 dvss 1.249f
C3746 por_ana_0.rstring_mux_0.vtrip6.n6 dvss 1.9489f
C3747 por_ana_0.rstring_mux_0.vtrip6.n7 dvss 1.58785f
C3748 por_ana_0.rstring_mux_0.vtrip6.t5 dvss 0.166356f
C3749 por_ana_0.rstring_mux_0.vtrip5.t1 dvss 0.169149f
C3750 por_ana_0.rstring_mux_0.vtrip5.n0 dvss 0.183575f
C3751 por_ana_0.rstring_mux_0.vtrip5.n1 dvss 0.120363f
C3752 por_ana_0.rstring_mux_0.vtrip5.n2 dvss 1.20735f
C3753 por_ana_0.rstring_mux_0.vtrip5.n3 dvss 0.183575f
C3754 por_ana_0.rstring_mux_0.vtrip5.n4 dvss 0.120363f
C3755 por_ana_0.rstring_mux_0.vtrip5.n5 dvss 0.742428f
C3756 por_ana_0.rstring_mux_0.vtrip5.n6 dvss 0.936052f
C3757 por_ana_0.rstring_mux_0.vtrip5.n7 dvss 2.7123f
C3758 por_ana_0.rstring_mux_0.vtrip5.t0 dvss 0.169167f
C3759 por_dig_0.net7.n0 dvss 0.642722f
C3760 por_dig_0.net7.n10 dvss 0.231554f
C3761 por_dig_0.net7.n17 dvss 0.396583f
C3762 por_dig_0.net7.n20 dvss 0.286976f
C3763 por_ana_0.ibias_gen_0.ibias0.n0 dvss 3.82913f
C3764 por_ana_0.ibias_gen_0.ibias0.n1 dvss 0.899038f
C3765 por_ana_0.ibias_gen_0.vp.n0 dvss 0.431943f
C3766 por_ana_0.ibias_gen_0.vp.t6 dvss 0.188332f
C3767 por_ana_0.ibias_gen_0.vp.n3 dvss 0.662608f
C3768 por_ana_0.ibias_gen_0.vp.t8 dvss 1.71268f
C3769 por_ana_0.ibias_gen_0.vp.n4 dvss 1.29098f
C3770 por_ana_0.ibias_gen_0.vp.t7 dvss 1.65245f
C3771 por_ana_0.ibias_gen_0.vp.n5 dvss 1.29098f
C3772 por_ana_0.ibias_gen_0.vp.t10 dvss 1.65245f
C3773 por_ana_0.ibias_gen_0.vp.n6 dvss 1.29098f
C3774 por_ana_0.ibias_gen_0.vp.t11 dvss 1.68256f
C3775 por_ana_0.ibias_gen_0.vp.n7 dvss 0.597984f
C3776 por_ana_0.ibias_gen_0.vp.t12 dvss 2.31092f
C3777 por_ana_0.ibias_gen_0.vp.t9 dvss 2.34104f
C3778 por_ana_0.ibias_gen_0.vp.n8 dvss 0.730243f
C3779 por_ana_0.ibias_gen_0.vp.n9 dvss 1.1851f
C3780 por_ana_0.ibias_gen_0.vp.n10 dvss 0.917156f
C3781 por_ana_0.ibias_gen_0.vp.n12 dvss 0.488746f
C3782 por_dig_0._034_.n8 dvss 0.174295f
C3783 por_dig_0._034_.n11 dvss 0.294368f
C3784 por_dig_0._034_.n14 dvss 0.158565f
C3785 por_ana_0.sky130_fd_sc_hvl__lsbuflv2hv_1_0[0|7].X dvss 0.106163f
C3786 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[6].t3 dvss 0.27812f
C3787 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[6].t4 dvss 0.278015f
C3788 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[6].n2 dvss 0.268193f
C3789 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[6].n5 dvss 1.26254f
C3790 por_ana_0.rstring_mux_0.vtrip_decoded_avdd[6].n6 dvss 0.65885f
C3791 por_ana_0.rstring_mux_0.vtrip2.t5 dvss 0.211519f
C3792 por_ana_0.rstring_mux_0.vtrip2.n0 dvss 0.229108f
C3793 por_ana_0.rstring_mux_0.vtrip2.n1 dvss 0.150216f
C3794 por_ana_0.rstring_mux_0.vtrip2.n2 dvss 0.947831f
C3795 por_ana_0.rstring_mux_0.vtrip2.n3 dvss 0.229108f
C3796 por_ana_0.rstring_mux_0.vtrip2.n4 dvss 0.150216f
C3797 por_ana_0.rstring_mux_0.vtrip2.n5 dvss 1.50485f
C3798 por_ana_0.rstring_mux_0.vtrip2.n6 dvss 2.43692f
C3799 por_ana_0.rstring_mux_0.vtrip2.n7 dvss 2.81264f
C3800 por_ana_0.rstring_mux_0.vtrip2.t2 dvss 0.898141f
C3801 por_ana_0.rstring_mux_0.vtrip3.t9 dvss 0.157727f
C3802 por_ana_0.rstring_mux_0.vtrip3.n0 dvss 0.17118f
C3803 por_ana_0.rstring_mux_0.vtrip3.n1 dvss 0.112235f
C3804 por_ana_0.rstring_mux_0.vtrip3.n2 dvss 0.753957f
C3805 por_ana_0.rstring_mux_0.vtrip3.n3 dvss 0.17118f
C3806 por_ana_0.rstring_mux_0.vtrip3.n4 dvss 0.112235f
C3807 por_ana_0.rstring_mux_0.vtrip3.n5 dvss 1.08769f
C3808 por_ana_0.rstring_mux_0.vtrip3.n6 dvss 0.877189f
C3809 por_ana_0.rstring_mux_0.vtrip3.n7 dvss 2.47396f
C3810 por_ana_0.rstring_mux_0.vtrip3.t4 dvss 0.157744f
C3811 dcomp.n30 dvss 0.585628f
C3812 por_ana_0.comparator_1.vpp.n0 dvss 5.51282f
C3813 por_ana_0.comparator_1.vpp.n1 dvss 4.2909f
C3814 por_ana_0.comparator_1.vpp.n2 dvss 8.02316f
C3815 por_ana_0.comparator_1.vpp.n3 dvss 1.27207f
C3816 por_ana_0.comparator_1.vpp.n4 dvss 1.27207f
C3817 por_ana_0.comparator_1.vpp.t10 dvss 1.40408f
C3818 por_ana_0.comparator_1.vpp.t6 dvss 1.40408f
C3819 por_ana_0.comparator_1.vpp.t4 dvss 1.40408f
C3820 por_ana_0.comparator_1.vpp.t0 dvss 1.40408f
C3821 por_ana_0.comparator_1.vpp.t12 dvss 1.40408f
C3822 por_ana_0.comparator_1.vpp.t8 dvss 1.40408f
C3823 por_ana_0.comparator_1.vpp.t2 dvss 1.40408f
C3824 por_ana_0.comparator_1.vpp.t14 dvss 1.40408f
C3825 por_ana_0.comparator_1.vpp.t62 dvss 1.49278f
C3826 por_ana_0.comparator_1.vpp.t48 dvss 1.30445f
C3827 por_ana_0.comparator_1.vpp.t50 dvss 1.49278f
C3828 por_ana_0.comparator_1.vpp.t55 dvss 1.30445f
C3829 por_ana_0.comparator_1.vpp.t51 dvss 1.49278f
C3830 por_ana_0.comparator_1.vpp.t56 dvss 1.30445f
C3831 por_ana_0.comparator_1.vpp.t52 dvss 1.49278f
C3832 por_ana_0.comparator_1.vpp.t57 dvss 1.30445f
C3833 por_ana_0.comparator_1.vpp.t53 dvss 1.49278f
C3834 por_ana_0.comparator_1.vpp.t58 dvss 1.30445f
C3835 por_ana_0.comparator_1.vpp.t60 dvss 1.49278f
C3836 por_ana_0.comparator_1.vpp.t61 dvss 1.30445f
C3837 por_ana_0.comparator_1.vpp.t54 dvss 1.49278f
C3838 por_ana_0.comparator_1.vpp.t59 dvss 1.30445f
C3839 por_ana_0.comparator_1.vpp.t47 dvss 1.49278f
C3840 por_ana_0.comparator_1.vpp.t49 dvss 1.30445f
C3841 por_dig_0.net23.n0 dvss 0.126275f
C3842 por_dig_0.net23.n7 dvss 0.170246f
C3843 por_dig_0.net23.n18 dvss 0.13607f
C3844 por_dig_0.net23.n23 dvss 0.154766f
C3845 por_dig_0.net23.n27 dvss 0.162338f
C3846 por_dig_0.net23.n28 dvss 0.129169f
C3847 osc_ck.n8 dvss 0.658829f
C3848 osc_ck.n9 dvss 0.434689f
C3849 osc_ck.n10 dvss 0.248882f
C3850 osc_ck.n11 dvss 3.52702f
C3851 osc_ck.n12 dvss 4.83809f
C3852 por.n30 dvss 0.566272f
C3853 avss.n1 dvss 0.63981f
C3854 avss.n7 dvss 2.65437f
C3855 avss.t156 dvss 6.89451f
C3856 avss.n8 dvss 7.70488f
C3857 avss.t364 dvss 6.60459f
C3858 avss.n9 dvss 0.206188f
C3859 avss.n10 dvss 0.206188f
C3860 avss.n11 dvss 0.289882f
C3861 avss.t34 dvss 0.455506f
C3862 avss.t165 dvss 6.60459f
C3863 avss.t234 dvss 9.11583f
C3864 avss.n12 dvss 0.294077f
C3865 avss.n13 dvss 0.294077f
C3866 avss.n14 dvss 0.172673f
C3867 avss.n15 dvss 0.143772f
C3868 avss.t339 dvss 0.216947f
C3869 avss.t383 dvss 0.212474f
C3870 avss.n16 dvss 0.865895f
C3871 avss.n17 dvss 0.204678f
C3872 avss.t341 dvss 9.492519f
C3873 avss.t244 dvss 11.5015f
C3874 avss.t323 dvss 9.492519f
C3875 avss.t163 dvss 5.75076f
C3876 avss.n18 dvss 9.492519f
C3877 avss.t218 dvss 5.75076f
C3878 avss.t325 dvss 9.492519f
C3879 avss.t248 dvss 9.46741f
C3880 avss.t396 dvss 3.46552f
C3881 avss.t335 dvss 8.06111f
C3882 avss.t305 dvss 9.11583f
C3883 avss.t217 dvss 5.47452f
C3884 avss.n19 dvss 0.394198f
C3885 avss.n20 dvss 0.394198f
C3886 avss.n21 dvss 0.231601f
C3887 avss.n22 dvss 0.12851f
C3888 avss.t97 dvss 0.348381f
C3889 avss.n23 dvss 0.341542f
C3890 avss.t70 dvss 0.3484f
C3891 avss.n24 dvss 0.296013f
C3892 avss.t39 dvss 0.348384f
C3893 avss.n25 dvss 0.645131f
C3894 avss.n26 dvss 2.02224f
C3895 avss.n27 dvss 1.02499f
C3896 avss.t105 dvss 4.08169f
C3897 avss.t107 dvss 0.15847f
C3898 avss.n28 dvss 1.54091f
C3899 avss.n29 dvss 0.399913f
C3900 avss.n30 dvss 0.638189f
C3901 avss.n31 dvss 0.150542f
C3902 avss.n32 dvss 0.162702f
C3903 avss.n33 dvss 1.25073f
C3904 avss.n34 dvss 1.25073f
C3905 avss.t57 dvss 4.08169f
C3906 avss.n35 dvss 0.162702f
C3907 avss.t58 dvss 0.200808f
C3908 avss.n36 dvss 1.54091f
C3909 avss.n37 dvss 0.457138f
C3910 avss.n38 dvss 0.450301f
C3911 avss.n40 dvss 0.920493f
C3912 avss.t115 dvss 4.08169f
C3913 avss.t117 dvss 0.15847f
C3914 avss.n41 dvss 1.54091f
C3915 avss.n42 dvss 0.399913f
C3916 avss.n44 dvss 0.690062f
C3917 avss.n45 dvss 0.690062f
C3918 avss.t338 dvss 2.05922f
C3919 avss.t382 dvss 9.492519f
C3920 avss.t319 dvss 6.47902f
C3921 avss.t35 dvss 7.4333f
C3922 avss.n46 dvss 6.47902f
C3923 avss.n47 dvss 1.08831f
C3924 avss.n48 dvss 1.08831f
C3925 avss.n49 dvss 8.259799f
C3926 avss.t337 dvss 4.84671f
C3927 avss.n50 dvss 1.71896f
C3928 avss.n51 dvss 1.71896f
C3929 avss.n52 dvss 1.71896f
C3930 avss.n53 dvss 2.73003f
C3931 avss.n54 dvss 1.72077f
C3932 avss.n55 dvss 0.606218f
C3933 avss.n56 dvss 3.82626f
C3934 avss.n57 dvss 0.834494f
C3935 avss.n58 dvss 0.403922f
C3936 avss.n59 dvss 0.96103f
C3937 avss.n60 dvss 0.786686f
C3938 avss.n61 dvss 0.781665f
C3939 avss.n62 dvss 0.781665f
C3940 avss.t81 dvss 0.148617p
C3941 avss.t27 dvss 16.2904f
C3942 avss.n63 dvss 3.28517f
C3943 avss.n64 dvss 29.959698f
C3944 avss.t104 dvss 1.06784f
C3945 avss.n65 dvss 0.206718f
C3946 avss.n66 dvss 0.206718f
C3947 avss.t298 dvss 5.55172f
C3948 avss.t40 dvss 5.04761f
C3949 avss.n69 dvss 1.89088f
C3950 avss.n70 dvss 11.654901f
C3951 avss.n71 dvss 37.1594f
C3952 avss.n72 dvss 0.943753f
C3953 avss.n73 dvss 0.943753f
C3954 avss.n74 dvss 0.570582f
C3955 avss.n75 dvss 0.623434f
C3956 avss.n76 dvss 0.61967f
C3957 avss.n77 dvss 1.09967f
C3958 avss.t331 dvss 1.13458f
C3959 avss.n78 dvss 0.96003f
C3960 avss.t276 dvss 3.60835f
C3961 avss.t42 dvss 0.791536f
C3962 avss.n79 dvss 3.31379f
C3963 avss.t280 dvss 0.232692f
C3964 avss.t268 dvss 0.376292f
C3965 avss.t272 dvss 0.376292f
C3966 avss.t278 dvss 0.656996f
C3967 avss.n80 dvss 0.512839f
C3968 avss.n81 dvss 0.220653f
C3969 avss.n82 dvss 0.104352f
C3970 avss.n83 dvss 0.108871f
C3971 avss.n85 dvss 0.202626f
C3972 avss.n89 dvss 0.203153f
C3973 avss.n91 dvss 0.11116f
C3974 avss.n93 dvss 0.198518f
C3975 avss.n95 dvss 0.134943f
C3976 avss.n99 dvss 2.15301f
C3977 avss.n101 dvss 0.262183f
C3978 avss.n102 dvss 0.468516f
C3979 avss.t95 dvss 1.11293f
C3980 avss.n103 dvss 5.56155f
C3981 avss.t44 dvss 1.11293f
C3982 avss.n104 dvss 0.551361f
C3983 avss.n106 dvss 0.468516f
C3984 avss.n108 dvss 0.134943f
C3985 avss.n110 dvss 0.124609f
C3986 avss.n111 dvss 0.467264f
C3987 avss.n112 dvss 31.0235f
C3988 avss.n113 dvss 1.08437f
C3989 avss.n114 dvss 0.148681f
C3990 avss.n115 dvss 0.214704f
C3991 avss.n116 dvss 0.112866f
C3992 avss.n117 dvss 0.250147f
C3993 avss.n118 dvss 0.839556f
C3994 avss.n119 dvss 0.13071f
C3995 avss.n120 dvss 0.839556f
C3996 avss.t320 dvss 3.37711f
C3997 avss.n132 dvss 0.212772f
C3998 avss.t385 dvss 0.267958f
C3999 avss.n133 dvss 1.72077f
C4000 avss.n134 dvss 54.083897f
C4001 avss.t166 dvss 9.57101f
C4002 avss.t409 dvss 11.4489f
C4003 avss.t245 dvss 11.4489f
C4004 avss.t353 dvss 11.4489f
C4005 avss.t177 dvss 11.3429f
C4006 avss.t309 dvss 5.42155f
C4007 avss.t310 dvss 2.99851f
C4008 avss.t173 dvss 2.69563f
C4009 avss.t73 dvss 5.08838f
C4010 avss.t30 dvss 3.33168f
C4011 avss.t155 dvss 2.69563f
C4012 avss.t31 dvss 4.75522f
C4013 avss.t87 dvss 3.66485f
C4014 avss.t242 dvss 2.69563f
C4015 avss.t5 dvss 2.86221f
C4016 avss.n135 dvss 2.69563f
C4017 avss.t2 dvss 2.86221f
C4018 avss.t214 dvss 2.69563f
C4019 avss.t51 dvss 4.08888f
C4020 avss.t238 dvss 4.33118f
C4021 avss.t287 dvss 2.69563f
C4022 avss.t237 dvss 3.75571f
C4023 avss.t109 dvss 4.66435f
C4024 avss.t149 dvss 2.69563f
C4025 avss.t378 dvss 3.42254f
C4026 avss.t379 dvss 4.99752f
C4027 avss.t367 dvss 2.69563f
C4028 avss.t123 dvss 3.08938f
C4029 avss.t259 dvss 5.33069f
C4030 avss.t160 dvss 2.69563f
C4031 avss.t260 dvss 2.75621f
C4032 avss.t79 dvss 5.39126f
C4033 avss.t373 dvss 2.96822f
C4034 avss.t0 dvss 2.69563f
C4035 avss.t374 dvss 5.11867f
C4036 avss.t114 dvss 3.30139f
C4037 avss.t360 dvss 2.69563f
C4038 avss.t229 dvss 4.7855f
C4039 avss.t226 dvss 3.63456f
C4040 avss.t312 dvss 2.69563f
C4041 avss.t60 dvss 4.45234f
C4042 avss.t221 dvss 3.96773f
C4043 avss.t286 dvss 2.69563f
C4044 avss.t222 dvss 4.11917f
C4045 avss.t94 dvss 4.3009f
C4046 avss.t361 dvss 2.69563f
C4047 avss.t315 dvss 3.786f
C4048 avss.t316 dvss 4.63406f
C4049 avss.t241 dvss 2.69563f
C4050 avss.t121 dvss 3.45283f
C4051 avss.t265 dvss 4.96723f
C4052 avss.t267 dvss 2.69563f
C4053 avss.t266 dvss 3.11966f
C4054 avss.t125 dvss 5.3004f
C4055 avss.t170 dvss 2.69563f
C4056 avss.t6 dvss 2.7865f
C4057 avss.t7 dvss 5.39126f
C4058 avss.t85 dvss 2.93794f
C4059 avss.t1 dvss 2.69563f
C4060 avss.t328 dvss 5.14896f
C4061 avss.t327 dvss 3.2711f
C4062 avss.t366 dvss 2.69563f
C4063 avss.t49 dvss 4.81579f
C4064 avss.t302 dvss 3.60427f
C4065 avss.t171 dvss 2.69563f
C4066 avss.t303 dvss 4.48262f
C4067 avss.t62 dvss 3.93744f
C4068 avss.t284 dvss 2.69563f
C4069 avss.t211 dvss 4.14946f
C4070 avss.t210 dvss 4.27061f
C4071 avss.t172 dvss 2.69563f
C4072 avss.t135 dvss 3.81629f
C4073 avss.t393 dvss 4.60378f
C4074 avss.t311 dvss 2.69563f
C4075 avss.t392 dvss 4.1646f
C4076 avss.t48 dvss 0.309333f
C4077 avss.t78 dvss 0.309333f
C4078 avss.t72 dvss 0.30935f
C4079 avss.n136 dvss 0.198885f
C4080 avss.t86 dvss 0.30935f
C4081 avss.n137 dvss 0.18977f
C4082 avss.t50 dvss 0.30935f
C4083 avss.n138 dvss 0.18977f
C4084 avss.t108 dvss 0.30935f
C4085 avss.n139 dvss 0.18977f
C4086 avss.t122 dvss 0.30935f
C4087 avss.n140 dvss 0.191982f
C4088 avss.n141 dvss 0.185132f
C4089 avss.t113 dvss 0.30935f
C4090 avss.n142 dvss 0.189053f
C4091 avss.t59 dvss 0.30935f
C4092 avss.n144 dvss 0.154279f
C4093 avss.t93 dvss 0.30935f
C4094 avss.n145 dvss 0.190139f
C4095 avss.t120 dvss 0.30935f
C4096 avss.n146 dvss 0.189902f
C4097 avss.t124 dvss 0.30935f
C4098 avss.n147 dvss 0.18977f
C4099 avss.t84 dvss 0.30935f
C4100 avss.n148 dvss 0.191982f
C4101 avss.n149 dvss 0.185161f
C4102 avss.t61 dvss 0.30935f
C4103 avss.n150 dvss 0.191932f
C4104 avss.t134 dvss 0.30935f
C4105 avss.n151 dvss 0.198092f
C4106 avss.n153 dvss 0.223929f
C4107 avss.n154 dvss 0.255905f
C4108 avss.n156 dvss 0.846866f
C4109 avss.n157 dvss 4.93694f
C4110 avss.t285 dvss 7.28426f
C4111 avss.t246 dvss 11.4489f
C4112 avss.t355 dvss 11.4489f
C4113 avss.t236 dvss 11.4489f
C4114 avss.t154 dvss 11.4489f
C4115 avss.t357 dvss 11.4489f
C4116 avss.t26 dvss 11.4489f
C4117 avss.t249 dvss 11.4489f
C4118 avss.t169 dvss 11.4489f
C4119 avss.t225 dvss 11.4489f
C4120 avss.t250 dvss 5.83044f
C4121 avss.n158 dvss 67.083496f
C4122 avss.n159 dvss 39.955f
C4123 avss.n208 dvss 0.797364f
C4124 avss.n211 dvss 0.624262f
C4125 avss.n219 dvss 0.331238f
C4126 avss.n220 dvss 0.325944f
C4127 avss.n231 dvss 0.331238f
C4128 avss.n232 dvss 0.325944f
C4129 avss.n243 dvss 0.331238f
C4130 avss.n244 dvss 0.325944f
C4131 avss.n255 dvss 0.331238f
C4132 avss.n256 dvss 0.325944f
C4133 avss.n267 dvss 0.331238f
C4134 avss.n268 dvss 0.325944f
C4135 avss.n279 dvss 0.331238f
C4136 avss.n280 dvss 0.325944f
C4137 avss.n291 dvss 0.331238f
C4138 avss.n292 dvss 0.325944f
C4139 avss.n303 dvss 0.331238f
C4140 avss.n304 dvss 0.325944f
C4141 avss.n315 dvss 0.331238f
C4142 avss.n316 dvss 0.325944f
C4143 avss.n327 dvss 0.331238f
C4144 avss.n328 dvss 0.325944f
C4145 avss.n339 dvss 0.331238f
C4146 avss.n340 dvss 0.325944f
C4147 avss.n351 dvss 0.331238f
C4148 avss.n352 dvss 0.325944f
C4149 avss.n363 dvss 0.331238f
C4150 avss.n364 dvss 0.325944f
C4151 avss.n375 dvss 0.331238f
C4152 avss.n376 dvss 0.325944f
C4153 avss.n387 dvss 0.331238f
C4154 avss.n388 dvss 0.325944f
C4155 avss.n398 dvss 0.400393f
C4156 avss.n399 dvss 13.372f
C4157 avss.n400 dvss 6.73702f
C4158 avss.t363 dvss 9.890409f
C4159 avss.t306 dvss 9.890409f
C4160 avss.t162 dvss 9.890409f
C4161 avss.t216 dvss 9.890409f
C4162 avss.t369 dvss 9.890409f
C4163 avss.t223 dvss 9.890409f
C4164 avss.t232 dvss 9.890409f
C4165 avss.t362 dvss 10.400599f
C4166 avss.n401 dvss 5.65588f
C4167 avss.t224 dvss 5.11867f
C4168 avss.n402 dvss 5.724431f
C4169 avss.n403 dvss 0.846866f
C4170 avss.n404 dvss 0.28388f
C4171 avss.n405 dvss 0.144238f
C4172 avss.n406 dvss 0.185618f
C4173 avss.n407 dvss 1.07574f
C4174 avss.n408 dvss 1.25652f
C4175 avss.n409 dvss 1.40932f
C4176 avss.n410 dvss 0.704704f
C4177 avss.n411 dvss 0.999198f
C4178 avss.t167 dvss 0.30501f
C4179 avss.n412 dvss 3.85937f
C4180 avss.n413 dvss 60.1687f
C4181 avss.t118 dvss 0.701065f
C4182 avss.n444 dvss 0.319421f
C4183 avss.n445 dvss 0.563618f
C4184 avss.n446 dvss 0.129748f
C4185 avss.n447 dvss 0.564264f
C4186 avss.n448 dvss 0.129651f
C4187 avss.n449 dvss 0.564264f
C4188 avss.n450 dvss 0.564264f
C4189 avss.n451 dvss 2.05868f
C4190 avss.n452 dvss 0.129947f
C4191 avss.n453 dvss 0.25932f
C4192 avss.n454 dvss 0.564494f
C4193 avss.n455 dvss 2.07333f
C4194 avss.n456 dvss 2.05868f
C4195 avss.n457 dvss 2.07333f
C4196 avss.n458 dvss 0.564494f
C4197 avss.n459 dvss 0.258921f
C4198 avss.n460 dvss 0.12965f
C4199 avss.n461 dvss 0.527136f
C4200 avss.n462 dvss 0.363835f
C4201 avss.n467 dvss 0.173733f
C4202 avss.n469 dvss 0.226335f
C4203 avss.t119 dvss 1.16016f
C4204 avss.n475 dvss 0.723326f
C4205 avss.n481 dvss 0.170755f
C4206 avss.n485 dvss 1.54769f
C4207 avss.n489 dvss 0.173733f
C4208 avss.n492 dvss 0.236327f
C4209 avss.n494 dvss 0.236327f
C4210 avss.n500 dvss 0.173733f
C4211 avss.n501 dvss 0.778266f
C4212 avss.n508 dvss 0.232277f
C4213 avss.n509 dvss 0.232277f
C4214 avss.n510 dvss 0.170755f
C4215 avss.n517 dvss 0.747219f
C4216 avss.n518 dvss 0.222282f
C4217 avss.n519 dvss 1.43984f
C4218 avss.n525 dvss 0.222282f
C4219 avss.n526 dvss 1.41357f
C4220 avss.n534 dvss 0.166387f
C4221 avss.n535 dvss 0.166387f
C4222 avss.n536 dvss 0.226335f
C4223 avss.n542 dvss 1.49434f
C4224 avss.n543 dvss 0.769369f
C4225 avss.n544 dvss 0.173733f
C4226 avss.n548 dvss 0.11956f
C4227 avss.n549 dvss 0.402612f
C4228 avss.n550 dvss 42.5165f
C4229 avss.n551 dvss 47.910896f
C4230 avss.n552 dvss 7.46744f
C4231 avss.t438 dvss 1.72444f
C4232 avss.n553 dvss 1.70136f
C4233 avss.t126 dvss 1.11293f
C4234 avss.n554 dvss 0.551361f
C4235 avss.n556 dvss 0.468516f
C4236 avss.n558 dvss 0.134943f
C4237 avss.n560 dvss 0.124609f
C4238 avss.n561 dvss 0.467264f
C4239 avss.n562 dvss 1.15844f
C4240 avss.n564 dvss 0.100806f
C4241 avss.n565 dvss 0.467264f
C4242 avss.n566 dvss 0.570582f
C4243 avss.n567 dvss 0.935393f
C4244 avss.n570 dvss 0.123765f
C4245 avss.n571 dvss 0.212263f
C4246 avss.n572 dvss 0.212263f
C4247 avss.t380 dvss 2.12763f
C4248 avss.n574 dvss 0.121845f
C4249 avss.n575 dvss 0.206718f
C4250 avss.n576 dvss 2.84055f
C4251 avss.t145 dvss 1.21806f
C4252 avss.n577 dvss 9.41524f
C4253 avss.n578 dvss 46.938198f
C4254 avss.n579 dvss 1.53903f
C4255 avss.n583 dvss 0.918491f
C4256 avss.n584 dvss 1.05784f
C4257 avss.n585 dvss 0.393201f
C4258 avss.n586 dvss 0.781737f
C4259 avss.n587 dvss 0.781737f
C4260 avss.n588 dvss 0.390874f
C4261 avss.n589 dvss 1.07763f
C4262 avss.n590 dvss 0.779327f
C4263 avss.n591 dvss 0.781665f
C4264 avss.n592 dvss 1.49376f
C4265 avss.t370 dvss 1.4485f
C4266 avss.t359 dvss 1.4485f
C4267 avss.t313 dvss 1.4485f
C4268 avss.t194 dvss 1.13164f
C4269 avss.t200 dvss 1.4485f
C4270 avss.t192 dvss 1.4485f
C4271 avss.t184 dvss 1.4485f
C4272 avss.t352 dvss 4.51147f
C4273 avss.n647 dvss 2.12748f
C4274 avss.n656 dvss 2.4896f
C4275 avss.t182 dvss 1.4485f
C4276 avss.n657 dvss 1.85589f
C4277 avss.n658 dvss 2.17274f
C4278 avss.t251 dvss 0.950575f
C4279 avss.t180 dvss 0.678982f
C4280 avss.n659 dvss 1.94642f
C4281 avss.n664 dvss 0.100969f
C4282 avss.n670 dvss 1.49376f
C4283 avss.n671 dvss 2.30854f
C4284 avss.t186 dvss 1.4485f
C4285 avss.n672 dvss 2.35381f
C4286 avss.t190 dvss 1.4485f
C4287 avss.n673 dvss 1.1769f
C4288 avss.t168 dvss 1.4485f
C4289 avss.n674 dvss 1.1769f
C4290 avss.n679 dvss 0.100969f
C4291 avss.n685 dvss 0.100969f
C4292 avss.n690 dvss 1.67482f
C4293 avss.n691 dvss 1.94642f
C4294 avss.t358 dvss 0.678982f
C4295 avss.t198 dvss 0.950575f
C4296 avss.n692 dvss 1.58429f
C4297 avss.n693 dvss 2.21801f
C4298 avss.n700 dvss 0.100969f
C4299 avss.n704 dvss 0.100969f
C4300 avss.n711 dvss 2.35381f
C4301 avss.t202 dvss 1.4485f
C4302 avss.n712 dvss 0.814777f
C4303 avss.t368 dvss 1.4485f
C4304 avss.t208 dvss 1.22217f
C4305 avss.n713 dvss 1.53903f
C4306 avss.n716 dvss 1.62956f
C4307 avss.t188 dvss 1.4485f
C4308 avss.t258 dvss 0.860044f
C4309 avss.n717 dvss 1.76536f
C4310 avss.n718 dvss 1.49376f
C4311 avss.n726 dvss 0.100969f
C4312 avss.n731 dvss 2.03695f
C4313 avss.n732 dvss 1.76536f
C4314 avss.t196 dvss 1.4485f
C4315 avss.n733 dvss 0.452653f
C4316 avss.t178 dvss 1.4485f
C4317 avss.n734 dvss 2.35381f
C4318 avss.n740 dvss 0.100969f
C4319 avss.n745 dvss 1.90115f
C4320 avss.t204 dvss 1.4485f
C4321 avss.n746 dvss 2.21801f
C4322 avss.n747 dvss 1.4485f
C4323 avss.t206 dvss 1.4485f
C4324 avss.n748 dvss 1.58429f
C4325 avss.n759 dvss 2.65558f
C4326 avss.t143 dvss 1.4485f
C4327 avss.n760 dvss 1.55412f
C4328 avss.n761 dvss 0.694069f
C4329 avss.t141 dvss 1.4485f
C4330 avss.n762 dvss 2.24819f
C4331 avss.n775 dvss 1.65973f
C4332 avss.t139 dvss 1.4485f
C4333 avss.n776 dvss 2.35381f
C4334 avss.t137 dvss 1.4485f
C4335 avss.t233 dvss 1.4485f
C4336 avss.n777 dvss 1.68991f
C4337 avss.n788 dvss 2.79138f
C4338 avss.t230 dvss 1.35796f
C4339 avss.n789 dvss 0.105618f
C4340 avss.n790 dvss 0.781737f
C4341 avss.n791 dvss 0.781665f
C4342 avss.n792 dvss 0.781665f
C4343 avss.n793 dvss 0.663999f
C4344 avss.n794 dvss 0.568078f
C4345 avss.n796 dvss 0.202626f
C4346 avss.n800 dvss 0.203153f
C4347 avss.n802 dvss 0.11116f
C4348 avss.n804 dvss 0.113222f
C4349 avss.n805 dvss 0.108871f
C4350 avss.n806 dvss 0.12866f
C4351 avss.n807 dvss 0.512839f
C4352 avss.n808 dvss 0.998447f
C4353 avss.t14 dvss 0.656996f
C4354 avss.t20 dvss 0.376292f
C4355 avss.t10 dvss 0.376292f
C4356 avss.t12 dvss 0.376292f
C4357 avss.t18 dvss 0.282216f
C4358 avss.n809 dvss 0.191392f
C4359 avss.n810 dvss 0.103916f
C4360 avss.n812 dvss 0.214925f
C4361 avss.n813 dvss 0.109922f
C4362 avss.t68 dvss 7.03696f
C4363 avss.n814 dvss 0.943753f
C4364 avss.n815 dvss 0.295739f
C4365 avss.n816 dvss 0.262183f
C4366 avss.n817 dvss 0.124609f
C4367 avss.t132 dvss 1.11293f
C4368 avss.n818 dvss 0.262183f
C4369 avss.t67 dvss 1.11293f
C4370 avss.n821 dvss 0.551361f
C4371 avss.t419 dvss 1.72444f
C4372 avss.n823 dvss 0.791962f
C4373 avss.t437 dvss 1.72444f
C4374 avss.n824 dvss 0.791962f
C4375 avss.t416 dvss 1.72444f
C4376 avss.n825 dvss 0.791962f
C4377 avss.t424 dvss 1.72444f
C4378 avss.n826 dvss 0.791962f
C4379 avss.t415 dvss 1.72444f
C4380 avss.n827 dvss 0.791962f
C4381 avss.t433 dvss 1.72444f
C4382 avss.n828 dvss 0.791962f
C4383 avss.t414 dvss 1.72444f
C4384 avss.n829 dvss 0.875609f
C4385 avss.n830 dvss 0.215816f
C4386 avss.n832 dvss 0.551361f
C4387 avss.n834 dvss 0.134943f
C4388 avss.n835 dvss 0.468516f
C4389 avss.n837 dvss 0.13562f
C4390 avss.n838 dvss 0.623434f
C4391 avss.n839 dvss 0.536805f
C4392 avss.t292 dvss 8.90292f
C4393 avss.t294 dvss 6.67719f
C4394 avss.t64 dvss 7.03696f
C4395 avss.t288 dvss 8.90292f
C4396 avss.t290 dvss 6.67719f
C4397 avss.n840 dvss 4.45146f
C4398 avss.n841 dvss 0.935393f
C4399 avss.n842 dvss 0.943753f
C4400 avss.n843 dvss 2.96211f
C4401 avss.n844 dvss 0.243423f
C4402 avss.t147 dvss 0.286129f
C4403 avss.t22 dvss 0.376292f
C4404 avss.t16 dvss 0.376292f
C4405 avss.t24 dvss 0.282216f
C4406 avss.n846 dvss 0.214925f
C4407 avss.n848 dvss 0.103916f
C4408 avss.n849 dvss 0.123762f
C4409 avss.n850 dvss 1.53958f
C4410 avss.n856 dvss 2.7612f
C4411 avss.t158 dvss 7.01616f
C4412 avss.t408 dvss 11.4069f
C4413 avss.t235 dvss 11.4069f
C4414 avss.t356 dvss 11.4069f
C4415 avss.t365 dvss 11.4069f
C4416 avss.t159 dvss 7.77059f
C4417 avss.t354 dvss 9.535951f
C4418 avss.t164 dvss 11.4069f
C4419 avss.t321 dvss 11.4069f
C4420 avss.t375 dvss 9.33979f
C4421 avss.n857 dvss 34.361603f
C4422 avss.t387 dvss 2.02766f
C4423 avss.n858 dvss 32.593002f
C4424 avss.n859 dvss 19.463f
C4425 avss.n860 dvss 15.231599f
C4426 avss.t55 dvss 23.4704f
C4427 avss.n861 dvss 0.651819f
C4428 avss.n862 dvss 0.651819f
C4429 avss.n863 dvss 0.202832f
C4430 avss.n864 dvss 0.202832f
C4431 avss.n865 dvss 0.680655f
C4432 avss.n866 dvss 0.350575f
C4433 avss.t56 dvss 0.153822f
C4434 avss.t54 dvss 1.80863f
C4435 avss.n867 dvss 1.60166f
C4436 avss.n868 dvss 0.703137f
C4437 avss.t110 dvss 2.31618f
C4438 avss.n869 dvss 1.84774f
C4439 avss.t75 dvss 0.153822f
C4440 avss.t74 dvss 1.80863f
C4441 avss.n870 dvss 1.60166f
C4442 avss.n871 dvss 0.705082f
C4443 avss.n872 dvss 0.492614f
C4444 avss.n873 dvss 0.196259f
C4445 avss.n874 dvss 0.196259f
C4446 avss.t152 dvss 4.88034f
C4447 avss.t151 dvss 5.99104f
C4448 avss.t153 dvss 5.99104f
C4449 avss.n875 dvss 0.398376f
C4450 avss.t150 dvss 50.6632f
C4451 avss.n877 dvss 0.392413f
C4452 avss.n878 dvss 0.403922f
C4453 avss.n879 dvss 0.796389f
C4454 avss.n880 dvss 0.702854f
C4455 avss.t314 dvss 0.232713f
C4456 avss.n881 dvss 1.07289f
C4457 avss.n882 dvss 0.710956f
C4458 avss.n883 dvss 0.700632f
C4459 avss.n884 dvss 0.586865f
C4460 avss.n885 dvss 0.781737f
C4461 avss.n886 dvss 22.0818f
C4462 avss.n887 dvss 16.7307f
C4463 avss.n888 dvss 0.645429f
C4464 avss.n889 dvss 0.379139f
C4465 avss.n890 dvss 0.660264f
C4466 avss.n891 dvss 0.680655f
C4467 avss.n892 dvss 0.625282f
C4468 avss.n893 dvss 0.366014f
C4469 avss.n894 dvss 0.645429f
C4470 avss.n895 dvss 23.692099f
C4471 avss.n896 dvss 30.689901f
C4472 avss.n897 dvss 15.702001f
C4473 avss.t256 dvss 0.793567f
C4474 avss.n898 dvss 1.3673f
C4475 avss.t252 dvss 2.15263f
C4476 avss.t254 dvss 1.2091f
C4477 avss.n899 dvss 1.11224f
C4478 avss.n900 dvss 0.206718f
C4479 avss.n903 dvss 0.295739f
C4480 avss.n904 dvss 0.536805f
C4481 avss.n905 dvss 0.61967f
C4482 avss.n907 dvss 2.15301f
C4483 avss.n908 dvss 0.208832f
C4484 avss.n909 dvss 0.100213f
C4485 avss.n910 dvss 0.111185f
C4486 avss.n911 dvss 0.309868f
C4487 avss.n912 dvss 1.23943f
C4488 avss.t63 dvss 1.11293f
C4489 avss.n913 dvss 0.551361f
C4490 avss.n916 dvss 0.262183f
C4491 avss.n917 dvss 0.262183f
C4492 avss.n918 dvss 0.218554f
C4493 avss.t418 dvss 1.71234f
C4494 avss.n919 dvss 0.867243f
C4495 avss.t436 dvss 1.71234f
C4496 avss.n920 dvss 0.777737f
C4497 avss.t421 dvss 1.71234f
C4498 avss.n921 dvss 0.777737f
C4499 avss.t425 dvss 1.71234f
C4500 avss.n922 dvss 0.777737f
C4501 avss.t422 dvss 1.71234f
C4502 avss.n923 dvss 0.777737f
C4503 avss.t439 dvss 1.71234f
C4504 avss.n924 dvss 0.777737f
C4505 avss.t423 dvss 1.71234f
C4506 avss.n925 dvss 0.777737f
C4507 avss.t440 dvss 1.71234f
C4508 avss.n926 dvss 0.830167f
C4509 avss.n927 dvss 3.93027f
C4510 avss.n928 dvss 10.9261f
C4511 avss.n929 dvss 12.2517f
C4512 avss.t429 dvss 0.138473f
C4513 avss.t432 dvss 0.138236f
C4514 avss.n930 dvss 0.13774f
C4515 avss.t431 dvss 0.138236f
C4516 avss.t103 dvss 0.135063f
C4517 avss.t41 dvss 0.135812f
C4518 avss.n932 dvss 0.284594f
C4519 avss.n933 dvss 0.134109f
C4520 avss.n934 dvss 4.41396f
C4521 avss.n935 dvss 4.74252f
C4522 avss.n936 dvss 0.208832f
C4523 avss.n937 dvss 0.100213f
C4524 avss.n938 dvss 0.111185f
C4525 avss.n939 dvss 0.37638f
C4526 avss.n940 dvss 1.23943f
C4527 avss.t99 dvss 1.11293f
C4528 avss.n941 dvss 0.551361f
C4529 avss.n944 dvss 0.262183f
C4530 avss.n945 dvss 0.262183f
C4531 avss.n946 dvss 0.218554f
C4532 avss.t430 dvss 1.71234f
C4533 avss.n947 dvss 0.867243f
C4534 avss.t413 dvss 1.71234f
C4535 avss.n948 dvss 0.777737f
C4536 avss.t443 dvss 1.71234f
C4537 avss.n949 dvss 0.777737f
C4538 avss.t434 dvss 1.71234f
C4539 avss.n950 dvss 0.777737f
C4540 avss.t417 dvss 1.71234f
C4541 avss.n951 dvss 0.777737f
C4542 avss.t435 dvss 1.71234f
C4543 avss.n952 dvss 0.777737f
C4544 avss.t420 dvss 1.71234f
C4545 avss.n953 dvss 0.777737f
C4546 avss.t444 dvss 1.71234f
C4547 avss.n954 dvss 0.830167f
C4548 avss.n955 dvss 3.94664f
C4549 avss.t442 dvss 1.72444f
C4550 avss.n956 dvss 1.70136f
C4551 avss.t412 dvss 1.72444f
C4552 avss.n957 dvss 0.791962f
C4553 avss.t428 dvss 1.72444f
C4554 avss.n958 dvss 0.791962f
C4555 avss.t411 dvss 1.72444f
C4556 avss.n959 dvss 0.791962f
C4557 avss.t427 dvss 1.72444f
C4558 avss.n960 dvss 0.791962f
C4559 avss.t441 dvss 1.72444f
C4560 avss.n961 dvss 0.791962f
C4561 avss.t410 dvss 1.72444f
C4562 avss.n962 dvss 0.791962f
C4563 avss.t426 dvss 1.72444f
C4564 avss.n963 dvss 0.875609f
C4565 avss.n964 dvss 0.215816f
C4566 avss.n966 dvss 0.551361f
C4567 avss.n968 dvss 0.134943f
C4568 avss.t111 dvss 1.11293f
C4569 avss.n969 dvss 0.551361f
C4570 avss.n971 dvss 0.124609f
C4571 avss.n972 dvss 0.467264f
C4572 avss.n973 dvss 0.262183f
C4573 avss.n975 dvss 1.15844f
C4574 avss.n976 dvss 0.191392f
C4575 avss.n977 dvss 0.103916f
C4576 avss.n978 dvss 0.214925f
C4577 avss.n980 dvss 0.12866f
C4578 avss.n982 dvss 0.214925f
C4579 avss.t45 dvss 2.54844f
C4580 avss.n984 dvss 0.604058f
C4581 avss.t296 dvss 3.72391f
C4582 avss.n985 dvss 3.10701f
C4583 avss.t274 dvss 2.69334f
C4584 avss.t100 dvss 3.10701f
C4585 avss.t282 dvss 4.22348f
C4586 avss.t270 dvss 4.27164f
C4587 avss.n987 dvss 1.5535f
C4588 avss.n988 dvss 0.935393f
C4589 avss.n989 dvss 0.536805f
C4590 avss.n991 dvss 0.295739f
C4591 avss.n993 dvss 0.295739f
C4592 avss.n994 dvss 0.536805f
C4593 avss.n995 dvss 0.935393f
C4594 avss.n996 dvss 3.89249f
C4595 avss.n997 dvss 0.212263f
C4596 avss.n999 dvss 0.121845f
C4597 avss.n1000 dvss 0.123765f
C4598 avss.n1001 dvss 0.212263f
C4599 avss.n1002 dvss 4.32707f
C4600 avss.n1003 dvss 34.63f
C4601 avss.n1004 dvss 38.7109f
C4602 avss.n1005 dvss 0.781737f
C4603 avss.n1006 dvss 0.580675f
C4604 avss.n1007 dvss 0.674107f
C4605 avss.n1008 dvss 0.77145f
C4606 avss.n1009 dvss 0.729086f
C4607 avss.n1010 dvss 7.69067f
C4608 avss.n1011 dvss 4.77871f
C4609 avss.n1012 dvss 0.13157f
C4610 avss.n1013 dvss 1.50175f
C4611 avss.n1014 dvss 1.5191f
C4612 avss.n1015 dvss 2.83673f
C4613 avss.n1016 dvss 2.83033f
C4614 avss.n1017 dvss 1.71896f
C4615 avss.n1018 dvss 1.72077f
C4616 avss.n1019 dvss 1.72077f
C4617 avss.n1020 dvss 1.65742f
C4618 avss.t398 dvss -1.12358f
C4619 avss.t71 dvss 5.09784f
C4620 avss.t176 dvss 4.47002f
C4621 avss.t343 dvss 6.65481f
C4622 avss.t98 dvss 7.30774f
C4623 avss.t247 dvss 4.47002f
C4624 avss.t340 dvss 6.10234f
C4625 avss.t384 dvss 4.59559f
C4626 avss.n1021 dvss 0.642362f
C4627 avss.n1022 dvss 1.08754f
C4628 avss.n1023 dvss 3.39019f
C4629 avss.n1024 dvss 1.08754f
C4630 avss.n1025 dvss 0.640638f
C4631 avss.n1026 dvss 0.742396f
C4632 avss.n1027 dvss 0.162702f
C4633 avss.n1028 dvss 1.25073f
C4634 avss.n1029 dvss 1.25073f
C4635 avss.t76 dvss 4.08169f
C4636 avss.n1030 dvss 0.162702f
C4637 avss.t77 dvss 0.200808f
C4638 avss.n1031 dvss 1.54091f
C4639 avss.n1032 dvss 0.457138f
C4640 avss.n1033 dvss 0.197783f
C4641 avss.n1034 dvss 0.501164f
C4642 avss.n1035 dvss 0.457138f
C4643 avss.t88 dvss 4.08169f
C4644 avss.n1036 dvss 1.54091f
C4645 avss.t89 dvss 0.200808f
C4646 avss.n1037 dvss 0.162702f
C4647 avss.n1038 dvss 1.25073f
C4648 avss.n1039 dvss 0.162702f
C4649 avss.n1040 dvss 1.25073f
C4650 avss.t129 dvss 4.08169f
C4651 avss.t131 dvss 0.15847f
C4652 avss.n1041 dvss 1.54091f
C4653 avss.n1042 dvss 0.399913f
C4654 avss.n1043 dvss 0.270268f
C4655 avss.n1044 dvss 0.500734f
C4656 avss.n1045 dvss 0.197352f
C4657 avss.n1046 dvss 0.270268f
C4658 avss.n1047 dvss 1.02499f
C4659 avss.n1048 dvss 1.02499f
C4660 avss.n1049 dvss 0.270268f
C4661 avss.t90 dvss 4.08169f
C4662 avss.t92 dvss 0.15847f
C4663 avss.n1050 dvss 1.54091f
C4664 avss.n1051 dvss 0.399913f
C4665 avss.n1052 dvss 0.162702f
C4666 avss.n1053 dvss 1.25073f
C4667 avss.n1054 dvss 1.25073f
C4668 avss.t52 dvss 4.08169f
C4669 avss.n1055 dvss 0.162702f
C4670 avss.t53 dvss 0.200808f
C4671 avss.n1056 dvss 1.54091f
C4672 avss.n1057 dvss 0.457138f
C4673 avss.n1058 dvss 0.150973f
C4674 avss.n1059 dvss 0.222383f
C4675 avss.n1060 dvss 0.457138f
C4676 avss.t36 dvss 4.08169f
C4677 avss.n1061 dvss 1.54091f
C4678 avss.t38 dvss 0.200808f
C4679 avss.n1062 dvss 0.162702f
C4680 avss.n1063 dvss 1.25073f
C4681 avss.n1064 dvss 0.162702f
C4682 avss.n1065 dvss 1.25073f
C4683 avss.t80 dvss 4.08169f
C4684 avss.t83 dvss 0.15847f
C4685 avss.n1066 dvss 1.54091f
C4686 avss.n1067 dvss 0.399913f
C4687 avss.n1068 dvss 0.270268f
C4688 avss.n1069 dvss 0.221953f
C4689 avss.n1070 dvss 0.44987f
C4690 avss.n1071 dvss 0.270268f
C4691 avss.n1072 dvss 1.04439f
C4692 avss.n1073 dvss 1.08301f
C4693 avss.n1074 dvss 0.856759f
C4694 avss.n1075 dvss 0.149546f
C4695 avss.n1076 dvss 0.202714f
C4696 avss.n1077 dvss 0.149546f
C4697 avss.n1078 dvss 0.12851f
C4698 avss.n1079 dvss 0.398376f
C4699 avss.n1080 dvss 6.40369f
C4700 avss.n1081 dvss 7.28262f
C4701 avss.n1082 dvss 0.296289f
C4702 avss.n1084 dvss 0.119748f
C4703 avss.n1085 dvss 0.109607f
C4704 avss.t336 dvss 0.212474f
C4705 avss.n1086 dvss 0.417142f
C4706 avss.n1087 dvss 0.155688f
C4707 avss.n1088 dvss 0.558435f
C4708 avss.t342 dvss 0.212474f
C4709 avss.n1089 dvss 0.417358f
C4710 avss.n1090 dvss 0.15455f
C4711 avss.n1091 dvss 0.119748f
C4712 avss.n1093 dvss 0.296289f
C4713 avss.n1094 dvss 2.23501f
C4714 avss.t37 dvss 6.05211f
C4715 avss.n1095 dvss 7.25751f
C4716 avss.n1096 dvss 0.205002f
C4717 avss.n1097 dvss 0.113055f
C4718 avss.n1098 dvss 0.298414f
C4719 avss.n1099 dvss 0.113551f
C4720 avss.n1100 dvss 0.205002f
C4721 avss.n1101 dvss 9.492519f
C4722 avss.t174 dvss 13.0585f
C4723 avss.t157 dvss 10.697901f
C4724 avss.n1102 dvss 20.218f
C4725 avss.t243 dvss 17.4983f
C4726 avss.t304 dvss 15.382699f
C4727 avss.t161 dvss 15.5227f
C4728 avss.t215 dvss 15.5227f
C4729 avss.t136 dvss 15.5227f
C4730 avss.t322 dvss 15.5227f
C4731 avss.t175 dvss 12.4633f
C4732 avss.n1103 dvss 17.4412f
C4733 avss.n1104 dvss 12.1641f
C4734 avss.t28 dvss 2.74842f
C4735 avss.n1110 dvss 0.156863f
C4736 avss.n1111 dvss 0.329806f
C4737 avss.n1112 dvss 0.617375f
C4738 por_dig_0.net22.n17 dvss 0.290913f
C4739 por_dig_0.net22.n18 dvss 0.220093f
C4740 por_dig_0.net22.n21 dvss 0.245438f
C4741 por_dig_0.net22.n26 dvss 0.125219f
C4742 por_dig_0.net22.n27 dvss 0.244466f
C4743 por_dig_0.clknet_1_1__leaf_osc_ck.n17 dvss 0.130985f
C4744 por_dig_0.clknet_1_1__leaf_osc_ck.n20 dvss 0.122095f
C4745 por_dig_0.clknet_1_1__leaf_osc_ck.n27 dvss 0.267282f
C4746 por_dig_0.clknet_1_1__leaf_osc_ck.n28 dvss 0.267987f
C4747 por_dig_0.clknet_1_1__leaf_osc_ck.n32 dvss 0.304204f
C4748 por_dig_0.clknet_1_1__leaf_osc_ck.n35 dvss 0.186102f
C4749 por_dig_0.clknet_1_1__leaf_osc_ck.n36 dvss 0.131031f
C4750 por_dig_0.clknet_1_1__leaf_osc_ck.n48 dvss 0.119959f
C4751 vbg_1v2.n0 dvss 0.46714f
C4752 vbg_1v2.n1 dvss 4.23283f
C4753 vbg_1v2.t16 dvss 1.96783f
C4754 vbg_1v2.t37 dvss 1.8832f
C4755 vbg_1v2.n2 dvss 1.56821f
C4756 vbg_1v2.t15 dvss 1.8832f
C4757 vbg_1v2.n3 dvss 0.828262f
C4758 vbg_1v2.t36 dvss 1.8832f
C4759 vbg_1v2.n4 dvss 0.828262f
C4760 vbg_1v2.t3 dvss 1.8832f
C4761 vbg_1v2.n5 dvss 0.828262f
C4762 vbg_1v2.t35 dvss 1.8832f
C4763 vbg_1v2.n6 dvss 0.828262f
C4764 vbg_1v2.t12 dvss 1.8832f
C4765 vbg_1v2.n7 dvss 0.828262f
C4766 vbg_1v2.t34 dvss 1.8832f
C4767 vbg_1v2.n8 dvss 0.979621f
C4768 vbg_1v2.t25 dvss 1.98466f
C4769 vbg_1v2.t43 dvss 1.89884f
C4770 vbg_1v2.n9 dvss 1.60346f
C4771 vbg_1v2.t24 dvss 1.89884f
C4772 vbg_1v2.n10 dvss 0.846485f
C4773 vbg_1v2.t42 dvss 1.89884f
C4774 vbg_1v2.n11 dvss 0.846485f
C4775 vbg_1v2.t10 dvss 1.89884f
C4776 vbg_1v2.n12 dvss 0.846485f
C4777 vbg_1v2.t41 dvss 1.89884f
C4778 vbg_1v2.n13 dvss 0.846485f
C4779 vbg_1v2.t21 dvss 1.89884f
C4780 vbg_1v2.n14 dvss 0.846485f
C4781 vbg_1v2.t40 dvss 1.89884f
C4782 vbg_1v2.n15 dvss 0.936128f
C4783 vbg_1v2.n16 dvss 0.767501f
C4784 vbg_1v2.n17 dvss 1.63958f
C4785 vbg_1v2.n18 dvss 1.09863f
C4786 vbg_1v2.t27 dvss 1.7581f
C4787 vbg_1v2.t19 dvss 1.60872f
C4788 vbg_1v2.n19 dvss 1.09417f
C4789 vbg_1v2.t39 dvss 1.7581f
C4790 vbg_1v2.n22 dvss 1.09417f
C4791 vbg_1v2.t31 dvss 1.60872f
C4792 vbg_1v2.n23 dvss 1.09417f
C4793 vbg_1v2.t14 dvss 1.7581f
C4794 vbg_1v2.n26 dvss 1.09417f
C4795 vbg_1v2.t7 dvss 1.60872f
C4796 vbg_1v2.n27 dvss 1.09417f
C4797 vbg_1v2.t38 dvss 1.7581f
C4798 vbg_1v2.n30 dvss 1.09417f
C4799 vbg_1v2.t30 dvss 1.60872f
C4800 vbg_1v2.n31 dvss 1.09417f
C4801 vbg_1v2.t13 dvss 1.7581f
C4802 vbg_1v2.n34 dvss 1.09417f
C4803 vbg_1v2.t6 dvss 1.60872f
C4804 vbg_1v2.n35 dvss 1.09417f
C4805 vbg_1v2.t26 dvss 1.7581f
C4806 vbg_1v2.n38 dvss 1.09417f
C4807 vbg_1v2.t17 dvss 1.60872f
C4808 vbg_1v2.n39 dvss 1.09417f
C4809 vbg_1v2.t33 dvss 1.7581f
C4810 vbg_1v2.n42 dvss 1.09417f
C4811 vbg_1v2.t29 dvss 1.60872f
C4812 vbg_1v2.n43 dvss 1.09417f
C4813 vbg_1v2.t11 dvss 1.7581f
C4814 vbg_1v2.n46 dvss 1.09417f
C4815 vbg_1v2.t4 dvss 1.60872f
C4816 vbg_1v2.n47 dvss 1.09417f
C4817 vbg_1v2.n48 dvss 1.37481f
C4818 vbg_1v2.n49 dvss 1.73642f
C4819 vbg_1v2.n50 dvss 0.108637f
C4820 vbg_1v2.n51 dvss 0.109088f
C4821 vbg_1v2.n52 dvss 0.109088f
C4822 vbg_1v2.n53 dvss 0.109088f
C4823 vbg_1v2.t20 dvss 0.316935f
C4824 vbg_1v2.n54 dvss 0.213144f
C4825 vbg_1v2.t23 dvss 0.316673f
C4826 vbg_1v2.n55 dvss 0.213144f
C4827 vbg_1v2.t18 dvss 0.316673f
C4828 vbg_1v2.n56 dvss 0.109088f
C4829 vbg_1v2.n57 dvss 0.109088f
C4830 vbg_1v2.t22 dvss 0.316673f
C4831 vbg_1v2.n58 dvss 0.109088f
C4832 vbg_1v2.t32 dvss 0.316673f
C4833 vbg_1v2.n59 dvss 0.109088f
C4834 vbg_1v2.n60 dvss 0.109088f
C4835 vbg_1v2.t5 dvss 0.316673f
C4836 vbg_1v2.n61 dvss 0.109088f
C4837 vbg_1v2.t9 dvss 0.316673f
C4838 vbg_1v2.n62 dvss 0.109088f
C4839 vbg_1v2.n63 dvss 0.109088f
C4840 vbg_1v2.t2 dvss 0.316673f
C4841 vbg_1v2.n64 dvss 0.109088f
C4842 vbg_1v2.t8 dvss 0.316673f
C4843 vbg_1v2.n65 dvss 0.108637f
C4844 vbg_1v2.n66 dvss 0.101228f
C4845 vbg_1v2.t28 dvss 0.316673f
C4846 vbg_1v2.n67 dvss 0.101228f
C4847 porb.n30 dvss 0.712335f
C4848 por_ana_0.comparator_1.n1.n0 dvss 0.795794f
C4849 por_ana_0.comparator_1.n1.n1 dvss 0.765455f
C4850 por_ana_0.comparator_1.n1.t16 dvss 0.177538f
C4851 por_ana_0.comparator_1.n1.t11 dvss 0.177346f
C4852 por_ana_0.comparator_1.n1.t5 dvss 0.177346f
C4853 por_ana_0.comparator_1.n1.t19 dvss 0.177346f
C4854 por_ana_0.comparator_1.n1.t12 dvss 0.177346f
C4855 por_ana_0.comparator_1.n1.t6 dvss 0.177346f
C4856 por_ana_0.comparator_1.n1.t18 dvss 0.177346f
C4857 por_ana_0.comparator_1.n1.t8 dvss 0.177346f
C4858 por_ana_0.comparator_1.n1.t14 dvss 0.172786f
C4859 por_ana_0.comparator_1.n1.t9 dvss 0.172595f
C4860 por_ana_0.comparator_1.n1.t17 dvss 0.172595f
C4861 por_ana_0.comparator_1.n1.t15 dvss 0.172595f
C4862 por_ana_0.comparator_1.n1.t10 dvss 0.172595f
C4863 por_ana_0.comparator_1.n1.t4 dvss 0.172595f
C4864 por_ana_0.comparator_1.n1.t13 dvss 0.172595f
C4865 por_ana_0.comparator_1.n1.t7 dvss 0.172595f
C4866 por_ana_0.comparator_1.n1.n3 dvss 0.590043f
C4867 por_ana_0.comparator_1.n1.n4 dvss 0.590765f
C4868 por_ana_0.comparator_1.n0.n0 dvss 1.12136f
C4869 por_ana_0.comparator_1.n0.t7 dvss 0.165842f
C4870 por_ana_0.comparator_1.n0.t5 dvss 0.165666f
C4871 por_ana_0.comparator_1.n0.n2 dvss 0.348475f
C4872 por_ana_0.comparator_1.n0.t8 dvss 0.161403f
C4873 por_ana_0.comparator_1.n0.t6 dvss 0.161228f
C4874 por_ana_0.comparator_1.n0.t2 dvss 0.151863f
C4875 dvdd.n0 dvss 4.315f
C4876 dvdd.n1 dvss 0.128259f
C4877 dvdd.n2 dvss 5.28458f
C4878 dvdd.t1802 dvss 0.124773f
C4879 dvdd.t1768 dvss 0.124547f
C4880 dvdd.t1745 dvss 0.124547f
C4881 dvdd.t1673 dvss 0.124773f
C4882 dvdd.t1564 dvss 0.124547f
C4883 dvdd.n328 dvss 0.686693f
C4884 dvdd.t1537 dvss 0.220006f
C4885 dvdd.t1780 dvss 0.104035f
C4886 dvdd.t1649 dvss 0.11597f
C4887 dvdd.t1593 dvss 0.219608f
C4888 dvdd.n611 dvss 0.244721f
C4889 dvdd.t1707 dvss 0.219608f
C4890 dvdd.n912 dvss 0.244721f
C4891 dvdd.n1201 dvss 0.244721f
C4892 dvdd.n1485 dvss 0.244721f
C4893 dvdd.n1786 dvss 0.244721f
C4894 dvdd.n2088 dvss 0.244721f
C4895 dvdd.t70 dvss 0.925901f
C4896 dvdd.t325 dvss 0.368746f
C4897 dvdd.n2147 dvss 0.337134f
C4898 dvdd.t668 dvss 0.12511f
C4899 dvdd.t737 dvss 0.167911f
C4900 dvdd.n2228 dvss 0.646984f
C4901 dvdd.n2358 dvss 0.244721f
C4902 dvdd.n2646 dvss 0.188939f
C4903 dvdd.n2647 dvss 5.04938f
C4904 dvdd.n2757 dvss 0.131822f
C4905 dvdd.n2758 dvss 0.468361f
C4906 dvdd.n2759 dvss 0.425937f
C4907 dvdd.n2802 dvss 0.434762f
C4908 dvdd.n2872 dvss 0.401794f
C4909 dvdd.n2929 dvss 0.338711f
C4910 dvdd.n2930 dvss 0.121734f
C4911 dvdd.n2931 dvss 0.264415f
C4912 dvdd.n2932 dvss 0.264362f
C4913 dvdd.n2933 dvss 0.990506f
C4914 dvdd.n2934 dvss 0.265145f
C4915 dvdd.n2935 dvss 1.00069f
C4916 dvdd.n2936 dvss 0.990298f
C4917 dvdd.n2937 dvss 1.00048f
C4918 dvdd.n2938 dvss 0.265092f
C4919 dvdd.n2939 dvss 0.12171f
C4920 dvdd.n2940 dvss 0.629012f
C4921 dvdd.n2941 dvss 0.174606f
C4922 dvdd.n2942 dvss 0.187177f
C4923 dvdd.n2969 dvss 0.100133f
C4924 dvdd.n3083 dvss 0.128231f
C4925 dvdd.n3094 dvss 0.559299f
C4926 dvdd.n3095 dvss 11.918799f
C4927 dvdd.n3096 dvss 6.38099f
C4928 dvdd.n3099 dvss 0.105395f
C4929 dvdd.n3100 dvss 0.742085f
C4930 dvdd.n3101 dvss 6.46094f
C4931 dvdd.n3102 dvss 0.890873f
C4932 dvdd.n3103 dvss 0.391202f
C4933 dvdd.n3104 dvss 0.849403f
C4934 dvdd.n3105 dvss 0.390614f
C4935 dvdd.n3106 dvss 0.849403f
C4936 dvdd.n3107 dvss 3.23911f
C4937 dvdd.n3108 dvss 0.852197f
C4938 dvdd.n3109 dvss 3.28186f
C4939 dvdd.n3110 dvss 3.23911f
C4940 dvdd.n3111 dvss 3.28186f
C4941 dvdd.n3112 dvss 0.852197f
C4942 dvdd.n3113 dvss 0.391202f
C4943 dvdd.n3114 dvss 0.390614f
C4944 dvdd.n3115 dvss 0.956515f
C4945 dvdd.n3116 dvss 0.860861f
C4946 dvdd.n3136 dvss 0.101374f
C4947 dvdd.n3142 dvss 0.184049f
C4948 dvdd.t1358 dvss 0.163124f
C4949 dvdd.t1356 dvss 0.121831f
C4950 dvdd.t1354 dvss 0.121831f
C4951 dvdd.t445 dvss 0.121831f
C4952 dvdd.t443 dvss 0.121831f
C4953 dvdd.t447 dvss 0.121831f
C4954 dvdd.t1288 dvss 0.141107f
C4955 dvdd.t1360 dvss 0.179661f
C4956 dvdd.t1362 dvss 0.198938f
C4957 dvdd.t1352 dvss 0.102168f
C4958 dvdd.t242 dvss 0.138408f
C4959 dvdd.t236 dvss 0.121831f
C4960 dvdd.t234 dvss 0.121831f
C4961 dvdd.t240 dvss 0.121831f
C4962 dvdd.t244 dvss 0.121831f
C4963 dvdd.t238 dvss 0.109878f
C4964 dvdd.t1283 dvss 0.113734f
C4965 dvdd.t1421 dvss 0.117204f
C4966 dvdd.t1423 dvss 0.115933f
C4967 dvdd.n3144 dvss 0.161458f
C4968 dvdd.n3154 dvss 1.22583f
C4969 dvdd.n3155 dvss 1.14836f
C4970 por_ana_0.ibias_gen_0.Mt4 dvss 1.11393f
C4971 por_ana_0.ibias_gen_0.vn0.n0 dvss 1.0805f
C4972 por_ana_0.ibias_gen_0.vn0.n1 dvss 1.39652f
C4973 por_ana_0.ibias_gen_0.vn0.n2 dvss 0.142325f
C4974 por_ana_0.ibias_gen_0.vn0.n3 dvss 0.874872f
C4975 por_ana_0.ibias_gen_0.vn0.t19 dvss 2.24075f
C4976 por_ana_0.ibias_gen_0.vn0.t2 dvss 2.19836f
C4977 por_ana_0.ibias_gen_0.vn0.n4 dvss 0.920525f
C4978 por_ana_0.ibias_gen_0.vn0.n5 dvss 0.111014f
C4979 por_ana_0.ibias_gen_0.vn0.n6 dvss 0.198283f
C4980 por_ana_0.ibias_gen_0.vn0.n7 dvss 0.161371f
C4981 por_ana_0.ibias_gen_0.vn0.t4 dvss 2.16084f
C4982 por_ana_0.ibias_gen_0.vn0.n8 dvss 1.01955f
C4983 por_ana_0.ibias_gen_0.vn0.n9 dvss 1.87632f
C4984 por_ana_0.ibias_gen_0.vn0.t20 dvss 2.16084f
C4985 por_ana_0.ibias_gen_0.vn0.n10 dvss 1.71213f
C4986 por_ana_0.ibias_gen_0.vn0.n11 dvss 0.975041f
C4987 por_ana_0.ibias_gen_0.vn0.t14 dvss 0.202556f
C4988 por_ana_0.ibias_gen_0.vn0.n12 dvss 0.12274f
C4989 por_ana_0.ibias_gen_0.vn0.n13 dvss 0.12274f
C4990 por_ana_0.ibias_gen_0.vn0.n14 dvss 0.12274f
C4991 por_ana_0.ibias_gen_0.vn0.n15 dvss 0.12274f
C4992 por_ana_0.ibias_gen_0.vn0.n16 dvss 0.12274f
C4993 por_ana_0.ibias_gen_0.vp0.n0 dvss 0.777153f
C4994 por_ana_0.ibias_gen_0.vp0.n1 dvss 0.217103f
C4995 por_ana_0.ibias_gen_0.vp0.n3 dvss 0.886385f
C4996 por_ana_0.ibias_gen_0.vp0.n5 dvss 0.157271f
C4997 por_ana_0.ibias_gen_0.vp0.t3 dvss 1.72871f
C4998 por_ana_0.ibias_gen_0.vp0.n6 dvss 1.47471f
C4999 por_ana_0.ibias_gen_0.vp0.n7 dvss 0.724776f
C5000 por_ana_0.ibias_gen_0.vp0.t12 dvss 1.76142f
C5001 por_ana_0.ibias_gen_0.vp0.t13 dvss 1.69947f
C5002 por_ana_0.ibias_gen_0.vp0.n8 dvss 1.47471f
C5003 por_ana_0.ibias_gen_0.vp0.n9 dvss 0.800719f
C5004 por_ana_0.ibias_gen_0.vp0.t1 dvss 1.69947f
C5005 por_ana_0.ibias_gen_0.vp0.n10 dvss 0.798648f
C5006 por_ana_0.ibias_gen_0.vp0.n11 dvss 0.128094f
C5007 por_ana_0.ibias_gen_0.vp0.n12 dvss 0.98287f
C5008 por_ana_0.ibias_gen_0.vp0.n13 dvss 1.07524f
C5009 por_ana_0.ibias_gen_0.vp0.n14 dvss 0.139118f
C5010 avdd.t615 dvss 0.874276f
C5011 avdd.n6 dvss 0.518139f
C5012 avdd.n12 dvss 0.26703f
C5013 avdd.n13 dvss 0.100963f
C5014 avdd.n14 dvss 0.948156f
C5015 avdd.t52 dvss 0.679404f
C5016 avdd.n15 dvss 0.421816f
C5017 avdd.n16 dvss 0.930405f
C5018 avdd.n17 dvss 0.556102f
C5019 avdd.n18 dvss 1.83502f
C5020 avdd.n19 dvss 1.83502f
C5021 avdd.n20 dvss 0.556102f
C5022 avdd.n21 dvss 0.930838f
C5023 avdd.n23 dvss 0.275544f
C5024 avdd.t619 dvss 0.436501f
C5025 avdd.n30 dvss 0.164106f
C5026 avdd.n31 dvss 0.726045f
C5027 avdd.n32 dvss 0.721072f
C5028 avdd.t503 dvss 0.159133f
C5029 avdd.t572 dvss 0.159133f
C5030 avdd.n41 dvss 0.26703f
C5031 avdd.n43 dvss 0.183998f
C5032 avdd.n49 dvss 0.164106f
C5033 avdd.n51 dvss 0.726045f
C5034 avdd.n52 dvss 0.721072f
C5035 avdd.t473 dvss 0.159133f
C5036 avdd.t518 dvss 0.159133f
C5037 avdd.n61 dvss 0.26703f
C5038 avdd.n63 dvss 0.183998f
C5039 avdd.n69 dvss 0.164106f
C5040 avdd.n71 dvss 0.726045f
C5041 avdd.n72 dvss 0.721072f
C5042 avdd.t435 dvss 0.159133f
C5043 avdd.t592 dvss 0.159133f
C5044 avdd.n81 dvss 0.26703f
C5045 avdd.n83 dvss 0.183998f
C5046 avdd.n89 dvss 0.164106f
C5047 avdd.n91 dvss 0.726045f
C5048 avdd.n92 dvss 0.721072f
C5049 avdd.t600 dvss 0.159133f
C5050 avdd.t449 dvss 0.159133f
C5051 avdd.n101 dvss 0.26703f
C5052 avdd.n103 dvss 0.183998f
C5053 avdd.n109 dvss 0.164106f
C5054 avdd.n111 dvss 0.726045f
C5055 avdd.n112 dvss 0.721072f
C5056 avdd.t258 dvss 0.159133f
C5057 avdd.t507 dvss 0.569672f
C5058 avdd.n121 dvss 0.26703f
C5059 avdd.n123 dvss 0.183998f
C5060 avdd.n124 dvss 0.193042f
C5061 avdd.n125 dvss 0.139218f
C5062 avdd.n127 dvss 0.26703f
C5063 avdd.n133 dvss 0.721072f
C5064 avdd.n134 dvss 0.726045f
C5065 avdd.n135 dvss 0.164106f
C5066 avdd.n139 dvss 0.183998f
C5067 avdd.n140 dvss 0.26703f
C5068 avdd.n145 dvss 0.726045f
C5069 avdd.n146 dvss 0.164106f
C5070 avdd.t0 dvss 0.159133f
C5071 avdd.n147 dvss 0.721072f
C5072 avdd.n150 dvss 0.183998f
C5073 avdd.n152 dvss 0.26703f
C5074 avdd.n158 dvss 0.721072f
C5075 avdd.n159 dvss 0.726045f
C5076 avdd.n160 dvss 0.164106f
C5077 avdd.n164 dvss 0.183998f
C5078 avdd.n165 dvss 0.26703f
C5079 avdd.n170 dvss 0.726045f
C5080 avdd.n171 dvss 0.164106f
C5081 avdd.t466 dvss 0.159133f
C5082 avdd.n172 dvss 0.721072f
C5083 avdd.n175 dvss 0.183998f
C5084 avdd.n177 dvss 0.26703f
C5085 avdd.n183 dvss 0.721072f
C5086 avdd.n184 dvss 0.726045f
C5087 avdd.n185 dvss 0.164106f
C5088 avdd.n189 dvss 0.183998f
C5089 avdd.n190 dvss 0.26703f
C5090 avdd.n195 dvss 0.726045f
C5091 avdd.n196 dvss 0.164106f
C5092 avdd.t423 dvss 0.159133f
C5093 avdd.n197 dvss 0.721072f
C5094 avdd.n200 dvss 0.183998f
C5095 avdd.n202 dvss 0.26703f
C5096 avdd.n208 dvss 0.721072f
C5097 avdd.n209 dvss 0.726045f
C5098 avdd.n210 dvss 0.164106f
C5099 avdd.n214 dvss 0.183998f
C5100 avdd.n215 dvss 0.26703f
C5101 avdd.n220 dvss 0.726045f
C5102 avdd.n221 dvss 0.164106f
C5103 avdd.t178 dvss 0.159133f
C5104 avdd.n222 dvss 0.721072f
C5105 avdd.n225 dvss 0.183998f
C5106 avdd.n227 dvss 0.26703f
C5107 avdd.n233 dvss 0.721072f
C5108 avdd.n234 dvss 0.726045f
C5109 avdd.n235 dvss 0.164106f
C5110 avdd.n239 dvss 0.183998f
C5111 avdd.n240 dvss 0.26703f
C5112 avdd.n245 dvss 0.726045f
C5113 avdd.n246 dvss 0.164106f
C5114 avdd.t390 dvss 0.159133f
C5115 avdd.n247 dvss 0.721072f
C5116 avdd.n250 dvss 0.183998f
C5117 avdd.n251 dvss 0.26703f
C5118 avdd.n257 dvss 0.902642f
C5119 avdd.t170 dvss 0.679404f
C5120 avdd.t39 dvss 0.679404f
C5121 avdd.t15 dvss 0.679404f
C5122 avdd.t72 dvss 0.679404f
C5123 avdd.t168 dvss 0.679404f
C5124 avdd.t156 dvss 0.679404f
C5125 avdd.t105 dvss 0.679404f
C5126 avdd.t37 dvss 0.679404f
C5127 avdd.t140 dvss 0.679404f
C5128 avdd.t66 dvss 0.679404f
C5129 avdd.t163 dvss 0.679404f
C5130 avdd.t117 dvss 0.679404f
C5131 avdd.t30 dvss 0.679404f
C5132 avdd.t98 dvss 0.679404f
C5133 avdd.n258 dvss 0.422925f
C5134 avdd.n259 dvss 0.422925f
C5135 avdd.n260 dvss 0.422925f
C5136 avdd.n261 dvss 0.422925f
C5137 avdd.n262 dvss 0.422925f
C5138 avdd.n263 dvss 0.422925f
C5139 avdd.n264 dvss 0.33011f
C5140 avdd.n266 dvss 0.417008f
C5141 avdd.n267 dvss 0.422925f
C5142 avdd.n268 dvss 0.422925f
C5143 avdd.n269 dvss 0.422925f
C5144 avdd.n270 dvss 0.422925f
C5145 avdd.n271 dvss 0.422925f
C5146 avdd.n272 dvss 0.434367f
C5147 avdd.n273 dvss 0.268917f
C5148 avdd.n274 dvss 2.17899f
C5149 avdd.n275 dvss 2.06497f
C5150 avdd.n276 dvss 12.359f
C5151 avdd.n277 dvss 0.718841f
C5152 avdd.n278 dvss 2.38231f
C5153 avdd.t49 dvss 2.50826f
C5154 avdd.n279 dvss 1.21434f
C5155 avdd.n280 dvss 0.186305f
C5156 avdd.n281 dvss 0.559858f
C5157 avdd.n282 dvss 0.166369f
C5158 avdd.n283 dvss 1.17335f
C5159 avdd.n284 dvss 1.24561f
C5160 avdd.n285 dvss 1.9778f
C5161 avdd.t3 dvss 42.410603f
C5162 avdd.n286 dvss 0.492917f
C5163 avdd.n287 dvss 2.37029f
C5164 avdd.n288 dvss 2.18197f
C5165 avdd.n289 dvss 1.34674f
C5166 avdd.n290 dvss 1.28101f
C5167 avdd.n291 dvss 0.172764f
C5168 avdd.n292 dvss 0.231603f
C5169 avdd.n293 dvss 0.392912f
C5170 avdd.n294 dvss 0.13548f
C5171 avdd.n295 dvss 0.146163f
C5172 avdd.t522 dvss 1.16861f
C5173 avdd.t574 dvss 1.61731f
C5174 avdd.n296 dvss 1.43163f
C5175 avdd.n297 dvss 0.392912f
C5176 avdd.t524 dvss 1.33066f
C5177 avdd.t520 dvss 1.46384f
C5178 avdd.n298 dvss 1.261f
C5179 avdd.n299 dvss 0.146163f
C5180 avdd.n300 dvss 0.13548f
C5181 avdd.n301 dvss 0.108276f
C5182 avdd.n302 dvss 0.728774f
C5183 avdd.n303 dvss 1.87701f
C5184 avdd.n304 dvss 1.34674f
C5185 avdd.t182 dvss 40.2424f
C5186 avdd.t191 dvss 53.6565f
C5187 avdd.t195 dvss 40.2424f
C5188 avdd.n305 dvss 1.24561f
C5189 avdd.n306 dvss 0.559858f
C5190 avdd.n308 dvss 0.22607f
C5191 avdd.n309 dvss 1.68642f
C5192 avdd.n310 dvss 1.55976f
C5193 avdd.n311 dvss 0.880079f
C5194 avdd.n313 dvss 0.402259f
C5195 avdd.n315 dvss 0.250756f
C5196 avdd.n317 dvss 0.250756f
C5197 avdd.n319 dvss 0.285234f
C5198 avdd.n321 dvss 0.285234f
C5199 avdd.n323 dvss 0.250756f
C5200 avdd.n325 dvss 0.250756f
C5201 avdd.n327 dvss 0.250756f
C5202 avdd.n329 dvss 0.250756f
C5203 avdd.n331 dvss 0.250756f
C5204 avdd.n333 dvss 0.22607f
C5205 avdd.n334 dvss 0.100634f
C5206 avdd.n336 dvss 0.216493f
C5207 avdd.n337 dvss 2.25352f
C5208 avdd.n338 dvss 0.76996f
C5209 avdd.n339 dvss 0.855701f
C5210 avdd.n340 dvss 0.868137f
C5211 avdd.n341 dvss 3.69144f
C5212 avdd.n342 dvss 3.69097f
C5213 avdd.n343 dvss 13.9263f
C5214 avdd.n344 dvss 0.897212f
C5215 avdd.n345 dvss 0.867474f
C5216 avdd.n346 dvss 0.787913f
C5217 avdd.n347 dvss 1.57577f
C5218 avdd.n348 dvss 0.76996f
C5219 avdd.n349 dvss 1.34561f
C5220 avdd.n350 dvss 0.100634f
C5221 avdd.n351 dvss 0.124246f
C5222 avdd.n352 dvss 0.119114f
C5223 avdd.n353 dvss 0.111744f
C5224 avdd.n354 dvss 0.686022f
C5225 avdd.n355 dvss 2.4847f
C5226 avdd.n356 dvss 2.74167f
C5227 avdd.n357 dvss 2.47899f
C5228 avdd.n358 dvss 0.694691f
C5229 avdd.n359 dvss 0.145776f
C5230 avdd.n360 dvss 0.206471f
C5231 avdd.t477 dvss 0.61622f
C5232 avdd.n361 dvss 0.471201f
C5233 avdd.t489 dvss 0.61622f
C5234 avdd.t485 dvss 0.821627f
C5235 avdd.t487 dvss 0.821627f
C5236 avdd.t491 dvss 0.821627f
C5237 avdd.t481 dvss 1.01635f
C5238 avdd.n362 dvss 1.34589f
C5239 avdd.t483 dvss 0.821627f
C5240 avdd.t479 dvss 0.821627f
C5241 avdd.t501 dvss 0.821627f
C5242 avdd.t499 dvss 1.01635f
C5243 avdd.n363 dvss 1.34589f
C5244 avdd.n364 dvss 0.164257f
C5245 avdd.n365 dvss 0.15095f
C5246 avdd.n366 dvss 0.277707f
C5247 avdd.n367 dvss 0.15095f
C5248 avdd.n369 dvss 0.250756f
C5249 avdd.n371 dvss 0.250756f
C5250 avdd.n373 dvss 0.250756f
C5251 avdd.n375 dvss 0.250756f
C5252 avdd.n377 dvss 0.250756f
C5253 avdd.n379 dvss 0.285234f
C5254 avdd.n381 dvss 0.285234f
C5255 avdd.n383 dvss 0.250756f
C5256 avdd.n385 dvss 0.250756f
C5257 avdd.n387 dvss 0.402259f
C5258 avdd.n388 dvss 3.16454f
C5259 avdd.n389 dvss 2.38231f
C5260 avdd.n390 dvss 0.148932f
C5261 avdd.n391 dvss 0.285234f
C5262 avdd.t77 dvss 2.49356f
C5263 avdd.n392 dvss 0.148932f
C5264 avdd.n393 dvss 0.250756f
C5265 avdd.t54 dvss 2.49417f
C5266 avdd.n394 dvss 0.148932f
C5267 avdd.t144 dvss 2.49417f
C5268 avdd.n395 dvss 1.2293f
C5269 avdd.n397 dvss 0.22607f
C5270 avdd.t146 dvss 2.49417f
C5271 avdd.n398 dvss 1.2293f
C5272 avdd.n400 dvss 0.250756f
C5273 avdd.n401 dvss 0.250756f
C5274 avdd.t41 dvss 2.49417f
C5275 avdd.n403 dvss 1.2293f
C5276 avdd.n404 dvss 0.148932f
C5277 avdd.t12 dvss 2.49417f
C5278 avdd.n406 dvss 1.2293f
C5279 avdd.n407 dvss 0.148932f
C5280 avdd.n408 dvss 0.148932f
C5281 avdd.n409 dvss 1.2293f
C5282 avdd.n411 dvss 0.250756f
C5283 avdd.t47 dvss 2.49417f
C5284 avdd.n412 dvss 1.2293f
C5285 avdd.n414 dvss 0.250756f
C5286 avdd.n415 dvss 0.285234f
C5287 avdd.t61 dvss 2.49417f
C5288 avdd.n417 dvss 1.2293f
C5289 avdd.n418 dvss 0.183411f
C5290 avdd.t59 dvss 2.49356f
C5291 avdd.n420 dvss 1.22491f
C5292 avdd.n421 dvss 0.183411f
C5293 avdd.n422 dvss 0.148932f
C5294 avdd.n423 dvss 1.22491f
C5295 avdd.n425 dvss 0.250756f
C5296 avdd.t84 dvss 2.49356f
C5297 avdd.n426 dvss 1.22491f
C5298 avdd.n428 dvss 0.250756f
C5299 avdd.n429 dvss 0.402259f
C5300 avdd.t127 dvss 2.49356f
C5301 avdd.n431 dvss 1.22491f
C5302 avdd.n432 dvss 0.300435f
C5303 avdd.n433 dvss 1.75773f
C5304 avdd.n434 dvss 0.726183f
C5305 avdd.n435 dvss 0.211116f
C5306 avdd.n437 dvss 0.249373f
C5307 avdd.n439 dvss 0.249373f
C5308 avdd.n441 dvss 0.249373f
C5309 avdd.n443 dvss 0.249373f
C5310 avdd.n444 dvss 0.26803f
C5311 avdd.n445 dvss 0.165336f
C5312 avdd.n446 dvss 0.252782f
C5313 avdd.n447 dvss 0.471201f
C5314 avdd.n448 dvss 1.94802f
C5315 avdd.n449 dvss 0.492917f
C5316 avdd.t180 dvss 53.6565f
C5317 avdd.t13 dvss 42.410603f
C5318 avdd.n450 dvss 0.729577f
C5319 avdd.n451 dvss 1.24399f
C5320 avdd.n452 dvss 17.1196f
C5321 avdd.n453 dvss 1.04267f
C5322 avdd.n454 dvss 0.623909f
C5323 avdd.n455 dvss 0.190125f
C5324 avdd.n456 dvss 0.215937f
C5325 avdd.n457 dvss 0.100634f
C5326 avdd.n458 dvss 0.186305f
C5327 avdd.t68 dvss 2.50826f
C5328 avdd.n459 dvss 1.21434f
C5329 avdd.n461 dvss 0.694776f
C5330 avdd.n462 dvss 1.79115f
C5331 avdd.n463 dvss 2.19062f
C5332 avdd.n464 dvss 1.72069f
C5333 avdd.n465 dvss 0.839994f
C5334 avdd.n466 dvss 0.856753f
C5335 avdd.n467 dvss 3.70598f
C5336 avdd.n468 dvss 14.160501f
C5337 avdd.n469 dvss 13.9244f
C5338 avdd.n470 dvss 14.160501f
C5339 avdd.n471 dvss 3.70598f
C5340 avdd.n472 dvss 0.856245f
C5341 avdd.n473 dvss 0.829338f
C5342 avdd.n474 dvss 1.72069f
C5343 avdd.n475 dvss 1.5498f
C5344 avdd.n476 dvss 1.71222f
C5345 avdd.n477 dvss 0.557216f
C5346 avdd.n478 dvss 1.01478f
C5347 avdd.n479 dvss 1.6913f
C5348 avdd.n480 dvss 0.528888f
C5349 avdd.n482 dvss 0.209965f
C5350 avdd.n483 dvss 0.100634f
C5351 avdd.n484 dvss 0.739559f
C5352 avdd.n485 dvss 1.88884f
C5353 avdd.n486 dvss 26.8282f
C5354 avdd.n487 dvss 1.88884f
C5355 avdd.n488 dvss 1.10725f
C5356 avdd.n489 dvss 0.67404f
C5357 avdd.n490 dvss 0.729577f
C5358 avdd.n491 dvss 1.24399f
C5359 avdd.n492 dvss 17.1196f
C5360 avdd.n493 dvss 1.04267f
C5361 avdd.n494 dvss 0.623909f
C5362 avdd.n495 dvss 0.125419f
C5363 avdd.n496 dvss 0.215937f
C5364 avdd.n497 dvss 0.100634f
C5365 avdd.t124 dvss 2.49417f
C5366 avdd.n498 dvss 1.2293f
C5367 avdd.n499 dvss 0.124246f
C5368 avdd.t132 dvss 2.49417f
C5369 avdd.n500 dvss 1.2293f
C5370 avdd.n501 dvss 0.148932f
C5371 avdd.t165 dvss 2.49417f
C5372 avdd.n502 dvss 1.2293f
C5373 avdd.n503 dvss 0.148932f
C5374 avdd.t121 dvss 2.49417f
C5375 avdd.n504 dvss 1.2293f
C5376 avdd.n505 dvss 0.148932f
C5377 avdd.t2 dvss 2.49417f
C5378 avdd.n506 dvss 1.2293f
C5379 avdd.n507 dvss 0.148932f
C5380 avdd.t172 dvss 2.49417f
C5381 avdd.n508 dvss 1.2293f
C5382 avdd.n509 dvss 0.148932f
C5383 avdd.t9 dvss 2.49417f
C5384 avdd.n510 dvss 1.2293f
C5385 avdd.n511 dvss 0.183411f
C5386 avdd.t6 dvss 2.49356f
C5387 avdd.n512 dvss 1.22491f
C5388 avdd.n513 dvss 0.183411f
C5389 avdd.t17 dvss 2.49356f
C5390 avdd.n514 dvss 1.22491f
C5391 avdd.n515 dvss 0.148932f
C5392 avdd.t20 dvss 2.49356f
C5393 avdd.n516 dvss 1.22491f
C5394 avdd.n517 dvss 0.148932f
C5395 avdd.t56 dvss 2.49356f
C5396 avdd.n518 dvss 1.22491f
C5397 avdd.n519 dvss 0.300435f
C5398 avdd.n520 dvss 1.15566f
C5399 avdd.n521 dvss 0.451263f
C5400 avdd.n522 dvss 0.913885f
C5401 avdd.n523 dvss 0.676728f
C5402 avdd.n524 dvss 22.408098f
C5403 avdd.n525 dvss 91.0925f
C5404 avdd.n526 dvss 2.38231f
C5405 avdd.t129 dvss 2.50826f
C5406 avdd.n527 dvss 1.21434f
C5407 avdd.n528 dvss 0.186305f
C5408 avdd.n529 dvss 0.559858f
C5409 avdd.n530 dvss 0.166369f
C5410 avdd.n531 dvss 1.17335f
C5411 avdd.n532 dvss 1.24561f
C5412 avdd.n533 dvss 1.9778f
C5413 avdd.t27 dvss 42.410603f
C5414 avdd.n534 dvss 0.492917f
C5415 avdd.n535 dvss 2.37029f
C5416 avdd.n536 dvss 2.18197f
C5417 avdd.n537 dvss 1.34674f
C5418 avdd.n538 dvss 1.28101f
C5419 avdd.n539 dvss 0.172764f
C5420 avdd.n540 dvss 0.231603f
C5421 avdd.n541 dvss 0.392912f
C5422 avdd.n542 dvss 0.13548f
C5423 avdd.n543 dvss 0.146163f
C5424 avdd.t607 dvss 1.16861f
C5425 avdd.t460 dvss 1.61731f
C5426 avdd.n544 dvss 1.43163f
C5427 avdd.n545 dvss 0.392912f
C5428 avdd.t609 dvss 1.33066f
C5429 avdd.t605 dvss 1.46384f
C5430 avdd.n546 dvss 1.261f
C5431 avdd.n547 dvss 0.146163f
C5432 avdd.n548 dvss 0.13548f
C5433 avdd.n549 dvss 0.108276f
C5434 avdd.n550 dvss 0.728774f
C5435 avdd.n551 dvss 1.87701f
C5436 avdd.n552 dvss 1.34674f
C5437 avdd.t403 dvss 40.2424f
C5438 avdd.t395 dvss 53.6565f
C5439 avdd.t392 dvss 40.2424f
C5440 avdd.n553 dvss 1.24561f
C5441 avdd.n554 dvss 0.559858f
C5442 avdd.n556 dvss 0.22607f
C5443 avdd.n557 dvss 1.68642f
C5444 avdd.n558 dvss 1.55976f
C5445 avdd.n559 dvss 0.880079f
C5446 avdd.n561 dvss 0.402259f
C5447 avdd.n563 dvss 0.250756f
C5448 avdd.n565 dvss 0.250756f
C5449 avdd.n567 dvss 0.285234f
C5450 avdd.n569 dvss 0.285234f
C5451 avdd.n571 dvss 0.250756f
C5452 avdd.n573 dvss 0.250756f
C5453 avdd.n575 dvss 0.250756f
C5454 avdd.n577 dvss 0.250756f
C5455 avdd.n579 dvss 0.250756f
C5456 avdd.n581 dvss 0.22607f
C5457 avdd.n582 dvss 0.100634f
C5458 avdd.n584 dvss 0.216493f
C5459 avdd.n585 dvss 2.25352f
C5460 avdd.n586 dvss 0.76996f
C5461 avdd.n587 dvss 0.855701f
C5462 avdd.n588 dvss 0.868137f
C5463 avdd.n589 dvss 3.69144f
C5464 avdd.n590 dvss 3.69097f
C5465 avdd.n591 dvss 13.9263f
C5466 avdd.n592 dvss 0.897212f
C5467 avdd.n593 dvss 0.867474f
C5468 avdd.n594 dvss 0.787913f
C5469 avdd.n595 dvss 1.57577f
C5470 avdd.n596 dvss 0.76996f
C5471 avdd.n597 dvss 1.34561f
C5472 avdd.n598 dvss 0.100634f
C5473 avdd.n599 dvss 0.124246f
C5474 avdd.n600 dvss 0.119114f
C5475 avdd.n601 dvss 0.111744f
C5476 avdd.n602 dvss 0.686022f
C5477 avdd.n603 dvss 2.4847f
C5478 avdd.n604 dvss 2.74167f
C5479 avdd.n605 dvss 2.47899f
C5480 avdd.n606 dvss 0.694691f
C5481 avdd.n607 dvss 0.145776f
C5482 avdd.n608 dvss 0.206471f
C5483 avdd.t536 dvss 0.61622f
C5484 avdd.n609 dvss 0.471201f
C5485 avdd.t530 dvss 0.61622f
C5486 avdd.t538 dvss 0.821627f
C5487 avdd.t528 dvss 0.821627f
C5488 avdd.t532 dvss 0.821627f
C5489 avdd.t540 dvss 1.01635f
C5490 avdd.n610 dvss 1.34589f
C5491 avdd.t542 dvss 0.821627f
C5492 avdd.t534 dvss 0.821627f
C5493 avdd.t546 dvss 0.821627f
C5494 avdd.t544 dvss 1.01635f
C5495 avdd.n611 dvss 1.34589f
C5496 avdd.n612 dvss 0.164257f
C5497 avdd.n613 dvss 0.15095f
C5498 avdd.n614 dvss 0.277707f
C5499 avdd.n615 dvss 0.15095f
C5500 avdd.t274 dvss 0.159133f
C5501 avdd.t278 dvss 0.159133f
C5502 avdd.t344 dvss 0.159133f
C5503 avdd.t340 dvss 0.159133f
C5504 avdd.n640 dvss 0.165764f
C5505 avdd.t324 dvss 0.159133f
C5506 avdd.n651 dvss 0.185655f
C5507 avdd.t350 dvss 0.159133f
C5508 avdd.n662 dvss 0.205547f
C5509 avdd.t352 dvss 0.368443f
C5510 avdd.n667 dvss 0.504724f
C5511 avdd.n668 dvss 0.144996f
C5512 avdd.n673 dvss 0.212178f
C5513 avdd.t348 dvss 0.159133f
C5514 avdd.n674 dvss 0.258591f
C5515 avdd.t322 dvss 0.159133f
C5516 avdd.n675 dvss 0.251961f
C5517 avdd.n676 dvss 0.165764f
C5518 avdd.n684 dvss 0.225439f
C5519 avdd.n685 dvss 0.192286f
C5520 avdd.t328 dvss 0.159133f
C5521 avdd.t330 dvss 0.159133f
C5522 avdd.n686 dvss 0.258591f
C5523 avdd.n694 dvss 0.232069f
C5524 avdd.t336 dvss 0.159133f
C5525 avdd.n695 dvss 0.24533f
C5526 avdd.n696 dvss 0.258591f
C5527 avdd.t338 dvss 0.159133f
C5528 avdd.n697 dvss 0.172394f
C5529 avdd.n705 dvss 0.205547f
C5530 avdd.n706 dvss 0.212178f
C5531 avdd.t346 dvss 0.159133f
C5532 avdd.t326 dvss 0.159133f
C5533 avdd.n707 dvss 0.258591f
C5534 avdd.n715 dvss 0.251961f
C5535 avdd.t332 dvss 0.159133f
C5536 avdd.n716 dvss 0.225439f
C5537 avdd.n717 dvss 0.258591f
C5538 avdd.t334 dvss 0.159133f
C5539 avdd.n718 dvss 0.192286f
C5540 avdd.n726 dvss 0.185655f
C5541 avdd.n727 dvss 0.232069f
C5542 avdd.t342 dvss 0.159133f
C5543 avdd.n728 dvss 0.172394f
C5544 avdd.n729 dvss 0.24533f
C5545 avdd.n737 dvss 0.305005f
C5546 avdd.n738 dvss 0.306663f
C5547 avdd.t280 dvss 0.159133f
C5548 avdd.n739 dvss 0.246988f
C5549 avdd.n740 dvss 0.170737f
C5550 avdd.n752 dvss 0.885361f
C5551 avdd.n753 dvss 0.487438f
C5552 avdd.n754 dvss 0.487438f
C5553 avdd.n755 dvss 0.487438f
C5554 avdd.n756 dvss 0.487438f
C5555 avdd.n757 dvss 0.487438f
C5556 avdd.n758 dvss 0.480812f
C5557 avdd.n759 dvss 0.32463f
C5558 avdd.n760 dvss 0.331226f
C5559 avdd.n762 dvss 0.444821f
C5560 avdd.n763 dvss 0.167175f
C5561 avdd.n769 dvss 0.230412f
C5562 avdd.n770 dvss 0.187313f
C5563 avdd.t276 dvss 0.159133f
C5564 avdd.n771 dvss 0.258591f
C5565 avdd.n774 dvss 0.190628f
C5566 avdd.n775 dvss 0.318266f
C5567 avdd.n776 dvss 0.313293f
C5568 avdd.t443 dvss 0.569672f
C5569 avdd.n777 dvss 0.193042f
C5570 avdd.n778 dvss 0.139218f
C5571 avdd.n786 dvss 0.324733f
C5572 avdd.n788 dvss 0.26703f
C5573 avdd.n790 dvss 1.73653f
C5574 avdd.n792 dvss 0.250756f
C5575 avdd.n794 dvss 0.250756f
C5576 avdd.n796 dvss 0.250756f
C5577 avdd.n798 dvss 0.250756f
C5578 avdd.n800 dvss 0.250756f
C5579 avdd.n802 dvss 0.285234f
C5580 avdd.n804 dvss 0.285234f
C5581 avdd.n806 dvss 0.250756f
C5582 avdd.n808 dvss 0.250756f
C5583 avdd.n810 dvss 0.402259f
C5584 avdd.n811 dvss 3.16454f
C5585 avdd.n812 dvss 2.38231f
C5586 avdd.n813 dvss 0.148932f
C5587 avdd.n814 dvss 0.285234f
C5588 avdd.t151 dvss 2.49356f
C5589 avdd.n815 dvss 0.148932f
C5590 avdd.n816 dvss 0.250756f
C5591 avdd.t94 dvss 2.49417f
C5592 avdd.n817 dvss 0.148932f
C5593 avdd.t70 dvss 2.49417f
C5594 avdd.n818 dvss 1.2293f
C5595 avdd.n820 dvss 0.22607f
C5596 avdd.t32 dvss 2.49417f
C5597 avdd.n821 dvss 1.2293f
C5598 avdd.n823 dvss 0.250756f
C5599 avdd.n824 dvss 0.250756f
C5600 avdd.t82 dvss 2.49417f
C5601 avdd.n826 dvss 1.2293f
C5602 avdd.n827 dvss 0.148932f
C5603 avdd.t86 dvss 2.49417f
C5604 avdd.n829 dvss 1.2293f
C5605 avdd.n830 dvss 0.148932f
C5606 avdd.n831 dvss 0.148932f
C5607 avdd.n832 dvss 1.2293f
C5608 avdd.n834 dvss 0.250756f
C5609 avdd.t96 dvss 2.49417f
C5610 avdd.n835 dvss 1.2293f
C5611 avdd.n837 dvss 0.250756f
C5612 avdd.n838 dvss 0.285234f
C5613 avdd.t142 dvss 2.49417f
C5614 avdd.n840 dvss 1.2293f
C5615 avdd.n841 dvss 0.183411f
C5616 avdd.t103 dvss 2.49356f
C5617 avdd.n843 dvss 1.22491f
C5618 avdd.n844 dvss 0.183411f
C5619 avdd.n845 dvss 0.148932f
C5620 avdd.n846 dvss 1.22491f
C5621 avdd.n848 dvss 0.250756f
C5622 avdd.t112 dvss 2.49356f
C5623 avdd.n849 dvss 1.22491f
C5624 avdd.n851 dvss 0.250756f
C5625 avdd.n852 dvss 0.402259f
C5626 avdd.t158 dvss 2.49356f
C5627 avdd.n854 dvss 1.22491f
C5628 avdd.n855 dvss 0.300435f
C5629 avdd.n856 dvss 1.14292f
C5630 avdd.n857 dvss 4.99779f
C5631 avdd.n858 dvss 0.70867f
C5632 avdd.n859 dvss 0.211116f
C5633 avdd.n861 dvss 0.249373f
C5634 avdd.n863 dvss 0.249373f
C5635 avdd.n865 dvss 0.249373f
C5636 avdd.n867 dvss 0.249373f
C5637 avdd.n868 dvss 0.26803f
C5638 avdd.n869 dvss 0.165336f
C5639 avdd.n870 dvss 0.252782f
C5640 avdd.n871 dvss 0.471201f
C5641 avdd.n872 dvss 1.94802f
C5642 avdd.n873 dvss 0.492917f
C5643 avdd.t401 dvss 53.6565f
C5644 avdd.t33 dvss 42.410603f
C5645 avdd.n874 dvss 0.729577f
C5646 avdd.n875 dvss 1.24399f
C5647 avdd.n876 dvss 17.1196f
C5648 avdd.n877 dvss 1.04267f
C5649 avdd.n878 dvss 0.623909f
C5650 avdd.n879 dvss 0.190125f
C5651 avdd.n880 dvss 0.215937f
C5652 avdd.n881 dvss 0.100634f
C5653 avdd.n882 dvss 0.186305f
C5654 avdd.t135 dvss 2.50826f
C5655 avdd.n883 dvss 1.21434f
C5656 avdd.n885 dvss 0.694776f
C5657 avdd.n886 dvss 1.79115f
C5658 avdd.n887 dvss 2.19062f
C5659 avdd.n888 dvss 1.72069f
C5660 avdd.n889 dvss 0.839994f
C5661 avdd.n890 dvss 0.856753f
C5662 avdd.n891 dvss 3.70598f
C5663 avdd.n892 dvss 14.160501f
C5664 avdd.n893 dvss 13.9244f
C5665 avdd.n894 dvss 14.160501f
C5666 avdd.n895 dvss 3.70598f
C5667 avdd.n896 dvss 0.856245f
C5668 avdd.n897 dvss 0.829338f
C5669 avdd.n898 dvss 1.72069f
C5670 avdd.n899 dvss 1.5498f
C5671 avdd.n900 dvss 1.71222f
C5672 avdd.n901 dvss 0.557216f
C5673 avdd.n902 dvss 1.01478f
C5674 avdd.n903 dvss 1.6913f
C5675 avdd.n904 dvss 0.528888f
C5676 avdd.n906 dvss 0.209965f
C5677 avdd.n907 dvss 0.100634f
C5678 avdd.n908 dvss 0.739559f
C5679 avdd.n909 dvss 1.88884f
C5680 avdd.n910 dvss 26.8282f
C5681 avdd.n911 dvss 1.88884f
C5682 avdd.n912 dvss 1.10725f
C5683 avdd.n913 dvss 0.67404f
C5684 avdd.n914 dvss 0.729577f
C5685 avdd.n915 dvss 1.24399f
C5686 avdd.n916 dvss 17.1196f
C5687 avdd.n917 dvss 1.04267f
C5688 avdd.n918 dvss 0.623909f
C5689 avdd.n919 dvss 0.125419f
C5690 avdd.n920 dvss 0.215937f
C5691 avdd.n921 dvss 0.100634f
C5692 avdd.t63 dvss 2.49417f
C5693 avdd.n922 dvss 1.2293f
C5694 avdd.n923 dvss 0.124246f
C5695 avdd.t26 dvss 2.49417f
C5696 avdd.n924 dvss 1.2293f
C5697 avdd.n925 dvss 0.148932f
C5698 avdd.t74 dvss 2.49417f
C5699 avdd.n926 dvss 1.2293f
C5700 avdd.n927 dvss 0.148932f
C5701 avdd.t79 dvss 2.49417f
C5702 avdd.n928 dvss 1.2293f
C5703 avdd.n929 dvss 0.148932f
C5704 avdd.t88 dvss 2.49417f
C5705 avdd.n930 dvss 1.2293f
C5706 avdd.n931 dvss 0.148932f
C5707 avdd.t91 dvss 2.49417f
C5708 avdd.n932 dvss 1.2293f
C5709 avdd.n933 dvss 0.148932f
C5710 avdd.t137 dvss 2.49417f
C5711 avdd.n934 dvss 1.2293f
C5712 avdd.n935 dvss 0.183411f
C5713 avdd.t100 dvss 2.49356f
C5714 avdd.n936 dvss 1.22491f
C5715 avdd.n937 dvss 0.183411f
C5716 avdd.t148 dvss 2.49356f
C5717 avdd.n938 dvss 1.22491f
C5718 avdd.n939 dvss 0.148932f
C5719 avdd.t109 dvss 2.49356f
C5720 avdd.n940 dvss 1.22491f
C5721 avdd.n941 dvss 0.148932f
C5722 avdd.t153 dvss 2.49356f
C5723 avdd.n942 dvss 1.22491f
C5724 avdd.n943 dvss 0.300435f
C5725 avdd.n944 dvss 1.15566f
C5726 avdd.n945 dvss 0.451263f
C5727 avdd.n946 dvss 0.913885f
C5728 avdd.n947 dvss 0.676728f
C5729 avdd.n948 dvss 2.79605f
C5730 avdd.n949 dvss 4.54006f
C5731 avdd.n950 dvss 2.59963f
C5732 avdd.n951 dvss 1.68087f
C5733 avdd.n952 dvss 11.4123f
C5734 avdd.n953 dvss 8.03533f
C5735 avdd.n954 dvss 43.8503f
C5736 avdd.n955 dvss 37.4434f
C5737 avdd.n956 dvss 3.83384f
C5738 avdd.n957 dvss 4.10081f
C5739 avdd.n958 dvss 0.92979f
C5740 avdd.n959 dvss 5.68455f
C5741 avdd.n960 dvss 2.00459f
C5742 avdd.n961 dvss 7.69575f
C5743 avdd.n962 dvss 12.6061f
C5744 avdd.n963 dvss 3.23933f
C5745 avdd.n964 dvss 0.57311f
C5746 avdd.n965 dvss 1.53187f
C5747 avdd.n966 dvss 6.22696f
C5748 avdd.n967 dvss 1.24963f
C5749 avdd.n968 dvss 6.95338f
C5750 avdd.n969 dvss 1.94924f
C5751 avdd.n970 dvss 1.9502f
C5752 avdd.n971 dvss 23.895699f
C5753 avdd.n972 dvss 6.23715f
C5754 avdd.n973 dvss 0.912934f
C5755 avdd.n974 dvss 0.916912f
C5756 avdd.n975 dvss 3.25426f
C5757 avdd.n976 dvss 1.3951f
C5758 avdd.n977 dvss 76.9928f
C5759 avdd.n978 dvss 0.601892f
C5760 avdd.n982 dvss 0.127422f
C5761 avdd.t292 dvss 1.73f
C5762 avdd.t307 dvss 0.708015f
C5763 avdd.t431 dvss 1.15646f
C5764 avdd.n1004 dvss 1.03159f
C5765 avdd.t286 dvss 1.73f
C5766 avdd.t288 dvss 0.708015f
C5767 avdd.t505 dvss 1.15646f
C5768 avdd.n1025 dvss 1.03159f
C5769 avdd.t556 dvss 1.73f
C5770 avdd.t588 dvss 0.708015f
C5771 avdd.t270 dvss 1.15646f
C5772 avdd.n1046 dvss 1.03159f
C5773 avdd.t419 dvss 1.73f
C5774 avdd.t421 dvss 0.708015f
C5775 avdd.t475 dvss 1.15646f
C5776 avdd.n1067 dvss 1.03159f
C5777 avdd.t317 dvss 1.73f
C5778 avdd.t315 dvss 0.708015f
C5779 avdd.t320 dvss 1.15646f
C5780 avdd.n1088 dvss 1.03159f
C5781 avdd.t302 dvss 1.73f
C5782 avdd.t300 dvss 0.708015f
C5783 avdd.t212 dvss 1.15646f
C5784 avdd.n1109 dvss 1.03159f
C5785 avdd.t453 dvss 1.73f
C5786 avdd.t512 dvss 0.708015f
C5787 avdd.t264 dvss 1.15646f
C5788 avdd.n1130 dvss 1.03159f
C5789 avdd.t298 dvss 1.73f
C5790 avdd.t296 dvss 0.708015f
C5791 avdd.t461 dvss 1.15646f
C5792 avdd.n1151 dvss 1.03159f
C5793 avdd.t445 dvss 1.56819f
C5794 avdd.t657 dvss 0.641792f
C5795 avdd.t216 dvss 1.09623f
C5796 avdd.n1166 dvss 1.34401f
C5797 avdd.n1175 dvss 0.194978f
C5798 avdd.n1181 dvss 0.935098f
C5799 avdd.n1193 dvss 9.62448f
C5800 avdd.n1194 dvss 5.78011f
C5801 avdd.n1203 dvss 0.194978f
C5802 avdd.n1209 dvss 1.21613f
C5803 avdd.n1218 dvss 0.194978f
C5804 avdd.n1224 dvss 1.21613f
C5805 avdd.n1233 dvss 0.194978f
C5806 avdd.n1239 dvss 1.21613f
C5807 avdd.n1248 dvss 0.194978f
C5808 avdd.n1254 dvss 1.21613f
C5809 avdd.n1263 dvss 0.194978f
C5810 avdd.n1269 dvss 1.21613f
C5811 avdd.n1278 dvss 0.194978f
C5812 avdd.n1284 dvss 1.21613f
C5813 avdd.n1293 dvss 0.194978f
C5814 avdd.n1299 dvss 1.21613f
C5815 avdd.n1308 dvss 0.194978f
C5816 avdd.n1314 dvss 1.21613f
C5817 avdd.t311 dvss 1.21817f
C5818 avdd.n1320 dvss 0.563133f
C5819 avdd.n1322 dvss 0.437355f
C5820 avdd.t294 dvss 0.231967f
C5821 avdd.n1323 dvss 0.258547f
C5822 avdd.n1324 dvss 0.372114f
C5823 avdd.t439 dvss 0.231967f
C5824 avdd.n1326 dvss 0.323788f
C5825 avdd.n1327 dvss 0.463934f
C5826 avdd.t441 dvss 1.13567f
C5827 avdd.t655 dvss 0.207804f
C5828 avdd.n1328 dvss 0.42044f
C5829 avdd.n1339 dvss 0.194978f
C5830 avdd.n1349 dvss 1.04718f
C5831 avdd.n1350 dvss 2.11501f
C5832 avdd.n1351 dvss 49.638897f
C5833 avdd.n1355 dvss 0.127422f
C5834 avdd.t210 dvss 1.73f
C5835 avdd.t208 dvss 0.708015f
C5836 avdd.t494 dvss 1.15646f
C5837 avdd.n1377 dvss 1.03159f
C5838 avdd.t268 dvss 1.73f
C5839 avdd.t266 dvss 0.708015f
C5840 avdd.t515 dvss 1.15646f
C5841 avdd.n1398 dvss 1.03159f
C5842 avdd.t254 dvss 1.73f
C5843 avdd.t256 dvss 0.708015f
C5844 avdd.t262 dvss 1.15646f
C5845 avdd.n1419 dvss 1.03159f
C5846 avdd.t284 dvss 1.73f
C5847 avdd.t282 dvss 0.708015f
C5848 avdd.t456 dvss 1.15646f
C5849 avdd.n1440 dvss 1.03159f
C5850 avdd.t565 dvss 1.73f
C5851 avdd.t567 dvss 0.708015f
C5852 avdd.t651 dvss 1.15646f
C5853 avdd.n1461 dvss 1.03159f
C5854 avdd.t313 dvss 1.73f
C5855 avdd.t563 dvss 0.708015f
C5856 avdd.t437 dvss 1.15646f
C5857 avdd.n1482 dvss 1.03159f
C5858 avdd.t596 dvss 1.73f
C5859 avdd.t598 dvss 0.708015f
C5860 avdd.t304 dvss 1.15646f
C5861 avdd.n1503 dvss 1.03159f
C5862 avdd.t309 dvss 1.73f
C5863 avdd.t510 dvss 0.708015f
C5864 avdd.t427 dvss 1.15646f
C5865 avdd.n1524 dvss 1.03159f
C5866 avdd.n1540 dvss 0.194978f
C5867 avdd.n1546 dvss 1.21613f
C5868 avdd.n1555 dvss 0.194978f
C5869 avdd.n1561 dvss 1.21613f
C5870 avdd.n1570 dvss 0.194978f
C5871 avdd.n1576 dvss 1.21613f
C5872 avdd.n1585 dvss 0.194978f
C5873 avdd.n1591 dvss 1.21613f
C5874 avdd.n1600 dvss 0.194978f
C5875 avdd.n1606 dvss 1.21613f
C5876 avdd.n1615 dvss 0.194978f
C5877 avdd.n1621 dvss 1.21613f
C5878 avdd.n1630 dvss 0.194978f
C5879 avdd.n1636 dvss 1.21613f
C5880 avdd.n1645 dvss 0.194978f
C5881 avdd.n1651 dvss 1.21613f
C5882 avdd.t272 dvss 1.2179f
C5883 avdd.n1657 dvss 0.560242f
C5884 avdd.n1659 dvss 0.434938f
C5885 avdd.t447 dvss 0.231967f
C5886 avdd.n1660 dvss 0.258547f
C5887 avdd.n1661 dvss 0.372114f
C5888 avdd.t252 dvss 0.231967f
C5889 avdd.n1663 dvss 0.323788f
C5890 avdd.n1664 dvss 0.463934f
C5891 avdd.t250 dvss 1.13567f
C5892 avdd.t497 dvss 0.207804f
C5893 avdd.n1665 dvss 0.42044f
C5894 avdd.n1676 dvss 0.194978f
C5895 avdd.n1686 dvss 1.07109f
C5896 avdd.n1687 dvss 0.907343f
C5897 avdd.n1689 dvss 1.05965f
C5898 avdd.n1690 dvss 5.4861f
C5899 avdd.n1691 dvss 19.7417f
C5900 avdd.n1692 dvss 64.6072f
C5901 avdd.n1693 dvss 81.356895f
C5902 avdd.n1694 dvss 82.178f
C5903 avdd.n1695 dvss 13.1971f
C5904 avdd.n1696 dvss 4.37046f
C5905 avdd.n1697 dvss 4.58552f
C5906 avdd.n1698 dvss 3.22329f
C5907 avdd.n1699 dvss 1.53528f
C5908 avdd.n1700 dvss 0.574676f
C5909 avdd.n1701 dvss 4.59175f
C5910 avdd.n1702 dvss 18.0441f
C5911 avdd.n1703 dvss 29.661901f
C5912 avdd.n1704 dvss 36.610397f
C5913 avdd.n1705 dvss 8.840321f
C5914 avdd.n1706 dvss 2.00388f
C5915 avdd.n1707 dvss 2.32847f
C5916 avdd.n1708 dvss 9.42348f
C5917 avdd.n1709 dvss 8.79056f
C5918 avdd.n1710 dvss 4.62764f
C5919 avdd.n1711 dvss 2.12896f
C5920 avdd.n1712 dvss 1.41065f
C5921 avdd.n1713 dvss 5.09092f
C5922 avdd.n1714 dvss 5.87451f
C5923 avdd.n1715 dvss 0.932463f
C5924 avdd.n1716 dvss 1.78015f
C5925 avdd.n1717 dvss 4.59618f
C5926 avdd.n1718 dvss 23.7499f
C5927 avdd.n1719 dvss 30.798101f
C5928 avdd.n1720 dvss 50.564198f
C5929 avdd.n1721 dvss 13.167f
C5930 avdd.n1722 dvss 1.30391f
C5931 avdd.n1723 dvss 2.04239f
C5932 avdd.n1724 dvss 5.68061f
C5933 avdd.n1725 dvss 3.2828f
C5934 avdd.n1726 dvss 1.32364f
C5935 avdd.n1727 dvss 32.9243f
C5936 avdd.n1728 dvss 33.77f
C5937 avdd.n1729 dvss 7.82596f
C5938 avdd.n1730 dvss 1.7031f
C5939 avdd.n1731 dvss 0.234737f
C5940 avdd.n1732 dvss 0.524002f
C5941 avdd.n1733 dvss 1.30139f
C5942 avdd.n1734 dvss 1.21593f
C5943 avdd.n1735 dvss 0.190607f
C5944 avdd.n1736 dvss 0.254316f
C5945 avdd.n1737 dvss 0.533778f
C5946 avdd.n1738 dvss 0.607078f
C5947 avdd.t576 dvss 4.05139f
C5948 avdd.t621 dvss 2.0257f
C5949 avdd.n1739 dvss 0.533778f
C5950 avdd.n1741 dvss 0.269334f
C5951 avdd.n1742 dvss 0.457234f
C5952 avdd.t382 dvss 5.21218f
C5953 avdd.t108 dvss 4.05139f
C5954 avdd.t575 dvss 4.05139f
C5955 avdd.t571 dvss 2.73128f
C5956 avdd.t623 dvss 2.53781f
C5957 avdd.n1743 dvss 0.248862f
C5958 avdd.n1744 dvss 5.96329f
C5959 avdd.t584 dvss 7.93208f
C5960 avdd.t388 dvss 5.21218f
C5961 avdd.t603 dvss 6.62334f
C5962 avdd.n1745 dvss 0.457234f
C5963 avdd.n1746 dvss 1.34129f
C5964 avdd.t580 dvss 0.387358f
C5965 avdd.n1747 dvss 0.958909f
C5966 avdd.t618 dvss 0.387358f
C5967 avdd.n1748 dvss 0.835825f
C5968 avdd.t175 dvss 0.774121f
C5969 avdd.n1749 dvss 0.701673f
C5970 avdd.t119 dvss 0.774012f
C5971 avdd.n1750 dvss 0.83081f
C5972 avdd.t107 dvss 0.774012f
C5973 avdd.n1751 dvss 0.935075f
C5974 avdd.n1752 dvss 0.143179f
C5975 avdd.n1753 dvss 0.433701f
C5976 avdd.t585 dvss 0.387358f
C5977 avdd.n1754 dvss 0.903763f
C5978 avdd.n1755 dvss 0.236257f
C5979 avdd.n1756 dvss 1.23797f
C5980 avdd.n1757 dvss 0.236257f
C5981 avdd.n1758 dvss 1.08511f
C5982 avdd.n1759 dvss 0.439835f
C5983 avdd.n1760 dvss 0.143179f
C5984 avdd.n1761 dvss 0.256686f
C5985 avdd.t35 dvss 1.2519f
C5986 avdd.n1762 dvss 2.61106f
C5987 avdd.t579 dvss 2.789f
C5988 avdd.t577 dvss 7.2834f
C5989 avdd.t611 dvss 7.693089f
C5990 avdd.t161 dvss 4.13105f
C5991 avdd.n1764 dvss 0.248862f
C5992 avdd.n1765 dvss 4.64317f
C5993 avdd.t617 dvss 4.75697f
C5994 avdd.n1766 dvss 2.83847f
C5995 avdd.n1767 dvss 2.83847f
C5996 avdd.n1768 dvss 1.66517f
C5997 avdd.n1769 dvss 1.64767f
C5998 avdd.n1770 dvss 1.59572f
C5999 avdd.t583 dvss 3.09545f
C6000 avdd.t176 dvss 4.05139f
C6001 avdd.t581 dvss 4.05139f
C6002 avdd.t570 dvss 4.56351f
C6003 avdd.n1771 dvss 2.61747f
C6004 avdd.t386 dvss 5.81251f
C6005 avdd.t384 dvss 8.45503f
C6006 avdd.t378 dvss 6.539629f
C6007 avdd.n1772 dvss 4.35975f
C6008 avdd.t380 dvss 6.539629f
C6009 avdd.t24 dvss 8.719501f
C6010 avdd.t550 dvss 8.719501f
C6011 avdd.t548 dvss 8.719501f
C6012 avdd.t115 dvss 8.719501f
C6013 avdd.t552 dvss 8.719501f
C6014 avdd.t554 dvss 8.719501f
C6015 avdd.t44 dvss 7.33424f
C6016 avdd.n1773 dvss 6.56865f
C6017 avdd.n1774 dvss 0.849471f
C6018 avdd.n1775 dvss 0.856818f
C6019 avdd.n1776 dvss 2.58152f
C6020 avdd.t23 dvss 3.90696f
C6021 avdd.n1777 dvss 1.44336f
C6022 avdd.n1778 dvss 1.59688f
C6023 avdd.n1779 dvss 0.3183f
C6024 avdd.t46 dvss 0.342639f
C6025 avdd.t43 dvss 4.00344f
C6026 avdd.n1780 dvss 3.54837f
C6027 avdd.n1781 dvss 0.636365f
C6028 avdd.n1782 dvss 0.197548f
C6029 avdd.n1783 dvss 1.31001f
C6030 avdd.n1784 dvss 1.31001f
C6031 avdd.n1785 dvss 0.197548f
C6032 avdd.t116 dvss 0.18489f
C6033 avdd.n1786 dvss 0.190362f
C6034 avdd.t114 dvss 3.99625f
C6035 avdd.n1787 dvss 3.52291f
C6036 avdd.n1788 dvss 1.25595f
C6037 avdd.n1789 dvss 0.18831f
C6038 avdd.t25 dvss 0.18489f
C6039 avdd.n1790 dvss 0.197548f
C6040 avdd.n1791 dvss 1.31048f
C6041 avdd.n1792 dvss 0.901982f
C6042 avdd.n1793 dvss 0.149534f
C6043 avdd.n1794 dvss 1.58632f
C6044 avdd.n1795 dvss 1.42287f
C6045 avdd.n1796 dvss 1.57524f
C6046 avdd.n1797 dvss 0.197548f
C6047 avdd.n1798 dvss 1.24585f
C6048 avdd.n1799 dvss 0.197548f
C6049 avdd.n1800 dvss 1.7148f
C6050 avdd.n1801 dvss 0.197548f
C6051 avdd.n1802 dvss 1.7148f
C6052 avdd.n1803 dvss 1.31001f
C6053 avdd.n1804 dvss 0.197548f
C6054 avdd.t162 dvss 0.435084f
C6055 avdd.t160 dvss 4.00344f
C6056 avdd.n1805 dvss 3.54837f
C6057 avdd.n1806 dvss 0.633566f
C6058 avdd.n1807 dvss 2.9201f
C6059 avdd.n1808 dvss 0.856818f
C6060 avdd.n1809 dvss 0.849471f
C6061 avdd.n1810 dvss 2.85615f
C6062 avdd.n1811 dvss 2.9118f
C6063 avdd.n1812 dvss 0.189272f
C6064 avdd.n1813 dvss 0.323131f
C6065 avdd.t36 dvss 2.40668f
C6066 avdd.n1814 dvss 0.323131f
C6067 avdd.n1815 dvss 0.580797f
C6068 avdd.n1816 dvss 0.247983f
C6069 avdd.n1817 dvss 0.138623f
C6070 avdd.n1818 dvss 0.183494f
C6071 avdd.n1819 dvss 0.472949f
C6072 avdd.t613 dvss 8.35315f
C6073 avdd.n1820 dvss 0.472949f
C6074 avdd.n1821 dvss 0.183494f
C6075 avdd.n1822 dvss 0.138623f
C6076 avdd.n1823 dvss 0.269334f
C6077 avdd.n1824 dvss 0.278479f
C6078 avdd.n1825 dvss 0.474664f
C6079 avdd.t120 dvss 2.98164f
C6080 avdd.n1826 dvss 0.474664f
C6081 avdd.n1827 dvss 0.26288f
C6082 avdd.n1828 dvss 0.204892f
C6083 avdd.n1829 dvss 1.34038f
C6084 avdd.n1830 dvss 1.94501f
C6085 avdd.n1831 dvss 12.9194f
C6086 avdd.n1832 dvss 27.136301f
C6087 avdd.n1833 dvss 16.504f
C6088 avdd.t219 dvss 0.410625f
C6089 avdd.n1834 dvss 0.783103f
C6090 avdd.n1835 dvss 0.674999f
C6091 avdd.n1836 dvss 0.272332f
C6092 avdd.n1837 dvss 0.261614f
C6093 avdd.n1838 dvss 0.851961f
C6094 avdd.n1839 dvss 0.261614f
C6095 avdd.n1840 dvss 0.851961f
C6096 avdd.n1841 dvss 0.261614f
C6097 avdd.n1842 dvss 0.851961f
C6098 avdd.n1843 dvss 0.261614f
C6099 avdd.n1844 dvss 0.851961f
C6100 avdd.n1845 dvss 0.261614f
C6101 avdd.n1846 dvss 0.851961f
C6102 avdd.n1847 dvss 0.261614f
C6103 avdd.n1848 dvss 0.851961f
C6104 avdd.n1849 dvss 0.261614f
C6105 avdd.n1850 dvss 0.851961f
C6106 avdd.t247 dvss 0.410625f
C6107 avdd.n1851 dvss 0.908053f
C6108 avdd.n1852 dvss 0.891458f
C6109 avdd.n1853 dvss 0.279066f
C6110 avdd.n1854 dvss 0.818269f
C6111 avdd.n1855 dvss 0.272332f
C6112 avdd.n1856 dvss 0.394608f
C6113 avdd.n1857 dvss 0.818269f
C6114 avdd.n1858 dvss 2.688f
C6115 avdd.t218 dvss 2.09379f
C6116 avdd.t222 dvss 1.7295f
C6117 avdd.t248 dvss 1.7295f
C6118 avdd.t244 dvss 1.7295f
C6119 avdd.t240 dvss 1.7295f
C6120 avdd.t228 dvss 1.7295f
C6121 avdd.t230 dvss 1.7295f
C6122 avdd.t226 dvss 1.29713f
C6123 avdd.n1859 dvss 0.864751f
C6124 avdd.t224 dvss 1.29713f
C6125 avdd.t238 dvss 1.7295f
C6126 avdd.t236 dvss 1.7295f
C6127 avdd.t242 dvss 1.7295f
C6128 avdd.t234 dvss 1.7295f
C6129 avdd.t232 dvss 1.7295f
C6130 avdd.t220 dvss 1.7295f
C6131 avdd.t246 dvss 2.09379f
C6132 avdd.n1860 dvss 2.688f
C6133 avdd.n1861 dvss 0.279066f
C6134 avdd.n1862 dvss 0.480793f
C6135 avdd.n1863 dvss 0.949341f
C6136 avdd.n1864 dvss 0.890518f
C6137 avdd.n1865 dvss 0.323876f
C6138 avdd.n1866 dvss 1.20838f
C6139 avdd.n1867 dvss 1.02121f
C6140 avdd.n1868 dvss 0.95743f
C6141 avdd.n1869 dvss 1.59047f
C6142 avdd.n1870 dvss 0.954262f
C6143 avdd.n1871 dvss 0.556102f
C6144 avdd.n1872 dvss 0.138715f
C6145 avdd.n1873 dvss 3.7117f
C6146 avdd.t434 dvss 2.09379f
C6147 avdd.t433 dvss 1.7295f
C6148 avdd.t171 dvss 1.7295f
C6149 avdd.t559 dvss 1.7295f
C6150 avdd.t558 dvss 1.7295f
C6151 avdd.t40 dvss 1.7295f
C6152 avdd.t458 dvss 1.7295f
C6153 avdd.t459 dvss 1.7295f
C6154 avdd.t16 dvss 1.7295f
C6155 avdd.t471 dvss 1.7295f
C6156 avdd.t470 dvss 1.7295f
C6157 avdd.t73 dvss 1.7295f
C6158 avdd.t261 dvss 1.7295f
C6159 avdd.t260 dvss 1.7295f
C6160 avdd.t169 dvss 1.7295f
C6161 avdd.t591 dvss 1.7295f
C6162 avdd.t590 dvss 1.7295f
C6163 avdd.t157 dvss 1.7295f
C6164 avdd.t465 dvss 1.7295f
C6165 avdd.t464 dvss 1.7295f
C6166 avdd.t106 dvss 1.7295f
C6167 avdd.t426 dvss 1.7295f
C6168 avdd.t425 dvss 1.7295f
C6169 avdd.t38 dvss 1.7295f
C6170 avdd.t653 dvss 1.7295f
C6171 avdd.t654 dvss 1.7295f
C6172 avdd.t141 dvss 1.7295f
C6173 avdd.t595 dvss 1.7295f
C6174 avdd.t594 dvss 1.7295f
C6175 avdd.t67 dvss 1.7295f
C6176 avdd.t469 dvss 1.7295f
C6177 avdd.t468 dvss 1.7295f
C6178 avdd.t164 dvss 1.7295f
C6179 avdd.t561 dvss 1.7295f
C6180 avdd.t560 dvss 1.7295f
C6181 avdd.t118 dvss 1.7295f
C6182 avdd.t451 dvss 1.7295f
C6183 avdd.t452 dvss 1.7295f
C6184 avdd.t31 dvss 1.7295f
C6185 avdd.t526 dvss 1.7295f
C6186 avdd.t527 dvss 1.7295f
C6187 avdd.t99 dvss 1.7295f
C6188 avdd.t215 dvss 1.7295f
C6189 avdd.t214 dvss 1.7295f
C6190 avdd.t53 dvss 1.7295f
C6191 avdd.t430 dvss 1.7295f
C6192 avdd.t429 dvss 2.09379f
C6193 avdd.n1874 dvss 3.7117f
C6194 avdd.n1875 dvss 0.138971f
C6195 avdd.n1876 dvss 0.555412f
C6196 avdd.n1877 dvss 0.260284f
C6197 avdd.n1878 dvss 1.13707f
C6198 avdd.n1879 dvss 0.864789f
C6199 por_ana_0.comparator_0.vpp.n0 dvss 5.66344f
C6200 por_ana_0.comparator_0.vpp.n1 dvss 4.40814f
C6201 por_ana_0.comparator_0.vpp.n2 dvss 8.24237f
C6202 por_ana_0.comparator_0.vpp.n3 dvss 1.30683f
C6203 por_ana_0.comparator_0.vpp.n4 dvss 1.30683f
C6204 por_ana_0.comparator_0.vpp.t8 dvss 1.44245f
C6205 por_ana_0.comparator_0.vpp.t2 dvss 1.44245f
C6206 por_ana_0.comparator_0.vpp.t10 dvss 1.44245f
C6207 por_ana_0.comparator_0.vpp.t4 dvss 1.44245f
C6208 por_ana_0.comparator_0.vpp.t14 dvss 1.44245f
C6209 por_ana_0.comparator_0.vpp.t12 dvss 1.44245f
C6210 por_ana_0.comparator_0.vpp.t6 dvss 1.44245f
C6211 por_ana_0.comparator_0.vpp.t0 dvss 1.44245f
C6212 por_ana_0.comparator_0.vpp.t60 dvss 1.53356f
C6213 por_ana_0.comparator_0.vpp.t58 dvss 1.34009f
C6214 por_ana_0.comparator_0.vpp.t48 dvss 1.53356f
C6215 por_ana_0.comparator_0.vpp.t61 dvss 1.34009f
C6216 por_ana_0.comparator_0.vpp.t62 dvss 1.53356f
C6217 por_ana_0.comparator_0.vpp.t59 dvss 1.34009f
C6218 por_ana_0.comparator_0.vpp.t53 dvss 1.53356f
C6219 por_ana_0.comparator_0.vpp.t50 dvss 1.34009f
C6220 por_ana_0.comparator_0.vpp.t49 dvss 1.53356f
C6221 por_ana_0.comparator_0.vpp.t47 dvss 1.34009f
C6222 por_ana_0.comparator_0.vpp.t54 dvss 1.53356f
C6223 por_ana_0.comparator_0.vpp.t55 dvss 1.34009f
C6224 por_ana_0.comparator_0.vpp.t56 dvss 1.53356f
C6225 por_ana_0.comparator_0.vpp.t57 dvss 1.34009f
C6226 por_ana_0.comparator_0.vpp.t51 dvss 1.53356f
C6227 por_ana_0.comparator_0.vpp.t52 dvss 1.34009f
.ends

