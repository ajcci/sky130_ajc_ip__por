magic
tech sky130A
magscale 1 2
timestamp 1712973328
<< error_s >>
rect 39827 23173 39828 23227
rect 39887 23123 39888 23173
rect 39887 22853 39888 22937
<< pwell >>
rect -1182 40391 42901 40527
rect -1182 -559 -1046 40391
rect 42765 -559 42901 40391
rect -1182 -695 42901 -559
<< psubdiff >>
rect -1146 40457 -1086 40491
rect 42805 40457 42865 40491
rect -1146 40431 -1112 40457
rect -1146 -625 -1112 -599
rect 42831 40431 42865 40457
rect 42831 -625 42865 -599
rect -1146 -659 -1086 -625
rect 42805 -659 42865 -625
<< psubdiffcont >>
rect -1086 40457 42805 40491
rect -1146 -599 -1112 40431
rect 42831 -599 42865 40431
rect -1086 -659 42805 -625
<< locali >>
rect -1146 40457 -1086 40491
rect 42805 40457 42865 40491
rect -1146 40431 -1112 40457
rect 42831 40431 42865 40457
rect 40265 27929 40313 27977
rect -1146 -625 -1112 -599
rect 42831 -625 42865 -599
rect -1146 -659 -1086 -625
rect 42805 -659 42865 -625
<< viali >>
rect -1086 40457 42805 40491
rect -1146 -556 -1112 40404
rect 27965 38035 29655 38069
rect 27965 37449 29655 37483
rect 42831 -567 42865 40393
rect -1086 -659 42805 -625
<< metal1 >>
rect 41177 40601 41325 40612
rect 41177 40531 41188 40601
rect -1186 40491 41188 40531
rect 41314 40531 41325 40601
rect 41314 40491 42905 40531
rect -1186 40457 -1086 40491
rect 42805 40457 42905 40491
rect -1186 40404 42905 40457
rect -1186 -556 -1146 40404
rect -1112 40393 42905 40404
rect -1112 40391 42831 40393
rect -1112 -556 -1046 40391
rect 27857 38069 29763 38081
rect 27857 38066 27965 38069
rect 27851 38014 27857 38066
rect 27909 38035 27965 38066
rect 29655 38035 29763 38069
rect 27909 38023 29763 38035
rect 27909 38014 27915 38023
rect 27857 37495 27915 38014
rect 28450 37791 28514 37797
rect 28133 37777 28197 37783
rect 28133 37725 28139 37777
rect 28191 37725 28197 37777
rect 28450 37739 28456 37791
rect 28508 37739 28514 37791
rect 28450 37733 28514 37739
rect 28771 37793 28835 37799
rect 28771 37741 28777 37793
rect 28829 37741 28835 37793
rect 28771 37735 28835 37741
rect 29087 37793 29151 37799
rect 29087 37741 29093 37793
rect 29145 37741 29151 37793
rect 29087 37735 29151 37741
rect 29407 37794 29471 37800
rect 29407 37742 29413 37794
rect 29465 37742 29471 37794
rect 29407 37736 29471 37742
rect 28133 37719 28197 37725
rect 27997 37627 28043 37659
rect 28313 37627 28359 37659
rect 28629 37627 28675 37659
rect 28945 37627 28991 37659
rect 29261 37627 29307 37659
rect 29577 37627 29623 37660
rect 27997 37581 28053 37627
rect 28145 37581 29475 37627
rect 29567 37581 29623 37627
rect 28053 37495 28145 37581
rect 29705 37495 29763 38023
rect 27857 37483 29763 37495
rect 27857 37449 27965 37483
rect 29655 37449 29763 37483
rect 27857 37437 29763 37449
rect 42223 27573 42301 27619
rect 42255 27563 42301 27573
rect 42067 27462 42131 27468
rect 42067 27410 42073 27462
rect 42125 27410 42131 27462
rect 42067 27404 42131 27410
rect 42255 27303 42301 27471
rect 42223 27257 42301 27303
rect 42134 27146 42198 27152
rect 42134 27094 42140 27146
rect 42192 27094 42198 27146
rect 42134 27088 42198 27094
rect 42255 26987 42301 27257
rect 42223 26941 42301 26987
rect 42024 26821 42088 26827
rect 42024 26769 42030 26821
rect 42082 26769 42088 26821
rect 42024 26763 42088 26769
rect 42255 26671 42301 26941
rect 42223 26625 42301 26671
rect 42084 26514 42158 26525
rect 42084 26462 42095 26514
rect 42147 26462 42158 26514
rect 42084 26451 42158 26462
rect 42255 26355 42301 26625
rect 42223 26309 42301 26355
rect 42104 26196 42178 26207
rect 42104 26144 42115 26196
rect 42167 26144 42178 26196
rect 42104 26133 42178 26144
rect 42255 26039 42301 26309
rect 42223 25993 42301 26039
rect 42096 25882 42170 25893
rect 42096 25830 42107 25882
rect 42159 25830 42170 25882
rect 42096 25819 42170 25830
rect 42255 25723 42301 25993
rect 42223 25677 42301 25723
rect 42134 25563 42198 25569
rect 42134 25511 42140 25563
rect 42192 25511 42198 25563
rect 42134 25505 42198 25511
rect 42255 25407 42301 25677
rect 42223 25388 42301 25407
rect 42765 25388 42831 40391
rect 42223 25361 42831 25388
rect 42255 25281 42831 25361
rect 42036 25247 42100 25253
rect 42036 25195 42042 25247
rect 42094 25195 42100 25247
rect 42036 25189 42100 25195
rect 42255 25193 42301 25281
rect 42255 25091 42301 25119
rect 42223 25045 42301 25091
rect 4280 348 4344 354
rect 4280 296 4286 348
rect 4338 296 4344 348
rect 4280 290 4344 296
rect 4136 179 4182 211
rect 4452 186 4498 211
rect 4452 180 4520 186
rect 4452 179 4462 180
rect 4136 133 4192 179
rect 4284 133 4350 179
rect 4442 133 4462 179
rect 4456 128 4462 133
rect 4514 128 4520 180
rect 4456 122 4520 128
rect -1186 -559 -1046 -556
rect 42765 -559 42831 25281
rect -1186 -567 42831 -559
rect 42865 -567 42905 40393
rect -1186 -625 42905 -567
rect -1186 -659 -1086 -625
rect 42805 -659 42905 -625
rect -1186 -699 42905 -659
<< via1 >>
rect 41188 40491 41314 40601
rect 41188 40475 41314 40491
rect 27857 38014 27909 38066
rect 28139 37725 28191 37777
rect 28456 37739 28508 37791
rect 28777 37741 28829 37793
rect 29093 37741 29145 37793
rect 29413 37742 29465 37794
rect 42073 27410 42125 27462
rect 42140 27094 42192 27146
rect 42030 26769 42082 26821
rect 42095 26462 42147 26514
rect 42115 26144 42167 26196
rect 42107 25830 42159 25882
rect 42140 25511 42192 25563
rect 42042 25195 42094 25247
rect 4286 296 4338 348
rect 4462 128 4514 180
<< metal2 >>
rect 1111 40272 1507 40292
rect 1111 39982 1131 40272
rect 1471 39982 1507 40272
rect 1111 39265 1507 39982
rect 1577 39865 1962 39896
rect 1577 39606 1599 39865
rect 1934 39606 1962 39865
rect 1577 39251 1962 39606
rect 10947 37781 11011 41282
rect 10938 37717 10947 37781
rect 11011 37717 11020 37781
rect 10947 32696 11011 37717
rect 10947 32632 11144 32696
rect 11080 32421 11144 32632
rect 11863 26526 11915 41282
rect 12176 38006 12236 41282
rect 12176 32368 12236 37946
rect 12176 32312 12178 32368
rect 12234 32312 12236 32368
rect 12176 32310 12236 32312
rect 12178 32303 12234 32310
rect 14069 23632 14078 23696
rect 14142 23632 14151 23696
rect 14947 23692 15011 41282
rect 24466 41068 24594 41077
rect 14947 23636 14951 23692
rect 15007 23636 15011 23692
rect 14947 23632 15011 23636
rect 19684 34398 19744 34407
rect 14951 23627 15007 23632
rect 4280 7138 4354 7147
rect 4280 7082 4289 7138
rect 4345 7082 4354 7138
rect 4280 7077 4354 7082
rect 10 -707 396 1690
rect 493 -110 893 1899
rect 4287 354 4347 7077
rect 15261 4203 15317 4210
rect 15259 4201 15319 4203
rect 15259 4145 15261 4201
rect 15317 4145 15319 4201
rect 15259 3495 15319 4145
rect 15157 3435 15319 3495
rect 18496 3531 18556 3540
rect 19684 3529 19744 34338
rect 24466 30961 24594 40940
rect 24666 40744 24794 40753
rect 24666 30932 24794 40616
rect 24320 30877 24380 30886
rect 26956 30851 27008 41282
rect 27302 39425 27358 41282
rect 19930 28201 19990 28210
rect 19921 28141 19930 28197
rect 19990 28141 19999 28197
rect 19930 4203 19990 28141
rect 21332 27822 21388 27829
rect 21330 27820 21390 27822
rect 21330 27764 21332 27820
rect 21388 27764 21390 27820
rect 21330 23716 21390 27764
rect 23126 27660 23182 27667
rect 23124 27658 23184 27660
rect 23124 27602 23126 27658
rect 23182 27602 23184 27658
rect 21508 26814 21564 26821
rect 21506 26812 21566 26814
rect 21506 26756 21508 26812
rect 21564 26756 21566 26812
rect 21506 22328 21566 26756
rect 23124 23396 23184 27602
rect 23637 26947 23693 26954
rect 23635 26945 23695 26947
rect 23635 26889 23637 26945
rect 23693 26889 23695 26945
rect 23635 23875 23695 26889
rect 24320 26680 24380 30817
rect 26883 30799 27008 30851
rect 27235 39369 27358 39425
rect 26802 30024 26858 30033
rect 26802 29959 26858 29968
rect 26785 28398 26845 28407
rect 26785 28329 26845 28338
rect 26787 27893 26843 28329
rect 26787 27837 26932 27893
rect 25396 27508 25452 27515
rect 24320 26624 24322 26680
rect 24378 26624 24380 26680
rect 24320 26622 24380 26624
rect 25394 27506 25454 27508
rect 25394 27450 25396 27506
rect 25452 27450 25454 27506
rect 24322 26615 24378 26622
rect 23448 23815 23695 23875
rect 23124 23336 23498 23396
rect 21337 22268 21566 22328
rect 21337 22054 21397 22268
rect 23438 22074 23498 23336
rect 25394 22642 25454 27450
rect 25556 27228 25612 27235
rect 25554 27226 25614 27228
rect 25554 27170 25556 27226
rect 25612 27170 25614 27226
rect 25554 23786 25614 27170
rect 27235 27158 27291 39369
rect 27692 34401 27752 41282
rect 27991 40491 28051 40500
rect 27991 40422 28051 40431
rect 27995 38618 28047 40422
rect 27857 38566 28047 38618
rect 28779 38586 28835 38593
rect 28777 38584 28837 38586
rect 27857 38066 27909 38566
rect 27857 38008 27909 38014
rect 28777 38528 28779 38584
rect 28835 38528 28837 38584
rect 28456 38006 28512 38013
rect 28454 38004 28514 38006
rect 28454 37948 28456 38004
rect 28512 37948 28514 38004
rect 28454 37797 28514 37948
rect 28777 37799 28837 38528
rect 29097 38432 29153 38439
rect 29095 38430 29155 38432
rect 29095 38374 29097 38430
rect 29153 38374 29155 38430
rect 29095 37799 29155 38374
rect 29410 38274 29466 38281
rect 29408 38272 29468 38274
rect 29408 38216 29410 38272
rect 29466 38216 29468 38272
rect 29408 37800 29468 38216
rect 28450 37791 28514 37797
rect 28131 37783 28187 37786
rect 28131 37777 28197 37783
rect 28191 37725 28197 37777
rect 28450 37739 28456 37791
rect 28508 37739 28514 37791
rect 28450 37733 28514 37739
rect 28771 37793 28837 37799
rect 28771 37741 28777 37793
rect 28829 37741 28837 37793
rect 28771 37736 28837 37741
rect 29087 37793 29155 37799
rect 29087 37741 29093 37793
rect 29145 37741 29155 37793
rect 29087 37739 29155 37741
rect 29407 37794 29471 37800
rect 29407 37742 29413 37794
rect 29465 37742 29471 37794
rect 28771 37735 28835 37736
rect 29087 37735 29151 37739
rect 29407 37736 29471 37742
rect 28187 37721 28197 37725
rect 28131 37719 28197 37721
rect 28131 37712 28187 37719
rect 27685 34396 27759 34401
rect 27685 34340 27694 34396
rect 27750 34340 27759 34396
rect 27685 34331 27759 34340
rect 29742 30313 29802 41282
rect 32348 38608 32376 41282
rect 32992 38615 33020 41282
rect 38788 38621 38816 41282
rect 41177 40603 41325 40612
rect 41177 40473 41186 40603
rect 41316 40473 41325 40603
rect 41177 40464 41325 40473
rect 32323 38586 32401 38595
rect 32323 38526 32332 38586
rect 32392 38526 32401 38586
rect 32323 38517 32401 38526
rect 32967 38432 33045 38441
rect 32967 38372 32976 38432
rect 33036 38372 33045 38432
rect 32967 38363 33045 38372
rect 38763 38274 38841 38283
rect 38763 38214 38772 38274
rect 38832 38214 38841 38274
rect 38763 38205 38841 38214
rect 31111 38144 31167 38151
rect 38119 38144 38197 38153
rect 31109 38142 31169 38144
rect 31109 38086 31111 38142
rect 31167 38086 31169 38142
rect 30945 37995 31001 38002
rect 30943 37993 31003 37995
rect 30943 37937 30945 37993
rect 31001 37937 31003 37993
rect 30810 37852 30866 37859
rect 30808 37850 30868 37852
rect 30808 37794 30810 37850
rect 30866 37794 30868 37850
rect 30657 37703 30713 37710
rect 30655 37701 30715 37703
rect 30655 37645 30657 37701
rect 30713 37645 30715 37701
rect 30112 37569 30168 37576
rect 30110 37567 30170 37569
rect 30110 37511 30112 37567
rect 30168 37511 30170 37567
rect 29963 35081 30019 35088
rect 27842 30026 27902 30035
rect 27842 28044 27902 29966
rect 29742 28396 29802 30253
rect 29742 28340 29744 28396
rect 29800 28340 29802 28396
rect 29742 28338 29802 28340
rect 29961 35079 30021 35081
rect 29961 35023 29963 35079
rect 30019 35023 30021 35079
rect 29744 28331 29800 28338
rect 27842 27988 27844 28044
rect 27900 27988 27902 28044
rect 27842 27986 27902 27988
rect 27844 27979 27900 27986
rect 27504 27368 27560 27375
rect 27502 27366 27562 27368
rect 27502 27310 27504 27366
rect 27560 27310 27562 27366
rect 27235 27102 27376 27158
rect 25394 22582 25614 22642
rect 25554 22032 25614 22582
rect 27502 22332 27562 27310
rect 27676 27088 27732 27095
rect 27674 27086 27734 27088
rect 27674 27030 27676 27086
rect 27732 27030 27734 27086
rect 27674 23750 27734 27030
rect 29961 25717 30021 35023
rect 29961 25648 30021 25657
rect 29783 23848 29839 23857
rect 29783 23783 29839 23792
rect 29776 22335 29832 22342
rect 30110 22335 30170 37511
rect 30502 37443 30558 37450
rect 30500 37441 30560 37443
rect 30500 37385 30502 37441
rect 30558 37385 30560 37441
rect 30266 37312 30322 37319
rect 30264 37310 30324 37312
rect 30264 37254 30266 37310
rect 30322 37254 30324 37310
rect 30264 23850 30324 37254
rect 30383 37187 30439 37194
rect 30264 23781 30324 23790
rect 30381 37185 30441 37187
rect 30381 37129 30383 37185
rect 30439 37129 30441 37185
rect 29774 22333 29834 22335
rect 27502 22272 27726 22332
rect 27666 22088 27726 22272
rect 29774 22277 29776 22333
rect 29832 22277 29834 22333
rect 29774 22108 29834 22277
rect 30110 22266 30170 22275
rect 30381 22306 30441 37129
rect 30500 26524 30560 37385
rect 30500 26455 30560 26464
rect 30655 26370 30715 37645
rect 30655 26301 30715 26310
rect 30808 26202 30868 37794
rect 30808 26133 30868 26142
rect 30943 26029 31003 37937
rect 30943 25960 31003 25969
rect 31109 25870 31169 38086
rect 38119 38084 38128 38144
rect 38188 38084 38197 38144
rect 38119 38075 38197 38084
rect 37475 37995 37553 38004
rect 37475 37935 37484 37995
rect 37544 37935 37553 37995
rect 37475 37926 37553 37935
rect 36831 37792 36840 37852
rect 36900 37792 36909 37852
rect 36187 37703 36265 37712
rect 36187 37643 36196 37703
rect 36256 37643 36265 37703
rect 36187 37634 36265 37643
rect 35543 37569 35621 37578
rect 35543 37509 35552 37569
rect 35612 37509 35621 37569
rect 35543 37500 35621 37509
rect 34908 37443 34968 37452
rect 34908 37374 34968 37383
rect 34255 37312 34333 37321
rect 34255 37252 34264 37312
rect 34324 37252 34333 37312
rect 34255 37243 34333 37252
rect 33611 37187 33689 37196
rect 33611 37127 33620 37187
rect 33680 37127 33689 37187
rect 33611 37118 33689 37127
rect 42249 33716 42316 33725
rect 42249 33660 42258 33716
rect 42314 33660 42316 33716
rect 42249 33655 42316 33660
rect 40462 33036 40536 33045
rect 40462 32980 40471 33036
rect 40527 32980 40536 33036
rect 40462 32975 40536 32980
rect 40469 32578 40529 32975
rect 40377 32518 40529 32578
rect 40377 32187 40437 32518
rect 40767 32358 40823 32365
rect 40765 32356 40825 32358
rect 40765 32300 40767 32356
rect 40823 32300 40825 32356
rect 40377 32127 40495 32187
rect 40293 30996 40367 31005
rect 40293 30940 40302 30996
rect 40358 30940 40367 30996
rect 40293 30935 40367 30940
rect 40300 28201 40360 30935
rect 40300 28132 40360 28141
rect 34908 27822 34968 27831
rect 34908 27753 34968 27762
rect 34255 27600 34264 27660
rect 34324 27600 34333 27660
rect 34924 27586 34952 27753
rect 37208 27508 37268 27517
rect 37208 27439 37268 27448
rect 37224 27368 37252 27439
rect 37484 27368 37544 27377
rect 37484 27299 37544 27308
rect 37500 27224 37528 27299
rect 38119 27168 38128 27228
rect 38188 27168 38197 27228
rect 38763 27088 38841 27097
rect 38763 27028 38772 27088
rect 38832 27028 38841 27088
rect 38763 27019 38841 27028
rect 33636 25882 33664 26991
rect 35568 26540 35596 27011
rect 35552 26531 35612 26540
rect 33854 26524 33910 26531
rect 33852 26522 33912 26524
rect 33852 26466 33854 26522
rect 33910 26466 33912 26522
rect 31897 25870 31953 25877
rect 33620 25873 33680 25882
rect 31109 25801 31169 25810
rect 31895 25868 31955 25870
rect 31895 25812 31897 25868
rect 31953 25812 31955 25868
rect 31895 23786 31955 25812
rect 33620 25804 33680 25813
rect 31892 22306 31948 22313
rect 30381 22237 30441 22246
rect 31890 22304 31950 22306
rect 31890 22248 31892 22304
rect 31948 22248 31950 22304
rect 31890 22097 31950 22248
rect 33852 22296 33912 26466
rect 35552 26462 35612 26471
rect 35943 26370 35999 26377
rect 35941 26368 36001 26370
rect 35941 26312 35943 26368
rect 35999 26312 36001 26368
rect 34007 26202 34063 26209
rect 34005 26200 34065 26202
rect 34005 26144 34007 26200
rect 34063 26144 34065 26200
rect 34005 23812 34065 26144
rect 35941 22315 36001 26312
rect 36212 26190 36240 26995
rect 39432 26956 39460 27250
rect 39416 26947 39476 26956
rect 39416 26878 39476 26887
rect 40076 26823 40104 27022
rect 40060 26814 40120 26823
rect 40060 26745 40120 26754
rect 40435 26682 40495 32127
rect 40765 28046 40825 32300
rect 41924 31676 41998 31685
rect 41924 31620 41933 31676
rect 41989 31620 41998 31676
rect 41924 31615 41998 31620
rect 40765 27977 40825 27986
rect 41931 26817 41991 31615
rect 42064 30316 42138 30325
rect 42064 30260 42073 30316
rect 42129 30260 42138 30316
rect 42064 30255 42138 30260
rect 42071 27468 42131 30255
rect 42067 27462 42131 27468
rect 42067 27410 42073 27462
rect 42125 27410 42131 27462
rect 42067 27404 42131 27410
rect 42071 27396 42131 27404
rect 42256 27154 42316 33655
rect 42124 27146 42316 27154
rect 42124 27094 42140 27146
rect 42192 27094 42316 27146
rect 42134 27088 42198 27094
rect 42024 26821 42088 26827
rect 42024 26817 42030 26821
rect 41931 26769 42030 26817
rect 42082 26817 42088 26821
rect 42082 26769 42091 26817
rect 41931 26757 42091 26769
rect 40435 26613 40495 26622
rect 42084 26516 42158 26525
rect 42084 26460 42093 26516
rect 42149 26460 42158 26516
rect 42084 26451 42158 26460
rect 42104 26198 42178 26207
rect 36196 26181 36256 26190
rect 42104 26142 42113 26198
rect 42169 26142 42178 26198
rect 42104 26133 42178 26142
rect 36196 26112 36256 26121
rect 36128 26027 36188 26029
rect 36121 25971 36130 26027
rect 36186 25971 36195 26027
rect 36128 23792 36188 25971
rect 42096 25884 42170 25893
rect 42096 25828 42105 25884
rect 42161 25828 42170 25884
rect 42096 25819 42170 25828
rect 38020 25717 38076 25724
rect 38018 25715 38078 25717
rect 38018 25659 38020 25715
rect 38076 25659 38078 25715
rect 38018 23197 38078 25659
rect 42151 25569 42211 25577
rect 42134 25563 42211 25569
rect 42134 25511 42140 25563
rect 42192 25511 42211 25563
rect 42134 25505 42211 25511
rect 42036 25252 42100 25253
rect 42036 25247 42105 25252
rect 42036 25195 42042 25247
rect 42094 25195 42105 25247
rect 42036 25189 42105 25195
rect 38213 23730 38222 23794
rect 38286 23730 38295 23794
rect 42041 23790 42105 25189
rect 42036 23734 42045 23790
rect 42101 23734 42110 23790
rect 42041 23730 42105 23734
rect 42151 23200 42211 25505
rect 38009 23137 38018 23197
rect 38078 23137 38087 23197
rect 42144 23195 42218 23200
rect 42144 23139 42153 23195
rect 42209 23139 42218 23195
rect 33852 22236 34060 22296
rect 35941 22255 36175 22315
rect 34000 22055 34060 22236
rect 36115 22040 36175 22255
rect 38018 22281 38078 23137
rect 42144 23130 42218 23139
rect 38018 22221 38276 22281
rect 38216 22103 38276 22221
rect 19930 4134 19990 4143
rect 19677 3473 19686 3529
rect 19742 3473 19751 3529
rect 19684 3471 19744 3473
rect 18496 3462 18556 3471
rect 4280 348 4347 354
rect 4280 296 4286 348
rect 4338 296 4347 348
rect 4280 290 4347 296
rect 493 -519 893 -510
rect 10 -1039 28 -707
rect 383 -1039 396 -707
rect 10 -1056 396 -1039
rect 4287 -1987 4347 290
rect 4456 180 4520 186
rect 4456 128 4462 180
rect 4514 128 4520 180
rect 4456 -1190 4520 128
rect 4456 -1263 4520 -1254
<< via2 >>
rect 1131 39982 1471 40272
rect 1599 39606 1934 39865
rect 10947 37717 11011 37781
rect 12176 37946 12236 38006
rect 12178 32312 12234 32368
rect 14078 23632 14142 23696
rect 24466 40940 24594 41068
rect 14951 23636 15007 23692
rect 19684 34338 19744 34398
rect 4289 7082 4345 7138
rect 15261 4145 15317 4201
rect 18496 3471 18556 3531
rect 24666 40616 24794 40744
rect 24320 30817 24380 30877
rect 19930 28141 19990 28201
rect 21332 27764 21388 27820
rect 23126 27602 23182 27658
rect 21508 26756 21564 26812
rect 23637 26889 23693 26945
rect 26802 29968 26858 30024
rect 26785 28338 26845 28398
rect 24322 26624 24378 26680
rect 25396 27450 25452 27506
rect 25556 27170 25612 27226
rect 27991 40431 28051 40491
rect 28779 38528 28835 38584
rect 28456 37948 28512 38004
rect 29097 38374 29153 38430
rect 29410 38216 29466 38272
rect 28131 37725 28139 37777
rect 28139 37725 28187 37777
rect 28131 37721 28187 37725
rect 27694 34340 27750 34396
rect 41186 40601 41316 40603
rect 41186 40475 41188 40601
rect 41188 40475 41314 40601
rect 41314 40475 41316 40601
rect 41186 40473 41316 40475
rect 32332 38526 32392 38586
rect 32976 38372 33036 38432
rect 38772 38214 38832 38274
rect 31111 38086 31167 38142
rect 30945 37937 31001 37993
rect 30810 37794 30866 37850
rect 30657 37645 30713 37701
rect 30112 37511 30168 37567
rect 29742 30253 29802 30313
rect 27842 29966 27902 30026
rect 29744 28340 29800 28396
rect 29963 35023 30019 35079
rect 27844 27988 27900 28044
rect 27504 27310 27560 27366
rect 27676 27030 27732 27086
rect 29961 25657 30021 25717
rect 29783 23792 29839 23848
rect 30502 37385 30558 37441
rect 30266 37254 30322 37310
rect 30264 23790 30324 23850
rect 30383 37129 30439 37185
rect 29776 22277 29832 22333
rect 30110 22275 30170 22335
rect 30500 26464 30560 26524
rect 30655 26310 30715 26370
rect 30808 26142 30868 26202
rect 30943 25969 31003 26029
rect 38128 38084 38188 38144
rect 37484 37935 37544 37995
rect 36840 37792 36900 37852
rect 36196 37643 36256 37703
rect 35552 37509 35612 37569
rect 34908 37383 34968 37443
rect 34264 37252 34324 37312
rect 33620 37127 33680 37187
rect 42258 33660 42314 33716
rect 40471 32980 40527 33036
rect 40767 32300 40823 32356
rect 40302 30940 40358 30996
rect 40300 28141 40360 28201
rect 34908 27762 34968 27822
rect 34264 27600 34324 27660
rect 37208 27448 37268 27508
rect 37484 27308 37544 27368
rect 38128 27168 38188 27228
rect 38772 27028 38832 27088
rect 33854 26466 33910 26522
rect 31109 25810 31169 25870
rect 31897 25812 31953 25868
rect 33620 25813 33680 25873
rect 30381 22246 30441 22306
rect 31892 22248 31948 22304
rect 35552 26471 35612 26531
rect 35943 26312 35999 26368
rect 34007 26144 34063 26200
rect 39416 26887 39476 26947
rect 40060 26754 40120 26814
rect 41933 31620 41989 31676
rect 40765 27986 40825 28046
rect 42073 30260 42129 30316
rect 40435 26622 40495 26682
rect 42093 26514 42149 26516
rect 42093 26462 42095 26514
rect 42095 26462 42147 26514
rect 42147 26462 42149 26514
rect 42093 26460 42149 26462
rect 36196 26121 36256 26181
rect 42113 26196 42169 26198
rect 42113 26144 42115 26196
rect 42115 26144 42167 26196
rect 42167 26144 42169 26196
rect 42113 26142 42169 26144
rect 36130 25971 36186 26027
rect 42105 25882 42161 25884
rect 42105 25830 42107 25882
rect 42107 25830 42159 25882
rect 42159 25830 42161 25882
rect 42105 25828 42161 25830
rect 38020 25659 38076 25715
rect 38222 23730 38286 23794
rect 42045 23734 42101 23790
rect 38018 23137 38078 23197
rect 42153 23139 42209 23195
rect 19930 4143 19990 4203
rect 19686 3473 19742 3529
rect 493 -510 893 -110
rect 28 -1039 383 -707
rect 4456 -1254 4520 -1190
<< metal3 >>
rect -1604 41276 43293 41282
rect -1604 40888 -1598 41276
rect -1210 41227 42899 41276
rect -1210 41068 34593 41227
rect -1210 40940 24466 41068
rect 24594 40940 34593 41068
rect -1210 40909 34593 40940
rect 34911 40909 42899 41227
rect -1210 40888 42899 40909
rect 43287 40888 43293 41276
rect -1604 40882 43293 40888
rect -1604 40816 43293 40822
rect -1604 40428 -1138 40816
rect -750 40779 42439 40816
rect -750 40744 35253 40779
rect -750 40616 24666 40744
rect 24794 40616 35253 40744
rect -750 40491 35253 40616
rect -750 40431 27991 40491
rect 28051 40461 35253 40491
rect 35571 40603 42439 40779
rect 35571 40473 41186 40603
rect 41316 40473 42439 40603
rect 35571 40461 42439 40473
rect 28051 40431 42439 40461
rect -750 40428 42439 40431
rect 42827 40428 43293 40816
rect -1604 40422 43293 40428
rect -1604 40356 43293 40362
rect -1604 39968 -678 40356
rect -290 40272 41979 40356
rect -290 39982 1131 40272
rect 1471 39982 41979 40272
rect -290 39968 41979 39982
rect 42367 39968 43293 40356
rect -1604 39962 43293 39968
rect -1604 39896 43293 39902
rect -1604 39508 -218 39896
rect 170 39865 41519 39896
rect 170 39606 1599 39865
rect 1934 39606 41519 39865
rect 170 39508 41519 39606
rect 41907 39508 43293 39896
rect -1604 39502 43293 39508
rect 947 39492 1357 39502
rect 28774 38586 28840 38589
rect 32327 38586 32397 38591
rect 28774 38584 32332 38586
rect 28774 38528 28779 38584
rect 28835 38528 32332 38584
rect 28774 38526 32332 38528
rect 32392 38526 32397 38586
rect 28774 38523 28840 38526
rect 32327 38521 32397 38526
rect 29092 38432 29158 38435
rect 32971 38432 33041 38437
rect 29092 38430 32976 38432
rect 29092 38374 29097 38430
rect 29153 38374 32976 38430
rect 29092 38372 32976 38374
rect 33036 38372 33041 38432
rect 29092 38369 29158 38372
rect 32971 38367 33041 38372
rect 29405 38274 29471 38277
rect 38767 38274 38837 38279
rect 29405 38272 38772 38274
rect 29405 38216 29410 38272
rect 29466 38216 38772 38272
rect 29405 38214 38772 38216
rect 38832 38214 38837 38274
rect 29405 38211 29471 38214
rect 38767 38209 38837 38214
rect 31106 38144 31172 38147
rect 38123 38144 38193 38149
rect 31106 38142 38128 38144
rect 31106 38086 31111 38142
rect 31167 38086 38128 38142
rect 31106 38084 38128 38086
rect 38188 38084 38193 38144
rect 31106 38081 31172 38084
rect 38123 38079 38193 38084
rect 12171 38006 12241 38011
rect 28451 38006 28517 38009
rect 12171 37946 12176 38006
rect 12236 38004 28517 38006
rect 12236 37948 28456 38004
rect 28512 37948 28517 38004
rect 12236 37946 28517 37948
rect 12171 37941 12241 37946
rect 28451 37943 28517 37946
rect 30940 37995 31006 37998
rect 37479 37995 37549 38000
rect 30940 37993 37484 37995
rect 30940 37937 30945 37993
rect 31001 37937 37484 37993
rect 30940 37935 37484 37937
rect 37544 37935 37549 37995
rect 30940 37932 31006 37935
rect 37479 37930 37549 37935
rect 30805 37852 30871 37855
rect 36835 37852 36905 37857
rect 30805 37850 36840 37852
rect 30805 37794 30810 37850
rect 30866 37794 36840 37850
rect 30805 37792 36840 37794
rect 36900 37792 36905 37852
rect 30805 37789 30871 37792
rect 36835 37787 36905 37792
rect 10942 37781 11016 37786
rect 28126 37781 28192 37782
rect 10942 37717 10947 37781
rect 11011 37777 28192 37781
rect 11011 37721 28131 37777
rect 28187 37721 28192 37777
rect 11011 37717 28192 37721
rect 10942 37712 11016 37717
rect 28126 37716 28192 37717
rect 30652 37703 30718 37706
rect 36191 37703 36261 37708
rect 30652 37701 36196 37703
rect 30652 37645 30657 37701
rect 30713 37645 36196 37701
rect 30652 37643 36196 37645
rect 36256 37643 36261 37703
rect 30652 37640 30718 37643
rect 36191 37638 36261 37643
rect 30107 37569 30173 37572
rect 35547 37569 35617 37574
rect 30107 37567 35552 37569
rect 30107 37511 30112 37567
rect 30168 37511 35552 37567
rect 30107 37509 35552 37511
rect 35612 37509 35617 37569
rect 30107 37506 30173 37509
rect 35547 37504 35617 37509
rect 30497 37443 30563 37446
rect 34903 37443 34973 37448
rect 30497 37441 34908 37443
rect 30497 37385 30502 37441
rect 30558 37385 34908 37441
rect 30497 37383 34908 37385
rect 34968 37383 34973 37443
rect 30497 37380 30563 37383
rect 34903 37378 34973 37383
rect 30261 37312 30327 37315
rect 34259 37312 34329 37317
rect 30261 37310 34264 37312
rect 30261 37254 30266 37310
rect 30322 37254 34264 37310
rect 30261 37252 34264 37254
rect 34324 37252 34329 37312
rect 30261 37249 30327 37252
rect 34259 37247 34329 37252
rect 30378 37187 30444 37190
rect 33615 37187 33685 37192
rect 30378 37185 33620 37187
rect 30378 37129 30383 37185
rect 30439 37129 33620 37185
rect 30378 37127 33620 37129
rect 33680 37127 33685 37187
rect 30378 37124 30444 37127
rect 33615 37122 33685 37127
rect 29958 35081 30024 35084
rect 29958 35079 30384 35081
rect 29958 35023 29963 35079
rect 30019 35075 30384 35079
rect 30019 35023 31282 35075
rect 29958 35021 31282 35023
rect 29958 35018 30024 35021
rect 19679 34398 19749 34403
rect 27689 34398 27755 34401
rect 19679 34338 19684 34398
rect 19744 34396 30674 34398
rect 19744 34340 27694 34396
rect 27750 34340 30674 34396
rect 19744 34338 30674 34340
rect 40676 34338 43293 34398
rect 19679 34333 19749 34338
rect 27689 34335 27755 34338
rect 42253 33718 42319 33721
rect 40679 33716 43293 33718
rect 40679 33660 42258 33716
rect 42314 33660 43293 33716
rect 40679 33658 43293 33660
rect 42253 33655 42319 33658
rect 40466 33036 40532 33041
rect 40466 32980 40471 33036
rect 40527 32980 40532 33036
rect 40466 32975 40532 32980
rect 12173 32370 12239 32373
rect 11246 32368 12239 32370
rect 11246 32312 12178 32368
rect 12234 32312 12239 32368
rect 40762 32358 40828 32361
rect 11246 32310 12239 32312
rect 12173 32307 12239 32310
rect 40633 32356 43293 32358
rect 40633 32300 40767 32356
rect 40823 32300 43293 32356
rect 40633 32298 43293 32300
rect 40762 32295 40828 32298
rect 41928 31678 41994 31681
rect 40674 31676 43293 31678
rect 40674 31620 41933 31676
rect 41989 31620 43293 31676
rect 40674 31618 43293 31620
rect 41928 31615 41994 31618
rect 40297 30996 40363 31001
rect 40297 30940 40302 30996
rect 40358 30940 40363 30996
rect 40297 30935 40363 30940
rect 24315 30877 24385 30882
rect 24315 30817 24320 30877
rect 24380 30817 25001 30877
rect 24315 30812 24385 30817
rect 42068 30318 42134 30321
rect 29737 30313 29807 30318
rect 40657 30316 43293 30318
rect 29737 30253 29742 30313
rect 29802 30253 30759 30313
rect 40657 30260 42073 30316
rect 42129 30260 43293 30316
rect 40657 30258 43293 30260
rect 42068 30255 42134 30258
rect 29737 30248 29807 30253
rect 26797 30026 26863 30029
rect 27837 30026 27907 30031
rect 26797 30024 27842 30026
rect 26797 29968 26802 30024
rect 26858 29968 27842 30024
rect 26797 29966 27842 29968
rect 27902 29966 27907 30026
rect 26797 29963 26863 29966
rect 27837 29961 27907 29966
rect 26780 28398 26850 28403
rect 29739 28398 29805 28401
rect 26780 28338 26785 28398
rect 26845 28396 29805 28398
rect 26845 28340 29744 28396
rect 29800 28340 29805 28396
rect 26845 28338 29805 28340
rect 26780 28333 26850 28338
rect 29739 28335 29805 28338
rect 19925 28201 19995 28206
rect 40295 28201 40365 28206
rect 19925 28141 19930 28201
rect 19990 28141 40300 28201
rect 40360 28141 40365 28201
rect 19925 28136 19995 28141
rect 40295 28136 40365 28141
rect 27839 28046 27905 28049
rect 40760 28046 40830 28051
rect 27839 28044 40765 28046
rect 27839 27988 27844 28044
rect 27900 27988 40765 28044
rect 27839 27986 40765 27988
rect 40825 27986 40830 28046
rect 27839 27983 27905 27986
rect 40760 27981 40830 27986
rect 21327 27822 21393 27825
rect 34903 27822 34973 27827
rect 21327 27820 34908 27822
rect 21327 27764 21332 27820
rect 21388 27764 34908 27820
rect 21327 27762 34908 27764
rect 34968 27762 34973 27822
rect 21327 27759 21393 27762
rect 34903 27757 34973 27762
rect 23121 27660 23187 27663
rect 34259 27660 34329 27665
rect 23121 27658 34264 27660
rect 23121 27602 23126 27658
rect 23182 27602 34264 27658
rect 23121 27600 34264 27602
rect 34324 27600 34329 27660
rect 23121 27597 23187 27600
rect 34259 27595 34329 27600
rect 25391 27508 25457 27511
rect 37203 27508 37273 27513
rect 25391 27506 37208 27508
rect 25391 27450 25396 27506
rect 25452 27450 37208 27506
rect 25391 27448 37208 27450
rect 37268 27448 37273 27508
rect 25391 27445 25457 27448
rect 37203 27443 37273 27448
rect 27499 27368 27565 27371
rect 37479 27368 37549 27373
rect 27499 27366 37484 27368
rect 27499 27310 27504 27366
rect 27560 27310 37484 27366
rect 27499 27308 37484 27310
rect 37544 27308 37549 27368
rect 27499 27305 27565 27308
rect 37479 27303 37549 27308
rect 25551 27228 25617 27231
rect 38123 27228 38193 27233
rect 25551 27226 38128 27228
rect 25551 27170 25556 27226
rect 25612 27170 38128 27226
rect 25551 27168 38128 27170
rect 38188 27168 38193 27228
rect 25551 27165 25617 27168
rect 38123 27163 38193 27168
rect 27671 27088 27737 27091
rect 38767 27088 38837 27093
rect 27671 27086 38772 27088
rect 27671 27030 27676 27086
rect 27732 27030 38772 27086
rect 27671 27028 38772 27030
rect 38832 27028 38837 27088
rect 27671 27025 27737 27028
rect 38767 27023 38837 27028
rect 23632 26947 23698 26950
rect 39411 26947 39481 26952
rect 23632 26945 39416 26947
rect 23632 26889 23637 26945
rect 23693 26889 39416 26945
rect 23632 26887 39416 26889
rect 39476 26887 39481 26947
rect 23632 26884 23698 26887
rect 39411 26882 39481 26887
rect 21503 26814 21569 26817
rect 40055 26814 40125 26819
rect 21503 26812 40060 26814
rect 21503 26756 21508 26812
rect 21564 26756 40060 26812
rect 21503 26754 40060 26756
rect 40120 26754 40125 26814
rect 21503 26751 21569 26754
rect 40055 26749 40125 26754
rect 24317 26682 24383 26685
rect 40430 26682 40500 26687
rect 24317 26680 40435 26682
rect 24317 26624 24322 26680
rect 24378 26624 40435 26680
rect 24317 26622 40435 26624
rect 40495 26622 40500 26682
rect 24317 26619 24383 26622
rect 40430 26617 40500 26622
rect 35547 26531 35617 26536
rect 30495 26524 30565 26529
rect 33849 26524 33915 26527
rect 30495 26464 30500 26524
rect 30560 26522 33915 26524
rect 30560 26466 33854 26522
rect 33910 26466 33915 26522
rect 35547 26471 35552 26531
rect 35612 26516 43293 26531
rect 35612 26471 42093 26516
rect 35547 26466 35617 26471
rect 30560 26464 33915 26466
rect 30495 26459 30565 26464
rect 33849 26461 33915 26464
rect 42084 26460 42093 26471
rect 42149 26471 43293 26516
rect 42149 26460 42158 26471
rect 42084 26451 42158 26460
rect 30650 26370 30720 26375
rect 35938 26370 36004 26373
rect 30650 26310 30655 26370
rect 30715 26368 36004 26370
rect 30715 26312 35943 26368
rect 35999 26312 36004 26368
rect 30715 26310 36004 26312
rect 30650 26305 30720 26310
rect 35938 26307 36004 26310
rect 30803 26202 30873 26207
rect 34002 26202 34068 26205
rect 30803 26142 30808 26202
rect 30868 26200 34068 26202
rect 30868 26144 34007 26200
rect 34063 26144 34068 26200
rect 42104 26198 42178 26207
rect 30868 26142 34068 26144
rect 30803 26137 30873 26142
rect 34002 26139 34068 26142
rect 36191 26181 36261 26186
rect 42104 26181 42113 26198
rect 36191 26121 36196 26181
rect 36256 26142 42113 26181
rect 42169 26181 42178 26198
rect 42169 26142 43293 26181
rect 36256 26121 43293 26142
rect 36191 26116 36261 26121
rect 30938 26029 31008 26034
rect 36125 26029 36191 26032
rect 30938 25969 30943 26029
rect 31003 26027 36191 26029
rect 31003 25971 36130 26027
rect 36186 25971 36191 26027
rect 31003 25969 36191 25971
rect 30938 25964 31008 25969
rect 36125 25966 36191 25969
rect 42096 25884 42170 25893
rect 31104 25870 31174 25875
rect 33615 25873 33685 25878
rect 42096 25873 42105 25884
rect 31892 25870 31958 25873
rect 31104 25810 31109 25870
rect 31169 25868 31958 25870
rect 31169 25812 31897 25868
rect 31953 25812 31958 25868
rect 31169 25810 31958 25812
rect 31104 25805 31174 25810
rect 31892 25807 31958 25810
rect 33615 25813 33620 25873
rect 33680 25828 42105 25873
rect 42161 25873 42170 25884
rect 42161 25828 43293 25873
rect 33680 25813 43293 25828
rect 33615 25808 33685 25813
rect 29956 25717 30026 25722
rect 38015 25717 38081 25720
rect 29956 25657 29961 25717
rect 30021 25715 38081 25717
rect 30021 25659 38020 25715
rect 38076 25659 38081 25715
rect 30021 25657 38081 25659
rect 29956 25652 30026 25657
rect 38015 25654 38081 25657
rect 29778 23850 29844 23853
rect 30259 23850 30329 23855
rect 29778 23848 30264 23850
rect 29778 23792 29783 23848
rect 29839 23792 30264 23848
rect 29778 23790 30264 23792
rect 30324 23790 30329 23850
rect 29778 23787 29844 23790
rect 30259 23785 30329 23790
rect 38217 23794 38291 23799
rect 42040 23794 42106 23795
rect 38217 23730 38222 23794
rect 38286 23790 43293 23794
rect 38286 23734 42045 23790
rect 42101 23734 43293 23790
rect 38286 23730 43293 23734
rect 38217 23725 38291 23730
rect 42040 23729 42106 23730
rect 14073 23696 14147 23701
rect 14946 23696 15012 23697
rect 14073 23632 14078 23696
rect 14142 23692 15012 23696
rect 14142 23636 14951 23692
rect 15007 23636 15012 23692
rect 14142 23632 15012 23636
rect 14073 23627 14147 23632
rect 14946 23631 15012 23632
rect 38013 23197 38083 23202
rect 42148 23197 42214 23200
rect 38013 23137 38018 23197
rect 38078 23195 43293 23197
rect 38078 23139 42153 23195
rect 42209 23139 43293 23195
rect 38078 23137 43293 23139
rect 38013 23132 38083 23137
rect 42148 23134 42214 23137
rect 29771 22335 29837 22338
rect 30105 22335 30175 22340
rect 29771 22333 30110 22335
rect 29771 22277 29776 22333
rect 29832 22277 30110 22333
rect 29771 22275 30110 22277
rect 30170 22275 30175 22335
rect 29771 22272 29837 22275
rect 30105 22270 30175 22275
rect 30376 22306 30446 22311
rect 31887 22306 31953 22309
rect 30376 22246 30381 22306
rect 30441 22304 31953 22306
rect 30441 22248 31892 22304
rect 31948 22248 31953 22304
rect 30441 22246 31953 22248
rect 30376 22241 30446 22246
rect 31887 22243 31953 22246
rect 4284 7138 4350 7143
rect 4284 7082 4289 7138
rect 4345 7082 4350 7138
rect 4284 7077 4350 7082
rect 15256 4203 15322 4206
rect 19925 4203 19995 4208
rect 15256 4201 19930 4203
rect 15256 4145 15261 4201
rect 15317 4145 19930 4201
rect 15256 4143 19930 4145
rect 19990 4143 19995 4203
rect 15256 4140 15322 4143
rect 19925 4138 19995 4143
rect 18491 3531 18561 3536
rect 19681 3531 19747 3534
rect 18491 3471 18496 3531
rect 18556 3529 19747 3531
rect 18556 3473 19686 3529
rect 19742 3473 19747 3529
rect 18556 3471 19747 3473
rect 18491 3466 18561 3471
rect 19681 3468 19747 3471
rect 488 -110 898 -105
rect 488 -207 493 -110
rect -1604 -213 493 -207
rect -1604 -601 -218 -213
rect 170 -510 493 -213
rect 893 -207 898 -110
rect 893 -213 43293 -207
rect 893 -510 41519 -213
rect 170 -601 41519 -510
rect 41907 -601 43293 -213
rect -1604 -607 43293 -601
rect -1604 -673 43293 -667
rect -1604 -1061 -678 -673
rect -290 -707 41979 -673
rect -290 -1039 28 -707
rect 383 -1039 41979 -707
rect -290 -1061 41979 -1039
rect 42367 -1061 43293 -673
rect -1604 -1067 43293 -1061
rect -1604 -1133 43293 -1127
rect -1604 -1521 -1138 -1133
rect -750 -1190 42439 -1133
rect -750 -1254 4456 -1190
rect 4520 -1254 42439 -1190
rect -750 -1521 42439 -1254
rect 42827 -1521 43293 -1133
rect -1604 -1527 43293 -1521
rect -1604 -1593 43293 -1587
rect -1604 -1981 -1598 -1593
rect -1210 -1981 42899 -1593
rect 43287 -1981 43293 -1593
rect -1604 -1987 43293 -1981
<< via3 >>
rect -1598 40888 -1210 41276
rect 34593 40909 34911 41227
rect 42899 40888 43287 41276
rect -1138 40428 -750 40816
rect 35253 40461 35571 40779
rect 42439 40428 42827 40816
rect -678 39968 -290 40356
rect 41979 39968 42367 40356
rect -218 39508 170 39896
rect 41519 39508 41907 39896
rect -218 -601 170 -213
rect 41519 -601 41907 -213
rect -678 -1061 -290 -673
rect 41979 -1061 42367 -673
rect -1138 -1521 -750 -1133
rect 42439 -1521 42827 -1133
rect -1598 -1981 -1210 -1593
rect 42899 -1981 43287 -1593
<< metal4 >>
rect -1604 41276 -1204 41283
rect -1604 40888 -1598 41276
rect -1210 40888 -1204 41276
rect -1604 -1593 -1204 40888
rect -1604 -1981 -1598 -1593
rect -1210 -1981 -1204 -1593
rect -1604 -1987 -1204 -1981
rect -1144 40816 -744 41283
rect -1144 40428 -1138 40816
rect -750 40428 -744 40816
rect -1144 -1133 -744 40428
rect -1144 -1521 -1138 -1133
rect -750 -1521 -744 -1133
rect -1144 -1987 -744 -1521
rect -684 40356 -284 41283
rect -684 39968 -678 40356
rect -290 39968 -284 40356
rect -684 -673 -284 39968
rect -684 -1061 -678 -673
rect -290 -1061 -284 -673
rect -684 -1987 -284 -1061
rect -224 39896 176 41283
rect -224 39508 -218 39896
rect 170 39508 176 39896
rect -224 7639 176 39508
rect 34592 41227 34912 41228
rect 34592 40909 34593 41227
rect 34911 40909 34912 41227
rect 34592 36728 34912 40909
rect 35252 40779 35572 40780
rect 35252 40461 35253 40779
rect 35571 40461 35572 40779
rect 35252 36621 35572 40461
rect 41513 39896 41913 41283
rect 41513 39508 41519 39896
rect 41907 39508 41913 39896
rect -224 7237 180 7639
rect -224 -213 176 7237
rect -224 -601 -218 -213
rect 170 -601 176 -213
rect -224 -1987 176 -601
rect 41513 -213 41913 39508
rect 41513 -601 41519 -213
rect 41907 -601 41913 -213
rect 41513 -1987 41913 -601
rect 41973 40356 42373 41283
rect 41973 39968 41979 40356
rect 42367 39968 42373 40356
rect 41973 -673 42373 39968
rect 41973 -1061 41979 -673
rect 42367 -1061 42373 -673
rect 41973 -1987 42373 -1061
rect 42433 40816 42833 41283
rect 42433 40428 42439 40816
rect 42827 40428 42833 40816
rect 42433 -1133 42833 40428
rect 42433 -1521 42439 -1133
rect 42827 -1521 42833 -1133
rect 42433 -1987 42833 -1521
rect 42893 41276 43293 41283
rect 42893 40888 42899 41276
rect 43287 40888 43293 41276
rect 42893 -1593 43293 40888
rect 42893 -1981 42899 -1593
rect 43287 -1981 43293 -1593
rect 42893 -1987 43293 -1981
use brownout_ana  brownout_ana_0 ~/chipalooza/sky130_ajc_ip__brownout/mag
timestamp 1712959001
transform 1 0 29373 0 1 25849
box -29373 -25849 12300 13900
use brownout_dig  brownout_dig_0 ~/chipalooza/sky130_ajc_ip__brownout/mag
timestamp 1712954807
transform 1 0 30384 0 1 26140
box 0 0 11173 13317
use sky130_fd_pr__nfet_g5v0d10v5_PXF6AN  sky130_fd_pr__nfet_g5v0d10v5_PXF6AN_0
timestamp 1712947988
transform 0 1 42123 -1 0 26332
box -1463 -358 1463 358
use sky130_fd_pr__nfet_g5v0d10v5_V6EN4F  sky130_fd_pr__nfet_g5v0d10v5_V6EN4F_0
timestamp 1712949175
transform 1 0 4317 0 1 311
box -357 -358 357 358
use sky130_fd_pr__nfet_g5v0d10v5_XTZQRT  sky130_fd_pr__nfet_g5v0d10v5_XTZQRT_0
timestamp 1712945108
transform 1 0 28810 0 1 37759
box -989 -358 989 358
<< labels >>
flabel metal3 1723 -1527 1723 -1527 0 FreeSans 1600 0 0 0 dvss
port 6 nsew
flabel metal3 1723 -1987 1723 -1987 0 FreeSans 1600 0 0 0 dvdd
port 4 nsew
flabel metal3 s 43093 30259 43293 30318 0 FreeSans 1600 0 0 0 force_dis_rc_osc
port 21 nsew
flabel metal3 s 43093 31618 43293 31678 0 FreeSans 1600 0 0 0 force_ena_rc_osc
port 19 nsew
flabel metal3 s 43093 33658 43293 33718 0 FreeSans 1600 0 0 0 force_short_oneshot
port 24 nsew
flabel metal3 s 43093 34338 43293 34398 0 FreeSans 1600 0 0 0 timed_out
port 22 nsew
flabel metal2 s 38788 41082 38816 41282 0 FreeSans 1600 90 0 0 vtrip[0]
port 16 nsew
flabel metal2 s 32992 41082 33020 41282 0 FreeSans 1600 90 0 0 vtrip[2]
port 14 nsew
flabel metal2 s 32348 41082 32376 41282 0 FreeSans 1600 90 0 0 vtrip[1]
port 15 nsew
flabel metal3 s 43093 25813 43293 25873 0 FreeSans 1600 0 0 0 otrip[0]
port 11 nsew
flabel metal3 s 43093 26471 43293 26531 0 FreeSans 1600 0 0 0 otrip[1]
port 10 nsew
flabel metal3 s 43093 26121 43293 26181 0 FreeSans 1600 0 0 0 otrip[2]
port 9 nsew
flabel metal3 s 43093 23730 43293 23794 0 FreeSans 1600 0 0 0 isrc_sel
port 25 nsew
flabel metal3 s 43093 23137 43293 23197 0 FreeSans 1600 0 0 0 ena
port 18 nsew
flabel metal2 s 10947 41082 11011 41282 0 FreeSans 1600 90 0 0 vbg_1v2
port 8 nsew
flabel metal2 s 14947 41082 15011 41282 0 FreeSans 1600 90 0 0 ibg_200n
port 26 nsew
flabel metal2 s 26956 41082 27008 41282 0 FreeSans 1600 90 0 0 outb
port 3 nsew
flabel metal2 s 27692 41082 27752 41282 0 FreeSans 1600 90 0 0 osc_ck
port 5 nsew
flabel metal3 s 43093 32298 43293 32358 0 FreeSans 1600 0 0 0 dcomp
port 7 nsew
flabel metal2 s 29742 41082 29802 41282 0 FreeSans 1600 90 0 0 brout_filt
port 13 nsew
flabel metal2 s 12176 41082 12236 41282 0 FreeSans 1600 90 0 0 vin_brout
port 17 nsew
flabel metal2 s 4287 -1987 4347 -1787 0 FreeSans 1600 90 0 0 vin_vunder
port 20 nsew
flabel metal2 s 27302 41082 27358 41282 0 FreeSans 1600 90 0 0 vunder
port 23 nsew
flabel metal3 1723 -607 1723 -607 0 FreeSans 1600 0 0 0 avss
port 2 nsew
flabel metal3 1723 -1067 1723 -1067 0 FreeSans 1600 0 0 0 avdd
port 1 nsew
flabel metal2 11863 41082 11915 41282 0 FreeSans 1600 90 0 0 itest
port 12 nsew
<< end >>
