* NGSPICE file created from por_ana_rcx.ext - technology: sky130A

.subckt por_ana_rcx otrip_decoded[1] otrip_decoded[0] itest ibg_200n osc_ck porb_h
+ por porb force_pdnb otrip_decoded[7] otrip_decoded[4] isrc_sel otrip_decoded[5]
+ otrip_decoded[2] vin vbg_1v2 pwup_filt dcomp por_unbuf otrip_decoded[3] otrip_decoded[6]
+ avss dvdd dvss avdd osc_ena
X0 a_n3778_7859# a_n3878_7771# dvss.t533 dvss.t532 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X1 a_8447_n11914# a_8069_n19314# avss.t132 sky130_fd_pr__res_xhigh_po_1p41 l=35
X2 avss.t40 comparator_1.n1 dcomp3v3 avss.t39 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.6
X3 comparator_1.vt avss.t410 comparator_1.vnn comparator_1.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=8
X4 a_n15745_n11914# a_n16123_n19314# avss.t43 sky130_fd_pr__res_xhigh_po_1p41 l=35
X5 rstring_mux_0.vtrip4.t2 rstring_mux_0.vtrip_decoded_avdd[4] comparator_0.vinn.t2 avss.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X6 avdd.t33 comparator_1.n1 dcomp3v3 avdd.t32 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X7 dvdd.t171 sky130_fd_sc_hd__inv_4_1.Y porb.t31 dvdd.t170 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 rstring_mux_0.vtrip_decoded_b_avdd[7] rstring_mux_0.vtrip_decoded_avdd[7] avss.t268 avss.t267 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X9 dvdd.t325 dvdd.t323 osc_ck.t7 dvdd.t324 sky130_fd_pr__pfet_01v8 ad=0.1475 pd=1.295 as=0.15 ps=1.3 w=1 l=0.18
X10 a_5346_n3990# a_4921_n3946# dvss.t110 dvss.t109 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X11 rc_osc_0.n.t5 dvdd.t321 rc_osc_0.m dvdd.t322 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X12 dvdd.t41 sky130_fd_sc_hd__inv_4_0.Y pwup_filt.t31 dvdd.t40 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13 avdd.t399 a_429_n2876# a_1122_n3990# avdd.t398 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.1365 ps=1.49 w=0.42 l=1
X14 rstring_mux_0.vtop.t17 a_n16123_n19314# avss.t323 sky130_fd_pr__res_xhigh_po_1p41 l=35
X15 comparator_0.vn avss.t230 comparator_0.ibias avss.t231 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X16 avss.t229 avss.t228 avss.t229 avss.t136 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=8
X17 dvss.t539 otrip_decoded[0].t0 a_n8119_n2964# dvss.t538 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X18 comparator_1.vpp rstring_mux_0.ena avdd.t528 avdd.t527 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X19 comparator_1.n0 comparator_1.vpp avdd.t652 avdd.t73 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X20 dvss.t720 a_7033_n3946# a_7458_n3990# dvss.t719 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X21 rstring_mux_0.otrip_decoded_b_avdd[1] rstring_mux_0.otrip_decoded_avdd[1] avss.t301 avss.t300 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X22 vin avdd.t394 vin avdd.t395 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=23.2 ps=169.28 w=5 l=0.6
X23 comparator_1.vt vbg_1v2.t0 comparator_1.vnn comparator_1.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X24 comparator_1.vpp comparator_1.vnn avdd.t90 avdd.t63 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X25 dcomp.t31 sky130_fd_sc_hd__inv_4_3.Y dvdd.t312 dvdd.t311 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X26 dvdd.t93 schmitt_trigger_0.in.t1 schmitt_trigger_0.m.t12 dvdd.t92 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X27 comparator_0.vnn comparator_0.vinn.t48 comparator_0.vt comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X28 a_3155_n11914# a_3533_n19314# avss.t244 sky130_fd_pr__res_xhigh_po_1p41 l=35
X29 a_n11209_n11914# a_n10831_n19314# avss.t394 sky130_fd_pr__res_xhigh_po_1p41 l=35
X30 comparator_1.vpp vin comparator_1.vt comparator_1.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X31 rstring_mux_0.otrip_decoded_avdd[5] a_n2588_n1478# avdd.t621 avdd.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.24375 ps=1.825 w=1.5 l=0.5
X32 dvdd.t280 a_10873_n2760# a_10873_n3956# dvdd.t278 sky130_fd_pr__pfet_01v8_hvt ad=0.2968 pd=2.77 as=0.2968 ps=2.77 w=1.12 l=0.15
X33 a_7458_n3990# a_7033_n3946# dvss.t718 dvss.t717 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X34 comparator_1.vpp comparator_1.vnn avdd.t89 avdd.t63 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X35 ibias_gen_0.vr.t4 ibias_gen_0.vn0.t19 ibias_gen_0.vp0.t11 avss.t67 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X36 avdd.t594 a_2541_n2876# a_3234_n3990# avdd.t593 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.1365 ps=1.49 w=0.42 l=1
X37 comparator_0.vpp comparator_0.vnn avdd.t204 avdd.t177 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X38 a_n26830_n2937# a_n27208_n10337# avss.t0 sky130_fd_pr__res_xhigh_po_1p41 l=35
X39 dvdd.t273 sky130_fd_sc_hd__inv_4_4.Y por.t31 dvdd.t272 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X40 dvss.t648 a_9145_n3946# a_9570_n3990# dvss.t647 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X41 comparator_0.vt comparator_0.vinn.t49 comparator_0.vnn comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X42 porb_h.t15 sky130_fd_sc_hvl__inv_16_0.A avss.t373 avss.t372 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X43 rstring_mux_0.vtrip_decoded_avdd[0] a_1636_n3212# dvss.t694 dvss.t693 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.121875 ps=1.075 w=0.75 l=0.5
X44 dvss.t114 a_6765_n2876# a_7972_n3212# dvss.t113 sky130_fd_pr__nfet_g5v0d10v5 ad=0.121875 pd=1.075 as=0.19875 ps=2.03 w=0.75 l=0.5
X45 avdd.t535 ibias_gen_0.isrc_sel ibias_gen_0.isrc_sel_b avdd.t534 sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=1
X46 a_n8951_9395# a_n8573_1995# avss.t310 sky130_fd_pr__res_xhigh_po_1p41 l=35
X47 itest.t1 ibias_gen_0.vp.t7 avdd.t425 avdd.t424 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X48 comparator_0.vinn.t47 avdd.t392 comparator_0.vinn.t47 avdd.t393 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=0.6
X49 comparator_1.vt vin comparator_1.vpp comparator_1.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X50 rstring_mux_0.vtrip7.t7 a_n247_n19314# avss.t269 sky130_fd_pr__res_xhigh_po_1p41 l=35
X51 dvss.t88 sky130_fd_sc_hd__inv_4_0.Y pwup_filt.t15 dvss.t87 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X52 comparator_1.vt vin comparator_1.vpp comparator_1.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X53 a_n24562_n2937# a_n24184_n10337# avss.t0 sky130_fd_pr__res_xhigh_po_1p41 l=35
X54 a_n21538_n2937# a_n21160_n10337# avss.t0 sky130_fd_pr__res_xhigh_po_1p41 l=35
X55 avdd.t626 a_4653_n2876# a_5346_n3990# avdd.t625 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.1365 ps=1.49 w=0.42 l=1
X56 vin avdd.t390 vin avdd.t391 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=0.6
X57 dvdd.t271 sky130_fd_sc_hd__inv_4_4.Y por.t30 dvdd.t270 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X58 rstring_mux_0.otrip_decoded_b_avdd[2] rstring_mux_0.otrip_decoded_avdd[2] avss.t341 avss.t340 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X59 a_6935_n11914# a_6557_n19314# avss.t322 sky130_fd_pr__res_xhigh_po_1p41 l=35
X60 avdd.t569 sky130_fd_sc_hvl__inv_16_0.A porb_h.t31 avdd.t568 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X61 avss.t331 rstring_mux_0.ena rstring_mux_0.ena_b avss.t330 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X62 a_n26830_n2937# a_n26452_n10337# avss.t0 sky130_fd_pr__res_xhigh_po_1p41 l=35
X63 a_n23806_n2937# a_n23428_n10337# avss.t0 sky130_fd_pr__res_xhigh_po_1p41 l=35
X64 comparator_0.vpp comparator_0.vnn avdd.t203 avdd.t177 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X65 rstring_mux_0.vtrip2.t7 rstring_mux_0.vtrip_decoded_avdd[2] comparator_0.vinn.t44 avss.t381 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X66 por.t15 sky130_fd_sc_hd__inv_4_4.Y dvss.t680 dvss.t679 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X67 rstring_mux_0.vtrip_decoded_avdd[2] a_3748_n3212# dvss.t692 dvss.t691 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.121875 ps=1.075 w=0.75 l=0.5
X68 a_n7326_n3990# a_n7751_n3946# dvss.t690 dvss.t689 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X69 a_6935_n11914# a_7313_n19314# avss.t387 sky130_fd_pr__res_xhigh_po_1p41 l=35
X70 a_n14989_n11914# a_n14611_n19314# avss.t321 sky130_fd_pr__res_xhigh_po_1p41 l=35
X71 a_n3649_n11914# a_n4027_n19314# avss.t251 sky130_fd_pr__res_xhigh_po_1p41 l=35
X72 dvdd.t241 vl sky130_fd_sc_hd__inv_4_3.Y dvdd.t240 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X73 avdd.t15 a_n3795_n1142# a_n2588_n1478# avdd.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0.24375 pd=1.825 as=0.3975 ps=3.53 w=1.5 l=0.5
X74 sky130_fd_sc_hvl__inv_1_0.A a_n2571_7523# dvss.t696 dvss.t695 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.121875 ps=1.075 w=0.75 l=0.5
X75 dvss.t758 sky130_fd_sc_hd__inv_4_3.Y dcomp.t15 dvss.t757 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X76 comparator_0.vnn comparator_0.vpp avdd.t618 avdd.t186 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X77 a_n4405_n11914# a_n4027_n19314# avss.t250 sky130_fd_pr__res_xhigh_po_1p41 l=35
X78 ibias_gen_0.vp1.t14 ibias_gen_0.vp1.t13 avdd.t98 avdd.t97 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X79 a_n15529_n2223# ibias_gen_0.isrc_sel_b ibias_gen_0.vn1.t7 avdd.t491 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X80 a_n1683_n1142# a_n1783_n1230# dvss.t613 dvss.t612 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X81 dvss.t319 dvss.t317 a_2441_n1230# dvss.t318 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X82 comparator_0.vpp comparator_0.vnn avdd.t202 avdd.t177 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X83 avdd.t493 a_n3102_n2256# a_n3795_n1142# avdd.t492 sky130_fd_pr__pfet_g5v0d10v5 ad=0.2142 pd=1.99 as=0.2142 ps=1.99 w=0.42 l=1
X84 avdd.t41 a_6765_n2876# a_7458_n3990# avdd.t40 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.1365 ps=1.49 w=0.42 l=1
X85 a_2809_n3946# a_2441_n2964# dvdd.t133 dvdd.t132 sky130_fd_pr__pfet_01v8_hvt ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X86 dvdd.t269 sky130_fd_sc_hd__inv_4_4.Y por.t29 dvdd.t268 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X87 dvdd.t169 sky130_fd_sc_hd__inv_4_1.Y porb.t30 dvdd.t168 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X88 dvss.t541 por_unbuf.t0 sky130_fd_sc_hd__inv_4_1.A dvss.t540 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X89 osc_ck.t2 osc_ena.t0 rc_osc_0.vr dvss.t477 sky130_fd_pr__nfet_01v8 ad=0.15 pd=1.3 as=0.1475 ps=1.295 w=1 l=0.18
X90 avdd.t201 comparator_0.vnn comparator_0.vnn avdd.t182 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X91 rstring_mux_0.otrip_decoded_b_avdd[6] rstring_mux_0.otrip_decoded_avdd[6] avdd.t495 avdd.t494 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X92 a_n10279_n24223# a_12321_n24601# dvss.t591 sky130_fd_pr__res_xhigh_po_1p41 l=111
X93 dcomp.t30 sky130_fd_sc_hd__inv_4_3.Y dvdd.t310 dvdd.t309 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X94 dvdd.t39 sky130_fd_sc_hd__inv_4_0.Y pwup_filt.t30 dvdd.t38 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X95 rstring_mux_0.vtrip3.t9 rstring_mux_0.vtrip_decoded_b_avdd[3] comparator_0.vinn.t36 avdd.t445 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X96 dvdd.t49 rc_osc_0.m rc_osc_0.n.t3 dvdd.t48 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X97 avss.t295 comparator_1.vn comparator_1.vn avss.t278 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X98 ibias_gen_0.vn0.t18 vbg_1v2.t1 ibias_gen_0.vstart.t10 avss.t128 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X99 rc_osc_0.m rc_osc_0.in dvdd.t219 dvdd.t218 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X100 ibias_gen_0.vr.t2 a_n20404_n10337# avss.t0 sky130_fd_pr__res_xhigh_po_1p41 l=35
X101 avdd.t439 a_n5907_n1142# a_n4700_n1478# avdd.t438 sky130_fd_pr__pfet_g5v0d10v5 ad=0.24375 pd=1.825 as=0.3975 ps=3.53 w=1.5 l=0.5
X102 comparator_1.ena_b rstring_mux_0.ena avdd.t526 avdd.t525 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X103 dvss.t521 sky130_fd_sc_hd__inv_4_1.Y porb.t15 dvss.t520 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X104 a_n13487_9395# a_n13109_1995# avss.t60 sky130_fd_pr__res_xhigh_po_1p41 l=35
X105 a_n3795_n1142# a_n3895_n1230# dvss.t373 dvss.t372 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X106 a_2541_n1142# a_2441_n1230# dvss.t52 dvss.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X107 a_7033_n3946# a_6665_n2964# dvdd.t127 dvdd.t126 sky130_fd_pr__pfet_01v8_hvt ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X108 sky130_fd_sc_hd__inv_4_1.Y sky130_fd_sc_hd__inv_4_1.A dvss.t599 dvss.t598 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X109 schmitt_trigger_0.m.t0 schmitt_trigger_0.out.t4 dvdd.t53 dvdd.t52 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X110 a_n14243_9395# a_n14621_1995# avss.t256 sky130_fd_pr__res_xhigh_po_1p41 l=35
X111 dvdd.t320 dvdd.t318 schmitt_trigger_0.m.t13 dvdd.t319 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X112 dvdd.t135 otrip_decoded[6].t0 a_n1783_n2964# dvdd.t134 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X113 avss.t38 comparator_1.n1 dcomp3v3 avss.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X114 dvss.t341 a_8877_n1142# a_10084_n1478# dvss.t175 sky130_fd_pr__nfet_g5v0d10v5 ad=0.121875 pd=1.075 as=0.19875 ps=2.03 w=0.75 l=0.5
X115 rstring_mux_0.vtrip_decoded_avdd[5] a_5860_n1478# avdd.t208 avdd.t207 sky130_fd_pr__pfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.24375 ps=1.825 w=1.5 l=0.5
X116 rstring_mux_0.otrip_decoded_b_avdd[1] rstring_mux_0.otrip_decoded_avdd[1] avdd.t487 avdd.t486 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X117 a_n7429_n11914# a_n7807_n19314# avss.t249 sky130_fd_pr__res_xhigh_po_1p41 l=35
X118 dvss.t710 a_2541_n2876# a_3748_n3212# dvss.t709 sky130_fd_pr__nfet_g5v0d10v5 ad=0.121875 pd=1.075 as=0.19875 ps=2.03 w=0.75 l=0.5
X119 comparator_0.vnn comparator_0.vpp avdd.t617 avdd.t186 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X120 avdd.t655 a_n8019_n1142# a_n6812_n1478# avdd.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=0.24375 pd=1.825 as=0.3975 ps=3.53 w=1.5 l=0.5
X121 dcomp3v3uv comparator_0.n1 avdd.t62 avdd.t61 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X122 comparator_0.vinn.t46 rstring_mux_0.vtrip_decoded_b_avdd[5] rstring_mux_0.vtrip5.t6 avdd.t579 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X123 rstring_mux_0.otrip_decoded_avdd[5] a_n2588_n1478# dvss.t722 dvss.t721 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.121875 ps=1.075 w=0.75 l=0.5
X124 avdd.t651 comparator_1.vpp comparator_1.vpp avdd.t65 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X125 a_4653_n1142# a_4553_n1230# dvss.t360 dvss.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X126 a_9145_n3946# a_8777_n2964# dvdd.t51 dvdd.t50 sky130_fd_pr__pfet_01v8_hvt ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X127 avdd.t200 comparator_0.vnn comparator_0.vnn avdd.t182 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X128 comparator_1.vt vbg_1v2.t2 comparator_1.vnn comparator_1.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X129 a_5423_n11914# a_5801_n19314# avss.t41 sky130_fd_pr__res_xhigh_po_1p41 l=35
X130 avdd.t88 comparator_1.vnn comparator_1.vpp avdd.t65 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X131 a_n3085_6745# a_n3510_6789# dvss.t456 dvss.t455 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X132 comparator_0.vnn comparator_0.vinn.t50 comparator_0.vt comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X133 dvss.t543 por_unbuf.t1 sky130_fd_sc_hd__inv_4_4.Y dvss.t542 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X134 dvdd.t69 otrip_decoded[4].t0 a_n3895_n2964# dvdd.t68 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X135 a_n11975_9395# a_n11597_1995# avss.t302 sky130_fd_pr__res_xhigh_po_1p41 l=35
X136 dvss.t86 sky130_fd_sc_hd__inv_4_0.Y pwup_filt.t14 dvss.t85 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X137 dvss.t316 dvss.t314 a_329_n1230# dvss.t315 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X138 a_697_n3946# a_329_n2964# dvdd.t43 dvdd.t42 sky130_fd_pr__pfet_01v8_hvt ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X139 avdd.t389 avdd.t387 avdd.t388 avdd.t221 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=8
X140 comparator_0.vpp comparator_0.vpp avdd.t616 avdd.t177 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X141 rstring_mux_0.vtrip1.t2 rstring_mux_0.vtrip2.t0 avss.t42 sky130_fd_pr__res_xhigh_po_1p41 l=35
X142 dvss.t313 dvss.t311 osc_ck.t1 dvss.t312 sky130_fd_pr__nfet_01v8 ad=0.1475 pd=1.295 as=0.15 ps=1.3 w=1 l=0.18
X143 comparator_1.vm comparator_1.vm avss.t285 avss.t284 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X144 dvdd.t267 sky130_fd_sc_hd__inv_4_4.Y por.t28 dvdd.t266 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X145 avdd.t443 a_429_n1142# a_1636_n1478# avdd.t442 sky130_fd_pr__pfet_g5v0d10v5 ad=0.24375 pd=1.825 as=0.3975 ps=3.53 w=1.5 l=0.5
X146 dvss.t724 a_4653_n2876# a_5860_n3212# dvss.t723 sky130_fd_pr__nfet_g5v0d10v5 ad=0.121875 pd=1.075 as=0.19875 ps=2.03 w=0.75 l=0.5
X147 avdd.t485 rstring_mux_0.ena_b rstring_mux_0.vtop.t16 avdd.t484 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X148 avdd.t421 comparator_0.n0 comparator_0.n1 avdd.t420 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X149 avdd.t199 comparator_0.vnn comparator_0.vpp avdd.t179 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X150 comparator_1.vpp comparator_1.vnn avdd.t87 avdd.t63 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X151 dvdd.t55 schmitt_trigger_0.out.t5 schmitt_trigger_0.m.t1 dvdd.t54 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X152 ibias_gen_0.vp0.t9 ibias_gen_0.vp0.t8 avdd.t403 avdd.t402 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X153 por.t14 sky130_fd_sc_hd__inv_4_4.Y dvss.t678 dvss.t677 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X154 rstring_mux_0.otrip_decoded_avdd[3] a_n4700_n1478# dvss.t571 dvss.t570 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.121875 ps=1.075 w=0.75 l=0.5
X155 avdd.t386 avdd.t385 avdd.t386 avdd.t240 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=8
X156 a_6765_n1142# a_6665_n1230# dvss.t588 dvss.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X157 rstring_mux_0.vtop.t15 rstring_mux_0.ena_b avdd.t483 avdd.t482 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X158 ibias_gen_0.ena_b rstring_mux_0.ena avss.t329 avss.t328 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=1
X159 rstring_mux_0.otrip_decoded_avdd[2] a_n4700_n3212# avdd.t417 avdd.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.24375 ps=1.825 w=1.5 l=0.5
X160 dvdd.t187 otrip_decoded[2].t0 a_n6007_n2964# dvdd.t186 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X161 vin rstring_mux_0.otrip_decoded_b_avdd[6] rstring_mux_0.vtrip6.t6 avdd.t451 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X162 avdd.t650 comparator_1.vpp comparator_1.vpp avdd.t65 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X163 porb_h.t14 sky130_fd_sc_hvl__inv_16_0.A avss.t371 avss.t370 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X164 avss.t227 avss.t225 avss.t226 avss.t146 sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0 ps=0 w=5 l=8
X165 dvss.t84 sky130_fd_sc_hd__inv_4_0.Y pwup_filt.t13 dvss.t83 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X166 a_10873_n2760# a_10514_n2760# dvss.t568 dvss.t565 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.105 ps=1.03 w=0.75 l=0.5
X167 a_887_n11914# a_509_n19314# avss.t386 sky130_fd_pr__res_xhigh_po_1p41 l=35
X168 comparator_0.vnn comparator_0.vpp avdd.t615 avdd.t186 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X169 avdd.t198 comparator_0.vnn comparator_0.vnn avdd.t182 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X170 ibias_gen_0.vp.t4 rstring_mux_0.ena avdd.t524 avdd.t523 sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=2
X171 avdd.t423 a_1122_n2256# a_429_n1142# avdd.t422 sky130_fd_pr__pfet_g5v0d10v5 ad=0.2142 pd=1.99 as=0.2142 ps=1.99 w=0.42 l=1
X172 osc_ck.t3 rc_osc_0.n.t6 dvss.t535 dvss.t534 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X173 avdd.t481 rstring_mux_0.ena_b rstring_mux_0.vtop.t14 avdd.t480 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X174 dvdd.t265 sky130_fd_sc_hd__inv_4_4.Y por.t27 dvdd.t264 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X175 comparator_0.vt vbg_1v2.t3 comparator_0.vpp comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X176 avdd.t427 ibias_gen_0.vp.t8 ibias_gen_0.ibias0 avdd.t426 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X177 dvss.t138 dcomp3v3uv a_10514_n2760# dvss.t137 sky130_fd_pr__nfet_g5v0d10v5 ad=0.178875 pd=1.26 as=0.1197 ps=1.41 w=0.42 l=0.5
X178 rstring_mux_0.vtrip_decoded_b_avdd[0] rstring_mux_0.vtrip_decoded_avdd[0] avss.t377 avss.t376 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X179 comparator_1.n1 comparator_1.n0 avss.t385 avss.t384 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.6
X180 ibias_gen_0.vn0.t6 ibias_gen_0.vn0.t5 ibias_gen_0.ve.t4 avss.t67 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X181 ibias_gen_0.vp.t3 ibias_gen_0.isrc_sel_b ibias_gen_0.vp0.t3 avss.t305 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X182 avss.t393 comparator_0.vn comparator_0.vt avss.t109 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X183 avdd.t384 avdd.t382 avdd.t383 avdd.t221 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=8
X184 comparator_0.vinn.t33 avdd.t380 vin avdd.t381 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X185 avss.t369 sky130_fd_sc_hvl__inv_16_0.A porb_h.t13 avss.t368 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X186 rstring_mux_0.vtop.t13 rstring_mux_0.ena_b avdd.t479 avdd.t478 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X187 comparator_1.vpp comparator_1.vnn avdd.t86 avdd.t63 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X188 ibias_gen_0.vp1.t0 ibias_gen_0.vn1.t10 avss.t119 avss.t117 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=8
X189 a_n5917_n11914# a_n6295_n19314# avss.t320 sky130_fd_pr__res_xhigh_po_1p41 l=35
X190 avdd.t197 comparator_0.vnn comparator_0.vpp avdd.t179 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X191 a_n7751_n2212# a_n8119_n1230# dvss.t626 dvss.t625 sky130_fd_pr__nfet_01v8 ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X192 rstring_mux_0.otrip_decoded_avdd[0] a_n6812_n3212# avdd.t499 avdd.t498 sky130_fd_pr__pfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.24375 ps=1.825 w=1.5 l=0.5
X193 rstring_mux_0.vtrip_decoded_b_avdd[4] rstring_mux_0.vtrip_decoded_avdd[4] avss.t23 avss.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X194 dvss.t82 sky130_fd_sc_hd__inv_4_0.Y pwup_filt.t12 dvss.t81 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X195 dvss.t519 sky130_fd_sc_hd__inv_4_1.Y porb.t14 dvss.t518 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X196 dvdd.t189 otrip_decoded[0].t1 a_n8119_n2964# dvdd.t188 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X197 vin rstring_mux_0.otrip_decoded_b_avdd[1] rstring_mux_0.vtrip1.t7 avdd.t414 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X198 rc_osc_0.in a_12321_n25357# dvss.t614 sky130_fd_pr__res_xhigh_po_1p41 l=111
X199 avdd.t567 sky130_fd_sc_hvl__inv_16_0.A porb_h.t30 avdd.t566 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X200 dcomp3v3 comparator_1.n1 avdd.t31 avdd.t30 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X201 sky130_fd_sc_hd__inv_4_1.Y sky130_fd_sc_hd__inv_4_1.A dvss.t597 dvss.t596 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X202 rstring_mux_0.vtrip_decoded_avdd[1] a_1636_n1478# avdd.t448 avdd.t442 sky130_fd_pr__pfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.24375 ps=1.825 w=1.5 l=0.5
X203 avdd.t504 a_6765_n1142# a_7972_n1478# avdd.t101 sky130_fd_pr__pfet_g5v0d10v5 ad=0.24375 pd=1.825 as=0.3975 ps=3.53 w=1.5 l=0.5
X204 avdd.t100 a_3234_n2256# a_2541_n1142# avdd.t99 sky130_fd_pr__pfet_g5v0d10v5 ad=0.2142 pd=1.99 as=0.2142 ps=1.99 w=0.42 l=1
X205 a_n8195_9395# schmitt_trigger_0.in.t0 avss.t71 sky130_fd_pr__res_xhigh_po_1p41 l=35
X206 rc_osc_0.vr dvdd.t316 rc_osc_0.ena_b dvdd.t317 sky130_fd_pr__pfet_01v8 ad=0.1475 pd=1.295 as=0.145 ps=1.29 w=1 l=0.5
X207 vin rstring_mux_0.otrip_decoded_avdd[0] rstring_mux_0.vtrip0.t5 avss.t314 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X208 comparator_0.vnn comparator_0.vpp avdd.t614 avdd.t186 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X209 a_n8951_9395# a_n9329_1995# avss.t315 sky130_fd_pr__res_xhigh_po_1p41 l=35
X210 avss.t224 avss.t222 avss.t223 avss.t146 sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0 ps=0 w=5 l=8
X211 dcomp.t29 sky130_fd_sc_hd__inv_4_3.Y dvdd.t308 dvdd.t307 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X212 vin avdd.t378 vin avdd.t379 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=0.6
X213 avdd.t85 comparator_1.vnn comparator_1.vnn avdd.t80 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X214 dvdd.t115 dvss.t770 a_2441_n1230# dvdd.t114 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X215 rstring_mux_0.otrip_decoded_b_avdd[4] rstring_mux_0.otrip_decoded_avdd[4] avss.t79 avss.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X216 avdd.t377 avdd.t376 avdd.t377 avdd.t240 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=8
X217 comparator_0.vinn.t34 avdd.t374 comparator_0.vinn.t34 avdd.t375 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=0.6
X218 avdd.t429 ibias_gen_0.vp.t9 itest.t0 avdd.t428 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X219 vin rstring_mux_0.otrip_decoded_avdd[4] rstring_mux_0.vtrip4.t6 avss.t77 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X220 avdd.t649 comparator_1.vpp comparator_1.vpp avdd.t65 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X221 porb_h.t29 sky130_fd_sc_hvl__inv_16_0.A avdd.t565 avdd.t564 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X222 ibias_gen_0.vstart.t9 vbg_1v2.t4 ibias_gen_0.vn0.t17 avss.t128 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X223 ibias_gen_0.isrc_sel_b avss.t220 ibias_gen_0.ena_b avss.t221 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X224 a_n1683_n1142# a_n1783_n1230# dvss.t611 dvss.t610 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X225 comparator_1.vn rstring_mux_0.ena ibias_gen_0.ibias0 avss.t327 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X226 comparator_0.vnn comparator_0.vpp avdd.t613 avdd.t186 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X227 comparator_1.vt vbg_1v2.t5 comparator_1.vnn comparator_1.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X228 comparator_0.vnn comparator_0.vinn.t51 comparator_0.vt comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X229 dvss.t531 a_n3878_7771# a_n3778_7859# dvss.t530 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X230 a_n20782_n2937# a_n21160_n10337# avss.t0 sky130_fd_pr__res_xhigh_po_1p41 l=35
X231 rstring_mux_0.vtrip_decoded_avdd[3] a_3748_n1478# avdd.t108 avdd.t107 sky130_fd_pr__pfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.24375 ps=1.825 w=1.5 l=0.5
X232 comparator_0.vnn comparator_0.vinn.t52 comparator_0.vt comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X233 dvss.t676 sky130_fd_sc_hd__inv_4_4.Y por.t13 dvss.t675 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X234 avdd.t104 a_5346_n2256# a_4653_n1142# avdd.t103 sky130_fd_pr__pfet_g5v0d10v5 ad=0.2142 pd=1.99 as=0.2142 ps=1.99 w=0.42 l=1
X235 comparator_1.vnn avss.t411 comparator_1.vt comparator_1.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=8
X236 avdd.t373 avdd.t371 avdd.t372 avdd.t230 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=8
X237 comparator_1.vnn avss.t412 comparator_1.vt comparator_1.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=8
X238 rstring_mux_0.vtop.t12 rstring_mux_0.ena_b avdd.t477 avdd.t476 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X239 sky130_fd_sc_hvl__inv_16_0.A sky130_fd_sc_hvl__inv_4_0.A avdd.t120 avdd.t119 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.4275 ps=3.57 w=1.5 l=0.5
X240 a_n3795_n1142# a_n3895_n1230# dvss.t371 dvss.t370 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X241 avdd.t84 comparator_1.vnn comparator_1.vnn avdd.t80 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X242 dcomp3v3uv comparator_0.n1 avss.t59 avss.t58 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X243 rstring_mux_0.vtrip5.t5 rstring_mux_0.vtrip_decoded_b_avdd[5] comparator_0.vinn.t45 avdd.t578 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X244 avdd.t96 ibias_gen_0.vp1.t11 ibias_gen_0.vp1.t12 avdd.t95 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X245 porb.t29 sky130_fd_sc_hd__inv_4_1.Y dvdd.t167 dvdd.t166 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X246 comparator_0.vinn.t7 rstring_mux_0.vtrip_decoded_avdd[3] rstring_mux_0.vtrip3.t2 avss.t75 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X247 rc_osc_0.m rc_osc_0.n.t7 dvdd.t175 dvdd.t174 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X248 rstring_mux_0.vtrip3.t7 rstring_mux_0.otrip_decoded_avdd[3] vin avss.t255 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X249 comparator_0.vinn.t27 rstring_mux_0.vtrip_decoded_b_avdd[7] rstring_mux_0.vtrip7.t9 avdd.t416 sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=0.6
X250 avdd.t648 comparator_1.vpp comparator_1.vpp avdd.t65 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X251 dvdd.t229 sky130_fd_sc_hd__inv_4_1.A sky130_fd_sc_hd__inv_4_1.Y dvdd.t228 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X252 avdd.t7 a_n3085_6745# a_n3778_7859# avdd.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=0.2142 pd=1.99 as=0.2142 ps=1.99 w=0.42 l=1
X253 dvss.t189 a_n6007_n1230# a_n5907_n1142# dvss.t188 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X254 dvss.t359 a_4553_n1230# a_4653_n1142# dvss.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X255 a_131_n11914# a_n247_n19314# avss.t97 sky130_fd_pr__res_xhigh_po_1p41 l=35
X256 avdd.t370 avdd.t369 avdd.t370 avdd.t240 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=8
X257 comparator_1.vn comparator_1.ena_b ibias_gen_0.ibias0 avdd.t446 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X258 avss.t121 ibias_gen_0.vn1.t11 ibias_gen_0.vp1.t1 avss.t120 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=8
X259 avdd.t124 a_7458_n2256# a_6765_n1142# avdd.t123 sky130_fd_pr__pfet_g5v0d10v5 ad=0.2142 pd=1.99 as=0.2142 ps=1.99 w=0.42 l=1
X260 rstring_mux_0.vtrip1.t1 rstring_mux_0.vtrip_decoded_avdd[1] comparator_0.vinn.t0 avss.t19 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X261 dvss.t80 sky130_fd_sc_hd__inv_4_0.Y pwup_filt.t11 dvss.t79 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X262 avdd.t612 comparator_0.vpp comparator_0.n0 avdd.t182 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X263 rc_osc_0.ena_b osc_ena.t1 dvdd.t137 dvdd.t136 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X264 comparator_0.vt avss.t413 comparator_0.vnn comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=8
X265 rstring_mux_0.vtrip0.t4 rstring_mux_0.otrip_decoded_avdd[0] vin avss.t313 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=0.6
X266 ibias_gen_0.vp1.t2 ibias_gen_0.vn1.t12 avss.t122 avss.t117 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=8
X267 rstring_mux_0.vtrip_decoded_avdd[6] a_7972_n3212# avdd.t509 avdd.t38 sky130_fd_pr__pfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.24375 ps=1.825 w=1.5 l=0.5
X268 comparator_0.vnn avss.t414 comparator_0.vt comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=8
X269 avss.t219 avss.t217 avss.t218 avss.t88 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=8
X270 ibias_gen_0.vp.t6 ibias_gen_0.isrc_sel ibias_gen_0.vp0.t5 avdd.t533 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X271 dvss.t756 sky130_fd_sc_hd__inv_4_3.Y dcomp.t14 dvss.t755 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X272 dvdd.t279 a_10873_n3956# sky130_fd_sc_hvl__lsbufhv2lv_1_1.X dvdd.t278 sky130_fd_pr__pfet_01v8_hvt ad=0.1568 pd=1.4 as=0.2968 ps=2.77 w=1.12 l=0.15
X273 dvdd.t263 sky130_fd_sc_hd__inv_4_4.Y por.t26 dvdd.t262 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X274 porb.t28 sky130_fd_sc_hd__inv_4_1.Y dvdd.t165 dvdd.t164 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X275 a_n5907_n1142# a_n6007_n1230# dvss.t187 dvss.t186 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X276 comparator_0.n1 comparator_0.n0 avss.t274 avss.t273 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.6
X277 comparator_1.vpp vin comparator_1.vt comparator_1.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X278 avss.t123 ibias_gen_0.vn1.t13 ibias_gen_0.vp1.t3 avss.t120 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=8
X279 comparator_0.vpp vbg_1v2.t6 comparator_0.vt comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X280 avss.t92 comparator_0.vm comparator_0.vm avss.t88 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X281 rstring_mux_0.vtrip4.t5 rstring_mux_0.otrip_decoded_avdd[4] vin avss.t76 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X282 dvdd.t113 dvss.t771 a_329_n1230# dvdd.t112 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X283 a_n10279_n22711# a_12321_n23089# dvss.t190 sky130_fd_pr__res_xhigh_po_1p41 l=111
X284 vin rstring_mux_0.otrip_decoded_avdd[2] rstring_mux_0.vtrip2.t5 avss.t339 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X285 a_n14999_9395# a_n14621_1995# avss.t103 sky130_fd_pr__res_xhigh_po_1p41 l=35
X286 dcomp3v3uv comparator_0.n1 avdd.t60 avdd.t59 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X287 comparator_0.vinn.t35 rstring_mux_0.vtrip_decoded_b_avdd[3] rstring_mux_0.vtrip3.t8 avdd.t444 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X288 avdd.t563 sky130_fd_sc_hvl__inv_16_0.A porb_h.t28 avdd.t562 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X289 dvdd.t239 vl sky130_fd_sc_hd__inv_4_3.Y dvdd.t238 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X290 avdd.t217 a_2541_n1142# a_3748_n1478# avdd.t107 sky130_fd_pr__pfet_g5v0d10v5 ad=0.24375 pd=1.825 as=0.3975 ps=3.53 w=1.5 l=0.5
X291 rstring_mux_0.vtrip0.t9 rstring_mux_0.vtrip_decoded_avdd[0] comparator_0.vinn.t41 avss.t375 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X292 rstring_mux_0.vtrip7.t4 rstring_mux_0.otrip_decoded_avdd[7] vin avss.t102 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X293 a_n10463_9395# a_n10085_1995# avss.t98 sky130_fd_pr__res_xhigh_po_1p41 l=35
X294 dvss.t624 a_n8119_n1230# a_n8019_n1142# dvss.t623 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X295 dvss.t587 a_6665_n1230# a_6765_n1142# dvss.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X296 avdd.t136 a_9570_n2256# a_8877_n1142# avdd.t135 sky130_fd_pr__pfet_g5v0d10v5 ad=0.2142 pd=1.99 as=0.2142 ps=1.99 w=0.42 l=1
X297 dvdd.t37 sky130_fd_sc_hd__inv_4_0.Y pwup_filt.t29 dvdd.t36 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X298 vin avdd.t367 vin avdd.t368 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=0.6
X299 dvss.t78 sky130_fd_sc_hd__inv_4_0.Y pwup_filt.t10 dvss.t77 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X300 dvss.t517 sky130_fd_sc_hd__inv_4_1.Y porb.t13 dvss.t516 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X301 comparator_0.vnn comparator_0.vnn avdd.t196 avdd.t186 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X302 comparator_0.vinn.t19 avss.t215 comparator_0.vinn.t19 avss.t216 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=0.6
X303 avdd.t83 comparator_1.vnn comparator_1.vnn avdd.t80 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X304 avdd.t342 avdd.t340 avdd.t342 avdd.t341 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=4
X305 dvss.t213 a_697_n2212# a_1122_n2256# dvss.t212 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X306 avdd.t366 avdd.t365 avdd.t366 avdd.t240 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=8
X307 a_8877_n1142# a_8777_n1230# dvss.t203 dvss.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X308 rc_osc_0.in dvss.t581 sky130_fd_pr__cap_mim_m3_2 l=30 w=30
X309 ibias_gen_0.vp.t0 avss.t213 ibias_gen_0.vp.t0 avss.t214 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=0.6
X310 comparator_1.vn comparator_1.vn avss.t294 avss.t284 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X311 dcomp.t28 sky130_fd_sc_hd__inv_4_3.Y dvdd.t306 dvdd.t305 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X312 dvss.t196 a_8877_n2876# a_10084_n3212# dvss.t195 sky130_fd_pr__nfet_g5v0d10v5 ad=0.121875 pd=1.075 as=0.19875 ps=2.03 w=0.75 l=0.5
X313 a_429_n1142# a_329_n1230# dvss.t422 dvss.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X314 rstring_mux_0.otrip_decoded_avdd[6] a_n476_n3212# avdd.t128 avdd.t127 sky130_fd_pr__pfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.24375 ps=1.825 w=1.5 l=0.5
X315 avdd.t364 avdd.t363 avdd.t364 avdd.t240 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=8
X316 porb_h.t12 sky130_fd_sc_hvl__inv_16_0.A avss.t367 avss.t366 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X317 a_n11975_9395# a_n12353_1995# avss.t104 sky130_fd_pr__res_xhigh_po_1p41 l=35
X318 avdd.t412 a_4653_n1142# a_5860_n1478# avdd.t207 sky130_fd_pr__pfet_g5v0d10v5 ad=0.24375 pd=1.825 as=0.3975 ps=3.53 w=1.5 l=0.5
X319 dvss.t202 a_8777_n1230# a_8877_n1142# dvss.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X320 comparator_0.vt comparator_0.vinn.t53 comparator_0.vnn comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X321 comparator_0.vinn.t23 rstring_mux_0.vtrip_decoded_avdd[5] rstring_mux_0.vtrip5.t4 avss.t248 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X322 avdd.t82 comparator_1.vnn comparator_1.vm avdd.t65 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X323 avdd.t490 ibias_gen_0.isrc_sel_b ibias_gen_0.vp0.t2 avdd.t489 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X324 schmitt_trigger_0.m.t11 schmitt_trigger_0.in.t2 dvdd.t91 dvdd.t90 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X325 dvss.t515 sky130_fd_sc_hd__inv_4_1.Y porb.t12 dvss.t514 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X326 avdd.t362 avdd.t361 avdd.t362 avdd.t234 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=8
X327 rstring_mux_0.otrip_decoded_b_avdd[0] rstring_mux_0.otrip_decoded_avdd[0] avss.t312 avss.t311 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X328 vin avdd.t359 vin avdd.t360 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=0.6
X329 comparator_1.vnn avss.t415 comparator_1.vt comparator_1.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=8
X330 rstring_mux_0.otrip_decoded_b_avdd[4] rstring_mux_0.otrip_decoded_avdd[4] avdd.t112 avdd.t111 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X331 avdd.t358 avdd.t356 avdd.t357 avdd.t230 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=8
X332 dvss.t674 sky130_fd_sc_hd__inv_4_4.Y por.t12 dvss.t673 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X333 a_9203_n11914# a_9581_n19314# avss.t106 sky130_fd_pr__res_xhigh_po_1p41 l=35
X334 avss.t365 sky130_fd_sc_hvl__inv_16_0.A porb_h.t11 avss.t364 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X335 dvss.t421 a_329_n1230# a_429_n1142# dvss.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X336 rc_osc_0.m rc_osc_0.in dvdd.t217 dvdd.t216 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X337 rc_osc_0.m rc_osc_0.in dvss.t580 dvss.t579 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.1475 ps=1.295 w=1 l=0.5
X338 rstring_mux_0.vtrip5.t8 rstring_mux_0.otrip_decoded_avdd[5] vin avss.t398 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X339 avdd.t401 ibias_gen_0.vp0.t6 ibias_gen_0.vp0.t7 avdd.t400 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X340 a_8877_n1142# a_8777_n1230# dvss.t201 dvss.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X341 a_n7751_n2212# a_n8119_n1230# dvdd.t233 dvdd.t232 sky130_fd_pr__pfet_01v8_hvt ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X342 comparator_0.vinn.t11 rstring_mux_0.vtrip_decoded_b_avdd[2] rstring_mux_0.vtrip2.t2 avdd.t138 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X343 avdd.t81 comparator_1.vnn comparator_1.vnn avdd.t80 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X344 rc_osc_0.n.t2 rc_osc_0.m dvdd.t47 dvdd.t46 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X345 a_n6673_n11914# a_n6295_n19314# avss.t105 sky130_fd_pr__res_xhigh_po_1p41 l=35
X346 comparator_0.vt comparator_0.vinn.t54 comparator_0.vnn comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X347 avdd.t79 comparator_1.vnn comparator_1.vpp avdd.t65 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X348 ibias_gen_0.vn0.t16 vbg_1v2.t7 ibias_gen_0.vstart.t8 avss.t128 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X349 a_5346_n2256# a_4921_n2212# dvss.t223 dvss.t222 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X350 avdd.t355 avdd.t353 avdd.t354 avdd.t230 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=8
X351 comparator_1.vpp comparator_1.vnn avdd.t78 avdd.t63 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X352 avdd.t532 ibias_gen_0.isrc_sel a_n16775_n2223# avdd.t531 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X353 rstring_mux_0.vtrip2.t4 rstring_mux_0.otrip_decoded_avdd[2] vin avss.t338 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X354 dvss.t513 sky130_fd_sc_hd__inv_4_1.Y porb.t11 dvss.t512 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X355 comparator_1.vm comparator_1.ena_b avss.t291 avss.t290 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X356 dvdd.t227 sky130_fd_sc_hd__inv_4_1.A sky130_fd_sc_hd__inv_4_1.Y dvdd.t226 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X357 dcomp3v3 comparator_1.n1 avss.t36 avss.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X358 dvss.t672 sky130_fd_sc_hd__inv_4_4.Y por.t11 dvss.t671 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X359 avdd.t522 rstring_mux_0.ena ibias_gen_0.vp1.t15 avdd.t521 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X360 avdd.t352 avdd.t351 avdd.t352 avdd.t234 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=8
X361 porb_h.t27 sky130_fd_sc_hvl__inv_16_0.A avdd.t561 avdd.t560 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X362 ibias_gen_0.vp1.t17 ibias_gen_0.isrc_sel avdd.t530 avdd.t529 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=2
X363 dcomp.t13 sky130_fd_sc_hd__inv_4_3.Y dvss.t754 dvss.t753 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X364 rstring_mux_0.ena a_10084_n3212# dvss.t194 dvss.t193 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.121875 ps=1.075 w=0.75 l=0.5
X365 rstring_mux_0.vtrip6.t5 rstring_mux_0.otrip_decoded_b_avdd[6] vin avdd.t450 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X366 comparator_1.vpp vin comparator_1.vt comparator_1.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X367 a_7458_n2256# a_7033_n2212# dvss.t235 dvss.t234 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X368 avdd.t146 a_n1683_n2876# a_n476_n3212# avdd.t127 sky130_fd_pr__pfet_g5v0d10v5 ad=0.24375 pd=1.825 as=0.3975 ps=3.53 w=1.5 l=0.5
X369 rstring_mux_0.vtrip5.t0 rstring_mux_0.vtrip4.t7 avss.t113 sky130_fd_pr__res_xhigh_po_1p41 l=35
X370 comparator_1.vpp vin comparator_1.vt comparator_1.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X371 comparator_0.vinn.t18 avss.t211 comparator_0.vinn.t18 avss.t212 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=0.6
X372 sky130_fd_sc_hd__inv_4_3.Y vl dvss.t637 dvss.t636 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X373 porb.t27 sky130_fd_sc_hd__inv_4_1.Y dvdd.t163 dvdd.t162 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X374 avdd.t143 a_n990_n3990# a_n1683_n2876# avdd.t142 sky130_fd_pr__pfet_g5v0d10v5 ad=0.2142 pd=1.99 as=0.2142 ps=1.99 w=0.42 l=1
X375 dvdd.t304 sky130_fd_sc_hd__inv_4_3.Y dcomp.t27 dvdd.t303 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X376 pwup_filt.t28 sky130_fd_sc_hd__inv_4_0.Y dvdd.t35 dvdd.t34 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X377 a_n1683_n2876# a_n1783_n2964# dvss.t353 dvss.t352 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X378 dvss.t310 dvss.t308 a_2441_n2964# dvss.t309 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X379 comparator_0.vn comparator_0.ena_b comparator_0.ibias avdd.t141 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X380 rc_osc_0.in dvss.t578 sky130_fd_pr__cap_mim_m3_2 l=30 w=30
X381 a_n9697_n11914# a_n10075_n19314# avss.t107 sky130_fd_pr__res_xhigh_po_1p41 l=35
X382 avss.t57 comparator_0.n1 dcomp3v3uv avss.t56 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X383 avdd.t350 avdd.t349 avdd.t350 avdd.t240 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=8
X384 comparator_0.vinn.t17 avss.t209 comparator_0.vinn.t17 avss.t210 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=0.6
X385 comparator_1.vnn comparator_1.vnn avdd.t77 avdd.t73 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X386 dvss.t670 sky130_fd_sc_hd__inv_4_4.Y por.t10 dvss.t669 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X387 comparator_1.vnn rstring_mux_0.ena avdd.t520 avdd.t519 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X388 dcomp3v3 comparator_1.n1 avdd.t29 avdd.t28 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X389 dvss.t76 sky130_fd_sc_hd__inv_4_0.Y pwup_filt.t9 dvss.t75 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X390 a_2541_n1142# a_2441_n1230# dvss.t51 dvss.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X391 a_n990_n2256# a_n1415_n2212# dvss.t246 dvss.t245 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X392 dvdd.t315 dvdd.t313 dvdd.t315 dvdd.t314 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.18
X393 a_n13477_n11914# a_n13099_n19314# avss.t114 sky130_fd_pr__res_xhigh_po_1p41 l=35
X394 dcomp.t12 sky130_fd_sc_hd__inv_4_3.Y dvss.t752 dvss.t751 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X395 sky130_fd_sc_hd__inv_4_0.Y schmitt_trigger_0.out.t6 dvdd.t57 dvdd.t56 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X396 a_n3795_n1142# a_n3895_n1230# dvss.t369 dvss.t368 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X397 dvss.t638 a_n1683_n1142# a_n476_n1478# dvss.t175 sky130_fd_pr__nfet_g5v0d10v5 ad=0.121875 pd=1.075 as=0.19875 ps=2.03 w=0.75 l=0.5
X398 avdd.t152 a_n5214_n2256# a_n5907_n1142# avdd.t151 sky130_fd_pr__pfet_g5v0d10v5 ad=0.2142 pd=1.99 as=0.2142 ps=1.99 w=0.42 l=1
X399 rstring_mux_0.vtrip1.t6 rstring_mux_0.otrip_decoded_b_avdd[1] vin avdd.t413 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X400 comparator_0.vinn.t16 avss.t207 comparator_0.vinn.t16 avss.t208 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=0.6
X401 comparator_0.vn comparator_0.ena_b avss.t112 avss.t111 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X402 porb_h.t10 sky130_fd_sc_hvl__inv_16_0.A avss.t363 avss.t362 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X403 ibias_gen_0.vp.t1 avdd.t347 ibias_gen_0.vp.t1 avdd.t348 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=0.6
X404 a_n10279_n24223# a_12321_n23845# dvss.t249 sky130_fd_pr__res_xhigh_po_1p41 l=111
X405 avdd.t118 sky130_fd_sc_hvl__inv_4_0.A sky130_fd_sc_hvl__inv_16_0.A avdd.t117 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X406 porb.t26 sky130_fd_sc_hd__inv_4_1.Y dvdd.t161 dvdd.t160 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X407 dvss.t760 a_n8019_n1142# a_n6812_n1478# dvss.t759 sky130_fd_pr__nfet_g5v0d10v5 ad=0.121875 pd=1.075 as=0.19875 ps=2.03 w=0.75 l=0.5
X408 dvss.t50 a_2441_n1230# a_2541_n1142# dvss.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X409 rstring_mux_0.otrip_decoded_b_avdd[5] rstring_mux_0.otrip_decoded_avdd[5] avss.t397 avss.t396 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X410 dcomp3v3uv comparator_0.n1 avss.t55 avss.t54 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X411 avdd.t346 avdd.t345 avdd.t346 avdd.t234 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=8
X412 pwup_filt.t27 sky130_fd_sc_hd__inv_4_0.Y dvdd.t33 dvdd.t32 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X413 a_n3795_n2876# a_n3895_n2964# dvss.t414 dvss.t413 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X414 a_2541_n2876# a_2441_n2964# dvss.t434 dvss.t433 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X415 comparator_0.vt comparator_0.vinn.t55 comparator_0.vnn comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X416 a_n26074_n2937# a_n26452_n10337# avss.t0 sky130_fd_pr__res_xhigh_po_1p41 l=35
X417 a_n23050_n2937# a_n23428_n10337# avss.t0 sky130_fd_pr__res_xhigh_po_1p41 l=35
X418 dvss.t258 a_10515_n2156# a_10874_n2222# dvss.t257 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.19875 ps=2.03 w=0.75 l=0.5
X419 a_n5161_n11914# a_n4783_n19314# avss.t116 sky130_fd_pr__res_xhigh_po_1p41 l=35
X420 a_n5907_n1142# a_n6007_n1230# dvss.t185 dvss.t184 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X421 rstring_mux_0.vtrip_decoded_avdd[3] a_3748_n1478# dvss.t177 dvss.t175 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.121875 ps=1.075 w=0.75 l=0.5
X422 comparator_0.vnn avss.t416 avdd.t170 avdd.t169 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X423 a_n5907_n1142# a_n6007_n1230# dvss.t183 dvss.t182 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X424 a_4653_n1142# a_4553_n1230# dvss.t358 dvss.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X425 avdd.t160 a_n7326_n2256# a_n8019_n1142# avdd.t159 sky130_fd_pr__pfet_g5v0d10v5 ad=0.2142 pd=1.99 as=0.2142 ps=1.99 w=0.42 l=1
X426 a_n5161_n11914# a_n5539_n19314# avss.t115 sky130_fd_pr__res_xhigh_po_1p41 l=35
X427 avdd.t647 comparator_1.vpp comparator_1.vnn avdd.t80 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X428 comparator_1.vnn comparator_1.vnn avdd.t76 avdd.t73 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X429 a_n25318_n2937# a_n25696_n10337# avss.t0 sky130_fd_pr__res_xhigh_po_1p41 l=35
X430 ibias_gen_0.vn1.t3 ibias_gen_0.vn1.t2 avss.t118 avss.t117 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=8
X431 dvss.t124 a_10515_n1026# a_10515_n2156# dvss.t123 sky130_fd_pr__nfet_g5v0d10v5 ad=0.178875 pd=1.26 as=0.1197 ps=1.41 w=0.42 l=0.5
X432 a_n1415_n2212# a_n1783_n1230# dvss.t609 dvss.t608 sky130_fd_pr__nfet_01v8 ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X433 dvss.t622 a_n8119_n1230# a_n8019_n1142# dvss.t621 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X434 a_4653_n2876# a_4553_n2964# dvss.t278 dvss.t277 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X435 dvss.t726 a_10873_n3956# sky130_fd_sc_hvl__lsbufhv2lv_1_1.X dvss.t725 sky130_fd_pr__nfet_01v8 ad=0.1961 pd=2.01 as=0.1961 ps=2.01 w=0.74 l=0.15
X436 rc_osc_0.in dvss.t577 sky130_fd_pr__cap_mim_m3_2 l=30 w=30
X437 avss.t34 comparator_1.n1 dcomp3v3 avss.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X438 a_10873_n3956# a_10514_n3890# dvss.t266 dvss.t265 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.178875 ps=1.26 w=0.75 l=0.5
X439 a_n8019_n1142# a_n8119_n1230# dvss.t620 dvss.t619 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X440 a_6765_n1142# a_6665_n1230# dvss.t586 dvss.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X441 dvss.t402 isrc_sel.t0 a_8777_n1230# dvss.t401 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X442 rstring_mux_0.vtrip2.t9 rstring_mux_0.otrip_decoded_b_avdd[2] vin avdd.t628 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X443 avdd.t344 avdd.t343 avdd.t344 avdd.t234 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=8
X444 a_n14999_9395# vl avss.t65 sky130_fd_pr__res_xhigh_po_1p41 l=35
X445 dvss.t511 sky130_fd_sc_hd__inv_4_1.Y porb.t10 dvss.t510 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X446 a_n8019_n1142# a_n8119_n1230# dvss.t618 dvss.t617 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X447 dvss.t307 dvss.t305 a_329_n2964# dvss.t306 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X448 rstring_mux_0.vtrip_decoded_b_avdd[6] rstring_mux_0.vtrip_decoded_avdd[6] avdd.t122 avdd.t121 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X449 rstring_mux_0.otrip_decoded_b_avdd[7] rstring_mux_0.otrip_decoded_avdd[7] avss.t101 avss.t100 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X450 avdd.t164 a_n3778_7859# a_n2571_7523# avdd.t163 sky130_fd_pr__pfet_g5v0d10v5 ad=0.24375 pd=1.825 as=0.3975 ps=3.53 w=1.5 l=0.5
X451 dvss.t668 sky130_fd_sc_hd__inv_4_4.Y por.t9 dvss.t667 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X452 avdd.t611 comparator_0.vpp comparator_0.vnn avdd.t182 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X453 a_n3527_n2212# a_n3895_n1230# dvss.t367 dvss.t366 sky130_fd_pr__nfet_01v8 ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X454 rstring_mux_0.otrip_decoded_avdd[4] a_n2588_n3212# avdd.t659 avdd.t155 sky130_fd_pr__pfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.24375 ps=1.825 w=1.5 l=0.5
X455 comparator_1.vnn avss.t417 comparator_1.vt comparator_1.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=8
X456 a_429_n1142# a_329_n1230# dvss.t420 dvss.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X457 a_10873_n2760# a_10514_n2760# dvss.t567 dvss.t565 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.178875 ps=1.26 w=0.75 l=0.5
X458 dcomp.t11 sky130_fd_sc_hd__inv_4_3.Y dvss.t750 dvss.t749 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X459 comparator_0.vinn.t15 avss.t205 comparator_0.vinn.t15 avss.t206 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=0.6
X460 rstring_mux_0.vtrip2.t1 rstring_mux_0.vtrip_decoded_b_avdd[2] comparator_0.vinn.t10 avdd.t137 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X461 sky130_fd_sc_hd__inv_4_1.A por_unbuf.t2 dvdd.t191 dvdd.t190 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X462 a_3911_n11914# a_4289_n19314# avss.t261 sky130_fd_pr__res_xhigh_po_1p41 l=35
X463 a_n10463_9395# a_n10841_1995# avss.t3 sky130_fd_pr__res_xhigh_po_1p41 l=35
X464 a_n3085_6745# a_n3510_6789# dvss.t454 dvss.t453 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X465 ibias_gen_0.vp1.t4 ibias_gen_0.vn1.t14 avss.t124 avss.t117 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=8
X466 a_n8941_n11914# a_n8563_n19314# avss.t263 sky130_fd_pr__res_xhigh_po_1p41 l=35
X467 a_n11965_n11914# a_n11587_n19314# avss.t14 sky130_fd_pr__res_xhigh_po_1p41 l=35
X468 a_6765_n2876# a_6665_n2964# dvss.t397 dvss.t396 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X469 rstring_mux_0.vtrip_decoded_b_avdd[6] rstring_mux_0.vtrip_decoded_avdd[6] avss.t96 avss.t95 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X470 comparator_0.vt vbg_1v2.t8 comparator_0.vpp comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X471 comparator_0.ena_b avss.t418 avdd.t168 avdd.t167 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X472 ibias_gen_0.vp0.t1 avdd.t337 avdd.t339 avdd.t338 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X473 avss.t204 avss.t202 avss.t203 avss.t193 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=8
X474 comparator_1.vnn vbg_1v2.t9 comparator_1.vt comparator_1.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X475 porb.t25 sky130_fd_sc_hd__inv_4_1.Y dvdd.t159 dvdd.t158 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X476 dvss.t334 a_2809_n2212# a_3234_n2256# dvss.t333 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X477 avdd.t336 avdd.t334 avdd.t335 avdd.t221 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=8
X478 comparator_1.vnn comparator_1.vnn avdd.t75 avdd.t73 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X479 sky130_fd_sc_hd__inv_4_3.Y vl dvss.t635 dvss.t634 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X480 dvss.t419 a_329_n1230# a_429_n1142# dvss.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X481 dvdd.t87 a_10874_n2222# vl dvdd.t66 sky130_fd_pr__pfet_01v8_hvt ad=0.1568 pd=1.4 as=0.2968 ps=2.77 w=1.12 l=0.15
X482 avdd.t646 comparator_1.vpp comparator_1.vnn avdd.t80 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X483 comparator_1.vnn vbg_1v2.t10 comparator_1.vt comparator_1.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X484 avss.t201 avss.t200 ibias_gen_0.vr.t0 avss.t67 sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=4
X485 dvdd.t302 sky130_fd_sc_hd__inv_4_3.Y dcomp.t26 dvdd.t301 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X486 pwup_filt.t26 sky130_fd_sc_hd__inv_4_0.Y dvdd.t31 dvdd.t30 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X487 avss.t53 comparator_0.n1 dcomp3v3uv avss.t52 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.6
X488 dvdd.t261 sky130_fd_sc_hd__inv_4_4.Y por.t25 dvdd.t260 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X489 avdd.t214 a_8877_n1142# a_10084_n1478# avdd.t213 sky130_fd_pr__pfet_g5v0d10v5 ad=0.24375 pd=1.825 as=0.3975 ps=3.53 w=1.5 l=0.5
X490 avdd.t195 comparator_0.vnn comparator_0.vpp avdd.t179 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X491 dvss.t452 a_n3510_6789# a_n3085_6745# dvss.t451 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X492 dvss.t666 sky130_fd_sc_hd__inv_4_4.Y por.t8 dvss.t665 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X493 a_n5639_n2212# a_n6007_n1230# dvss.t181 dvss.t180 sky130_fd_pr__nfet_01v8 ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X494 comparator_0.vpp comparator_0.vpp avdd.t610 avdd.t177 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X495 comparator_0.vinn.t32 avdd.t332 comparator_0.vinn.t32 avdd.t333 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=0.6
X496 a_n9707_9395# a_n9329_1995# avss.t10 sky130_fd_pr__res_xhigh_po_1p41 l=35
X497 rstring_mux_0.otrip_decoded_b_avdd[2] rstring_mux_0.otrip_decoded_avdd[2] avdd.t537 avdd.t536 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X498 comparator_0.vt vbg_1v2.t11 comparator_0.vpp comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X499 comparator_1.vt vbg_1v2.t12 comparator_1.vnn comparator_1.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X500 sky130_fd_sc_hd__inv_4_0.Y schmitt_trigger_0.out.t7 dvdd.t59 dvdd.t58 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X501 avdd.t609 comparator_0.vpp comparator_0.vnn avdd.t182 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X502 dvdd.t95 schmitt_trigger_0.m.t14 schmitt_trigger_0.out.t3 dvdd.t94 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X503 rstring_mux_0.vtop.t11 rstring_mux_0.ena_b avdd.t475 avdd.t474 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=0.6
X504 porb.t24 sky130_fd_sc_hd__inv_4_1.Y dvdd.t157 dvdd.t156 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X505 a_n7751_n3946# a_n8119_n2964# dvss.t708 dvss.t707 sky130_fd_pr__nfet_01v8 ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X506 a_9570_n2256# a_9145_n2212# dvss.t33 dvss.t32 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X507 dvdd.t300 sky130_fd_sc_hd__inv_4_3.Y dcomp.t25 dvdd.t299 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X508 porb_h.t26 sky130_fd_sc_hvl__inv_16_0.A avdd.t559 avdd.t558 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X509 dvss.t256 a_10515_n2156# a_10874_n2222# dvss.t255 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.19875 ps=2.03 w=0.75 l=0.5
X510 a_n14989_n11914# a_n15367_n19314# avss.t8 sky130_fd_pr__res_xhigh_po_1p41 l=35
X511 comparator_1.vnn comparator_1.vnn avdd.t74 avdd.t73 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X512 comparator_1.n0 comparator_1.ena_b avss.t289 avss.t288 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X513 sky130_fd_sc_hvl__inv_4_0.A sky130_fd_sc_hvl__inv_1_0.A avss.t389 avss.t388 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X514 avdd.t331 avdd.t329 avdd.t331 avdd.t330 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=4
X515 avdd.t156 a_n3795_n2876# a_n2588_n3212# avdd.t155 sky130_fd_pr__pfet_g5v0d10v5 ad=0.24375 pd=1.825 as=0.3975 ps=3.53 w=1.5 l=0.5
X516 a_7458_n2256# a_7033_n2212# dvss.t233 dvss.t232 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X517 a_10514_n3890# a_10514_n2760# avdd.t447 avdd.t45 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.1197 ps=1.41 w=0.42 l=0.5
X518 a_7691_n11914# a_8069_n19314# avss.t407 sky130_fd_pr__res_xhigh_po_1p41 l=35
X519 dcomp3v3 comparator_1.n1 avss.t32 avss.t31 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X520 a_n10279_n24979# a_12321_n25357# dvss.t765 sky130_fd_pr__res_xhigh_po_1p41 l=111
X521 a_n15745_n11914# a_n15367_n19314# avss.t277 sky130_fd_pr__res_xhigh_po_1p41 l=35
X522 dvss.t607 a_n1783_n1230# a_n1683_n1142# dvss.t606 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X523 dvss.t415 a_4653_n1142# a_5860_n1478# dvss.t175 sky130_fd_pr__nfet_g5v0d10v5 ad=0.121875 pd=1.075 as=0.19875 ps=2.03 w=0.75 l=0.5
X524 avdd.t174 a_n3102_n3990# a_n3795_n2876# avdd.t173 sky130_fd_pr__pfet_g5v0d10v5 ad=0.2142 pd=1.99 as=0.2142 ps=1.99 w=0.42 l=1
X525 a_n3510_6789# a_n3878_7771# dvdd.t173 dvdd.t172 sky130_fd_pr__pfet_01v8_hvt ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X526 rstring_mux_0.vtrip7.t8 rstring_mux_0.vtrip_decoded_b_avdd[7] comparator_0.vinn.t26 avdd.t415 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X527 avdd.t512 a_n1683_n1142# a_n990_n2256# avdd.t511 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.1365 ps=1.49 w=0.42 l=1
X528 avdd.t328 avdd.t326 avdd.t327 avdd.t221 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=8
X529 a_n1683_n2876# a_n1783_n2964# dvss.t351 dvss.t350 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X530 sky130_fd_sc_hvl__inv_16_0.A sky130_fd_sc_hvl__inv_4_0.A avdd.t116 avdd.t115 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X531 ibias_gen_0.ena_b rstring_mux_0.ena avdd.t518 avdd.t517 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=1
X532 a_n3102_n2256# a_n3527_n2212# dvss.t11 dvss.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X533 avdd.t194 comparator_0.vnn comparator_0.vpp avdd.t179 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X534 avdd.t325 avdd.t324 avdd.t325 avdd.t234 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=8
X535 comparator_1.vm comparator_1.vnn avdd.t72 avdd.t63 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X536 avss.t199 avss.t198 avss.t199 avss.t136 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=8
X537 dvdd.t298 sky130_fd_sc_hd__inv_4_3.Y dcomp.t24 dvdd.t297 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X538 a_2541_n1142# a_2441_n1230# dvss.t49 dvss.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X539 ibias_gen_0.isrc_sel a_10084_n1478# avdd.t210 avdd.t209 sky130_fd_pr__pfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.24375 ps=1.825 w=1.5 l=0.5
X540 dvss.t304 dvss.t302 a_4553_n1230# dvss.t303 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X541 comparator_0.vpp comparator_0.vpp avdd.t608 avdd.t177 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X542 a_2399_n11914# a_2777_n19314# avss.t66 sky130_fd_pr__res_xhigh_po_1p41 l=35
X543 a_10515_n1026# dcomp3v3 avdd.t43 avdd.t42 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.1197 ps=1.41 w=0.42 l=0.5
X544 avdd.t3 a_n5907_n2876# a_n4700_n3212# avdd.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0.24375 pd=1.825 as=0.3975 ps=3.53 w=1.5 l=0.5
X545 comparator_0.vt comparator_0.vinn.t56 comparator_0.vnn comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X546 porb_h.t9 sky130_fd_sc_hvl__inv_16_0.A avss.t361 avss.t360 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X547 ibias_gen_0.vn0.t15 vbg_1v2.t13 ibias_gen_0.vstart.t7 avss.t128 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X548 schmitt_trigger_0.out.t2 schmitt_trigger_0.m.t15 dvdd.t97 dvdd.t96 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X549 a_9570_n2256# a_9145_n2212# dvss.t31 dvss.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X550 a_3155_n11914# a_2777_n19314# avss.t258 sky130_fd_pr__res_xhigh_po_1p41 l=35
X551 a_n10453_n11914# a_n10831_n19314# avss.t64 sky130_fd_pr__res_xhigh_po_1p41 l=35
X552 rstring_mux_0.vtrip_decoded_avdd[5] a_5860_n1478# dvss.t339 dvss.t175 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.121875 ps=1.075 w=0.75 l=0.5
X553 dvss.t9 a_n3527_n2212# a_n3102_n2256# dvss.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X554 dvss.t244 a_n1415_n2212# a_n990_n2256# dvss.t243 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X555 a_4921_n2212# a_4553_n1230# dvss.t357 dvss.t356 sky130_fd_pr__nfet_01v8 ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X556 avdd.t114 sky130_fd_sc_hvl__inv_4_0.A sky130_fd_sc_hvl__inv_16_0.A avdd.t113 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.21 ps=1.78 w=1.5 l=0.5
X557 comparator_1.vnn avss.t419 comparator_1.vt comparator_1.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=8
X558 dvss.t365 a_n3895_n1230# a_n3795_n1142# dvss.t364 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X559 rstring_mux_0.vtop.t10 rstring_mux_0.ena_b avdd.t473 avdd.t472 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X560 a_n3795_n2876# a_n3895_n2964# dvss.t412 dvss.t411 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X561 avss.t359 sky130_fd_sc_hvl__inv_16_0.A porb_h.t8 avss.t358 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X562 sky130_fd_sc_hd__inv_4_1.A por_unbuf.t3 dvdd.t193 dvdd.t192 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X563 a_n5214_n2256# a_n5639_n2212# dvss.t44 dvss.t43 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X564 rstring_mux_0.vtrip_decoded_avdd[4] a_5860_n3212# avdd.t453 avdd.t452 sky130_fd_pr__pfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.24375 ps=1.825 w=1.5 l=0.5
X565 comparator_0.vt avss.t420 comparator_0.vnn comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=8
X566 dvss.t301 dvss.t299 a_6665_n1230# dvss.t300 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X567 a_131_n11914# a_509_n19314# avss.t13 sky130_fd_pr__res_xhigh_po_1p41 l=35
X568 rc_osc_0.in dvss.t576 sky130_fd_pr__cap_mim_m3_2 l=30 w=30
X569 comparator_0.vt vbg_1v2.t14 comparator_0.vpp comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X570 avdd.t645 comparator_1.vpp comparator_1.vnn avdd.t80 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X571 comparator_1.vnn vbg_1v2.t15 comparator_1.vt comparator_1.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X572 a_n3778_7859# a_n3878_7771# dvss.t529 dvss.t528 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X573 a_4653_n1142# a_4553_n1230# dvss.t355 dvss.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X574 a_n990_n2256# a_n1415_n2212# dvss.t242 dvss.t241 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X575 a_n1415_n2212# a_n1783_n1230# dvdd.t231 dvdd.t230 sky130_fd_pr__pfet_01v8_hvt ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X576 dvss.t385 a_n6007_n2964# a_n5907_n2876# dvss.t384 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X577 dvss.t276 a_4553_n2964# a_4653_n2876# dvss.t275 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X578 por.t24 sky130_fd_sc_hd__inv_4_4.Y dvdd.t259 dvdd.t258 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X579 dcomp.t10 sky130_fd_sc_hd__inv_4_3.Y dvss.t748 dvss.t747 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X580 avdd.t658 a_n8019_n2876# a_n6812_n3212# avdd.t498 sky130_fd_pr__pfet_g5v0d10v5 ad=0.24375 pd=1.825 as=0.3975 ps=3.53 w=1.5 l=0.5
X581 ibias_gen_0.vp1.t16 ibias_gen_0.isrc_sel ibias_gen_0.vp.t5 avss.t337 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X582 schmitt_trigger_0.m.t6 schmitt_trigger_0.in.t3 dvss.t166 dvss.t165 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X583 avdd.t323 avdd.t321 avdd.t322 avdd.t221 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=8
X584 comparator_0.vpp comparator_0.vpp avdd.t607 avdd.t177 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X585 comparator_1.vt avss.t421 comparator_1.vnn comparator_1.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=8
X586 ibias_gen_0.vstart.t6 vbg_1v2.t16 ibias_gen_0.vn0.t14 avss.t128 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X587 dvss.t298 dvss.t296 schmitt_trigger_0.m.t4 dvss.t297 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X588 dvss.t585 a_6665_n1230# a_6765_n1142# dvss.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X589 rstring_mux_0.vtrip_decoded_avdd[7] a_7972_n1478# dvss.t176 dvss.t175 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.121875 ps=1.075 w=0.75 l=0.5
X590 dvss.t42 a_n5639_n2212# a_n5214_n2256# dvss.t41 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X591 dvss.t575 rc_osc_0.in rc_osc_0.m dvss.t574 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X592 rstring_mux_0.vtop.t9 rstring_mux_0.ena_b avdd.t471 avdd.t470 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X593 avdd.t644 comparator_1.vpp comparator_1.vnn avdd.t80 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X594 comparator_1.vt vbg_1v2.t17 comparator_1.vnn comparator_1.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X595 dvss.t664 sky130_fd_sc_hd__inv_4_4.Y por.t7 dvss.t663 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X596 dvdd.t215 rc_osc_0.in rc_osc_0.m dvdd.t214 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X597 rc_osc_0.in dvss.t573 sky130_fd_pr__cap_mim_m3_2 l=30 w=30
X598 comparator_0.vt avss.t422 comparator_0.vnn comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=8
X599 comparator_1.vt avss.t423 comparator_1.vnn comparator_1.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=8
X600 dvss.t527 a_n3878_7771# a_n3778_7859# dvss.t526 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X601 comparator_0.vnn avss.t424 comparator_0.vt comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=8
X602 avss.t91 comparator_0.vm comparator_0.n0 avss.t88 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X603 avdd.t193 comparator_0.vnn comparator_0.vpp avdd.t179 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X604 avdd.t320 avdd.t319 avdd.t320 avdd.t234 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=8
X605 comparator_1.vt vbg_1v2.t18 comparator_1.vnn comparator_1.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X606 sky130_fd_sc_hd__inv_4_4.Y por_unbuf.t4 dvdd.t195 dvdd.t194 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X607 a_n5907_n2876# a_n6007_n2964# dvss.t383 dvss.t382 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X608 dvdd.t111 dvss.t772 a_2441_n2964# dvdd.t110 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X609 comparator_0.vnn comparator_0.vinn.t57 comparator_0.vt comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X610 ibias_gen_0.isrc_sel_b avdd.t317 ibias_gen_0.ena_b avdd.t318 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X611 pwup_filt.t25 sky130_fd_sc_hd__inv_4_0.Y dvdd.t29 dvdd.t28 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X612 dvdd.t117 isrc_sel.t1 a_8777_n1230# dvdd.t116 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X613 dvdd.t45 rc_osc_0.m rc_osc_0.n.t1 dvdd.t44 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X614 comparator_0.vn comparator_0.vn avss.t392 avss.t109 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X615 a_n7326_n2256# a_n7751_n2212# dvss.t466 dvss.t465 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X616 a_6179_n11914# a_6557_n19314# avss.t241 sky130_fd_pr__res_xhigh_po_1p41 l=35
X617 a_n14233_n11914# a_n13855_n19314# avss.t70 sky130_fd_pr__res_xhigh_po_1p41 l=35
X618 comparator_0.vpp vbg_1v2.t19 comparator_0.vt comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X619 avdd.t397 a_429_n2876# a_1636_n3212# avdd.t396 sky130_fd_pr__pfet_g5v0d10v5 ad=0.24375 pd=1.825 as=0.3975 ps=3.53 w=1.5 l=0.5
X620 dvss.t264 a_10514_n3890# a_10873_n3956# dvss.t263 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.19875 ps=2.03 w=0.75 l=0.5
X621 comparator_0.vinn.t40 rstring_mux_0.vtrip_decoded_b_avdd[0] rstring_mux_0.vtrip0.t7 avdd.t508 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X622 a_n23050_n2937# a_n22672_n10337# avss.t0 sky130_fd_pr__res_xhigh_po_1p41 l=35
X623 a_6765_n1142# a_6665_n1230# dvss.t584 dvss.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X624 a_n3527_n2212# a_n3895_n1230# dvdd.t123 dvdd.t122 sky130_fd_pr__pfet_01v8_hvt ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X625 comparator_1.vnn comparator_1.vpp avdd.t643 avdd.t73 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X626 dvss.t74 sky130_fd_sc_hd__inv_4_0.Y pwup_filt.t8 dvss.t73 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X627 dvss.t706 a_n8119_n2964# a_n8019_n2876# dvss.t705 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X628 dvss.t395 a_6665_n2964# a_6765_n2876# dvss.t394 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X629 a_n14233_n11914# a_n14611_n19314# avss.t264 sky130_fd_pr__res_xhigh_po_1p41 l=35
X630 a_n13487_9395# a_n13865_1995# avss.t6 sky130_fd_pr__res_xhigh_po_1p41 l=35
X631 por.t23 sky130_fd_sc_hd__inv_4_4.Y dvdd.t257 dvdd.t256 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X632 avdd.t316 avdd.t314 avdd.t315 avdd.t230 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=8
X633 dvdd.t296 sky130_fd_sc_hd__inv_4_3.Y dcomp.t23 dvdd.t295 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X634 a_1122_n2256# a_697_n2212# dvss.t211 dvss.t210 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X635 a_n22294_n2937# a_n21916_n10337# avss.t0 sky130_fd_pr__res_xhigh_po_1p41 l=35
X636 schmitt_trigger_0.m.t10 schmitt_trigger_0.in.t4 dvdd.t73 dvdd.t72 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X637 dvss.t200 a_8777_n1230# a_8877_n1142# dvss.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X638 dvss.t464 a_n7751_n2212# a_n7326_n2256# dvss.t463 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X639 dvss.t489 a_697_n3946# a_1122_n3990# dvss.t488 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X640 rstring_mux_0.vtrip4.t4 rstring_mux_0.otrip_decoded_b_avdd[4] vin avdd.t110 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X641 a_8877_n2876# a_8777_n2964# dvss.t136 dvss.t135 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X642 comparator_0.vinn.t37 rstring_mux_0.vtrip_decoded_b_avdd[4] rstring_mux_0.vtrip4.t9 avdd.t497 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X643 porb.t23 sky130_fd_sc_hd__inv_4_1.Y dvdd.t155 dvdd.t154 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X644 avdd.t212 a_8877_n1142# a_9570_n2256# avdd.t211 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.1365 ps=1.49 w=0.42 l=1
X645 dcomp.t9 sky130_fd_sc_hd__inv_4_3.Y dvss.t746 dvss.t745 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X646 avdd.t313 avdd.t311 avdd.t312 avdd.t221 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=8
X647 dvss.t321 a_n3778_7859# a_n2571_7523# dvss.t320 sky130_fd_pr__nfet_g5v0d10v5 ad=0.121875 pd=1.075 as=0.19875 ps=2.03 w=0.75 l=0.5
X648 a_1643_n11914# a_1265_n19314# avss.t63 sky130_fd_pr__res_xhigh_po_1p41 l=35
X649 vin avss.t196 vin avss.t197 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=23.2 ps=169.28 w=5 l=0.6
X650 porb.t9 sky130_fd_sc_hd__inv_4_1.Y dvss.t509 dvss.t508 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X651 avdd.t35 a_1122_n3990# a_429_n2876# avdd.t34 sky130_fd_pr__pfet_g5v0d10v5 ad=0.2142 pd=1.99 as=0.2142 ps=1.99 w=0.42 l=1
X652 comparator_0.n1 comparator_0.n0 avdd.t419 avdd.t418 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.6
X653 avdd.t192 comparator_0.vnn comparator_0.vpp avdd.t179 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X654 avss.t357 sky130_fd_sc_hvl__inv_16_0.A porb_h.t7 avss.t356 sky130_fd_pr__nfet_g5v0d10v5 ad=0.2025 pd=2.04 as=0.105 ps=1.03 w=0.75 l=0.5
X655 dvdd.t197 por_unbuf.t5 a_n3878_7771# dvdd.t196 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X656 dvss.t168 schmitt_trigger_0.in.t5 schmitt_trigger_0.m.t5 dvss.t167 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X657 a_429_n2876# a_329_n2964# dvss.t100 dvss.t99 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X658 dvss.t595 sky130_fd_sc_hd__inv_4_1.A sky130_fd_sc_hd__inv_4_1.Y dvss.t594 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X659 a_8877_n1142# a_8777_n1230# dvss.t199 dvss.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X660 a_n5639_n2212# a_n6007_n1230# dvdd.t82 dvdd.t81 sky130_fd_pr__pfet_01v8_hvt ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X661 dvss.t134 a_8777_n2964# a_8877_n2876# dvss.t133 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X662 a_1643_n11914# a_2021_n19314# avss.t7 sky130_fd_pr__res_xhigh_po_1p41 l=35
X663 dvdd.t213 rc_osc_0.in rc_osc_0.m dvdd.t212 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X664 avdd.t310 avdd.t308 avdd.t309 avdd.t221 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=8
X665 rstring_mux_0.vtop.t8 rstring_mux_0.ena_b avdd.t469 avdd.t468 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X666 porb_h.t6 sky130_fd_sc_hvl__inv_16_0.A avss.t355 avss.t354 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.19875 ps=2.03 w=0.75 l=0.5
X667 comparator_0.vt comparator_0.vinn.t58 comparator_0.vnn comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X668 avss.t195 avss.t192 avss.t194 avss.t193 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=8
X669 dvdd.t294 sky130_fd_sc_hd__inv_4_3.Y dcomp.t22 dvdd.t293 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X670 pwup_filt.t24 sky130_fd_sc_hd__inv_4_0.Y dvdd.t27 dvdd.t26 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X671 a_3234_n2256# a_2809_n2212# dvss.t332 dvss.t331 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X672 rstring_mux_0.vtrip_decoded_b_avdd[1] rstring_mux_0.vtrip_decoded_avdd[1] avdd.t9 avdd.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X673 avss.t403 a_9581_n19314# avss.t402 sky130_fd_pr__res_xhigh_po_1p41 l=35
X674 comparator_0.vt comparator_0.vinn.t59 comparator_0.vnn comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X675 avdd.t191 comparator_0.vnn comparator_0.vpp avdd.t179 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X676 comparator_0.vnn comparator_0.vnn avdd.t190 avdd.t186 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X677 avdd.t585 comparator_1.n0 comparator_1.n1 avdd.t584 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X678 a_n11219_9395# a_n10841_1995# avss.t15 sky130_fd_pr__res_xhigh_po_1p41 l=35
X679 dvss.t98 a_329_n2964# a_429_n2876# dvss.t97 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X680 avdd.t307 avdd.t305 avdd.t306 avdd.t230 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=8
X681 a_8877_n2876# a_8777_n2964# dvss.t132 dvss.t131 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X682 avdd.t467 rstring_mux_0.ena_b rstring_mux_0.vtop.t7 avdd.t466 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X683 comparator_1.vt vin comparator_1.vpp comparator_1.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X684 ibias_gen_0.vp0.t4 rstring_mux_0.ena avdd.t516 avdd.t515 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X685 comparator_0.vinn.t31 avdd.t303 comparator_0.vinn.t31 avdd.t304 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=0.6
X686 porb.t8 sky130_fd_sc_hd__inv_4_1.Y dvss.t507 dvss.t506 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X687 rstring_mux_0.vtrip_decoded_avdd[0] a_1636_n3212# avdd.t580 avdd.t396 sky130_fd_pr__pfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.24375 ps=1.825 w=1.5 l=0.5
X688 avdd.t39 a_6765_n2876# a_7972_n3212# avdd.t38 sky130_fd_pr__pfet_g5v0d10v5 ad=0.24375 pd=1.825 as=0.3975 ps=3.53 w=1.5 l=0.5
X689 avdd.t620 a_3234_n3990# a_2541_n2876# avdd.t619 sky130_fd_pr__pfet_g5v0d10v5 ad=0.2142 pd=1.99 as=0.2142 ps=1.99 w=0.42 l=1
X690 rstring_mux_0.vtrip_decoded_b_avdd[5] rstring_mux_0.vtrip_decoded_avdd[5] avdd.t206 avdd.t205 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X691 rstring_mux_0.vtrip_decoded_b_avdd[1] rstring_mux_0.vtrip_decoded_avdd[1] avss.t18 avss.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X692 comparator_1.vnn comparator_1.vpp avdd.t642 avdd.t73 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X693 avss.t383 comparator_1.n0 comparator_1.n1 avss.t382 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X694 comparator_1.vt vin comparator_1.vpp comparator_1.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X695 a_5346_n3990# a_4921_n3946# dvss.t108 dvss.t107 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X696 porb_h.t25 sky130_fd_sc_hvl__inv_16_0.A avdd.t557 avdd.t556 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X697 ibias_gen_0.vn0.t3 ibias_gen_0.ena_b avss.t319 avss.t318 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X698 dvss.t627 a_6765_n1142# a_7972_n1478# dvss.t175 sky130_fd_pr__nfet_g5v0d10v5 ad=0.121875 pd=1.075 as=0.19875 ps=2.03 w=0.75 l=0.5
X699 dvdd.t109 dvss.t773 a_329_n2964# dvdd.t108 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X700 comparator_0.vt avss.t425 comparator_0.vnn comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=8
X701 avss.t51 comparator_0.n1 dcomp3v3uv avss.t50 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X702 a_10515_n2156# a_10515_n1026# avdd.t44 avdd.t42 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.1197 ps=1.41 w=0.42 l=0.5
X703 rstring_mux_0.vtop.t6 rstring_mux_0.ena_b avdd.t465 avdd.t464 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X704 avdd.t58 comparator_0.n1 dcomp3v3uv avdd.t57 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X705 vin rstring_mux_0.otrip_decoded_avdd[1] rstring_mux_0.vtrip1.t9 avss.t299 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X706 a_n10279_n22711# a_12321_n22333# dvss.t324 sky130_fd_pr__res_xhigh_po_1p41 l=111
X707 dcomp3v3 comparator_1.n1 avdd.t27 avdd.t26 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X708 a_n9707_9395# a_n10085_1995# avss.t408 sky130_fd_pr__res_xhigh_po_1p41 l=35
X709 por.t22 sky130_fd_sc_hd__inv_4_4.Y dvdd.t255 dvdd.t254 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X710 avdd.t437 a_n5907_n1142# a_n5214_n2256# avdd.t436 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.1365 ps=1.49 w=0.42 l=1
X711 dvss.t605 a_n1783_n1230# a_n1683_n1142# dvss.t604 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X712 avdd.t555 sky130_fd_sc_hvl__inv_16_0.A porb_h.t24 avdd.t554 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X713 a_5423_n11914# a_5045_n19314# avss.t260 sky130_fd_pr__res_xhigh_po_1p41 l=35
X714 avdd.t302 avdd.t301 avdd.t302 avdd.t234 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=8
X715 avdd.t300 avdd.t298 avdd.t299 avdd.t230 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=8
X716 comparator_1.vt avss.t426 comparator_1.vnn comparator_1.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=8
X717 a_n12721_n11914# a_n13099_n19314# avss.t242 sky130_fd_pr__res_xhigh_po_1p41 l=35
X718 comparator_0.vm comparator_0.vnn avdd.t189 avdd.t177 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X719 dvss.t633 vl sky130_fd_sc_hd__inv_4_3.Y dvss.t632 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X720 dvdd.t107 dvss.t774 a_4553_n1230# dvdd.t106 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X721 rstring_mux_0.vtrip_decoded_avdd[2] a_3748_n3212# avdd.t577 avdd.t576 sky130_fd_pr__pfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.24375 ps=1.825 w=1.5 l=0.5
X722 rstring_mux_0.vtrip3.t0 rstring_mux_0.vtrip4.t0 avss.t2 sky130_fd_pr__res_xhigh_po_1p41 l=35
X723 avdd.t37 a_5346_n3990# a_4653_n2876# avdd.t36 sky130_fd_pr__pfet_g5v0d10v5 ad=0.2142 pd=1.99 as=0.2142 ps=1.99 w=0.42 l=1
X724 a_7458_n3990# a_7033_n3946# dvss.t716 dvss.t715 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X725 schmitt_trigger_0.in.t6 dvss.t169 sky130_fd_pr__cap_mim_m3_2 l=30 w=30
X726 porb.t22 sky130_fd_sc_hd__inv_4_1.Y dvdd.t153 dvdd.t152 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X727 rstring_mux_0.otrip_decoded_b_avdd[3] rstring_mux_0.otrip_decoded_avdd[3] avss.t254 avss.t253 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X728 vin avdd.t296 vin avdd.t297 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=0.6
X729 sky130_fd_sc_hd__inv_4_4.Y por_unbuf.t6 dvdd.t199 dvdd.t198 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X730 rstring_mux_0.vtrip3.t5 rstring_mux_0.vtrip2.t3 avss.t243 sky130_fd_pr__res_xhigh_po_1p41 l=35
X731 avss.t191 avss.t189 avss.t190 avss.t146 sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0 ps=0 w=5 l=8
X732 a_n1683_n1142# a_n1783_n1230# dvss.t603 dvss.t602 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X733 rc_osc_0.m rc_osc_0.n.t8 dvdd.t177 dvdd.t176 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X734 vin avss.t187 vin avss.t188 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=0.6
X735 comparator_1.ena_b rstring_mux_0.ena avss.t326 avss.t325 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X736 avdd.t295 avdd.t294 avdd.t295 avdd.t234 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=8
X737 pwup_filt.t7 sky130_fd_sc_hd__inv_4_0.Y dvss.t72 dvss.t71 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X738 a_4921_n2212# a_4553_n1230# dvdd.t121 dvdd.t120 sky130_fd_pr__pfet_01v8_hvt ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X739 dcomp3v3uv comparator_0.n1 avdd.t56 avdd.t55 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X740 comparator_0.vnn comparator_0.vnn avdd.t188 avdd.t186 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X741 avdd.t293 avdd.t291 avdd.t292 avdd.t230 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=8
X742 a_9570_n2256# a_9145_n2212# dvss.t29 dvss.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X743 dvss.t262 a_10514_n3890# a_10873_n3956# dvss.t261 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.19875 ps=2.03 w=0.75 l=0.5
X744 dvdd.t61 schmitt_trigger_0.out.t8 sky130_fd_sc_hd__inv_4_0.Y dvdd.t60 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X745 comparator_0.vt vbg_1v2.t20 comparator_0.vpp comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X746 comparator_1.vnn vbg_1v2.t21 comparator_1.vt comparator_1.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X747 dvss.t48 a_2441_n1230# a_2541_n1142# dvss.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X748 dvss.t240 a_n1415_n2212# a_n990_n2256# dvss.t239 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X749 schmitt_trigger_0.in.t7 dvss.t170 sky130_fd_pr__cap_mim_m3_2 l=30 w=30
X750 avdd.t71 comparator_1.vnn comparator_1.vpp avdd.t65 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X751 ibias_gen_0.vn1.t4 avss.t185 ibias_gen_0.vp1.t8 avss.t186 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X752 dcomp.t8 sky130_fd_sc_hd__inv_4_3.Y dvss.t744 dvss.t743 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X753 avdd.t654 a_n8019_n1142# a_n7326_n2256# avdd.t653 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.1365 ps=1.49 w=0.42 l=1
X754 dvss.t363 a_n3895_n1230# a_n3795_n1142# dvss.t362 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X755 sky130_fd_sc_hd__inv_4_0.Y schmitt_trigger_0.out.t9 dvss.t154 dvss.t153 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X756 dvdd.t151 sky130_fd_sc_hd__inv_4_1.Y porb.t21 dvdd.t150 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X757 a_2541_n2876# a_2441_n2964# dvss.t432 dvss.t431 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X758 a_n990_n3990# a_n1415_n3946# dvss.t23 dvss.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X759 avdd.t290 avdd.t288 avdd.t289 avdd.t221 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=8
X760 comparator_0.vinn.t9 rstring_mux_0.vtrip_decoded_avdd[6] rstring_mux_0.vtrip6.t4 avss.t94 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X761 ibias_gen_0.vn0.t13 vbg_1v2.t22 ibias_gen_0.vstart.t5 avss.t129 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X762 dvdd.t105 dvss.t775 a_6665_n1230# dvdd.t104 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X763 a_n3795_n2876# a_n3895_n2964# dvss.t410 dvss.t409 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X764 avss.t353 sky130_fd_sc_hvl__inv_16_0.A porb_h.t5 avss.t352 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X765 avdd.t162 a_n3778_7859# a_n3085_6745# avdd.t161 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.1365 ps=1.49 w=0.42 l=1
X766 dvss.t559 a_n5907_n1142# a_n4700_n1478# dvss.t558 sky130_fd_pr__nfet_g5v0d10v5 ad=0.121875 pd=1.075 as=0.19875 ps=2.03 w=0.75 l=0.5
X767 a_n5214_n2256# a_n5639_n2212# dvss.t40 dvss.t39 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X768 a_n7751_n3946# a_n8119_n2964# dvdd.t275 dvdd.t274 sky130_fd_pr__pfet_01v8_hvt ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X769 avdd.t587 a_7458_n3990# a_6765_n2876# avdd.t586 sky130_fd_pr__pfet_g5v0d10v5 ad=0.2142 pd=1.99 as=0.2142 ps=1.99 w=0.42 l=1
X770 rc_osc_0.vr dvss.t293 dvss.t295 dvss.t294 sky130_fd_pr__nfet_01v8 ad=0.1475 pd=1.295 as=0.145 ps=1.29 w=1 l=0.6
X771 avdd.t606 comparator_0.vpp comparator_0.vpp avdd.t179 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X772 a_n3102_n2256# a_n3527_n2212# dvss.t7 dvss.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X773 a_n990_n2256# a_n1415_n2212# dvss.t238 dvss.t237 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X774 dvss.t251 a_10874_n2222# vl dvss.t250 sky130_fd_pr__nfet_01v8 ad=0.1961 pd=2.01 as=0.1961 ps=2.01 w=0.74 l=0.15
X775 avss.t283 comparator_1.vm comparator_1.n0 avss.t282 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X776 dvdd.t75 schmitt_trigger_0.in.t8 schmitt_trigger_0.m.t9 dvdd.t74 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X777 pwup_filt.t23 sky130_fd_sc_hd__inv_4_0.Y dvdd.t25 dvdd.t24 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X778 vin rstring_mux_0.otrip_decoded_b_avdd[2] rstring_mux_0.vtrip2.t8 avdd.t627 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X779 a_8447_n11914# a_8825_n19314# avss.t9 sky130_fd_pr__res_xhigh_po_1p41 l=35
X780 pwup_filt.t6 sky130_fd_sc_hd__inv_4_0.Y dvss.t70 dvss.t69 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X781 rstring_mux_0.vtrip_decoded_avdd[1] a_1636_n1478# dvss.t569 dvss.t175 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.121875 ps=1.075 w=0.75 l=0.5
X782 dvss.t430 a_2441_n2964# a_2541_n2876# dvss.t429 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X783 rstring_mux_0.vtrip0.t6 rstring_mux_0.vtrip_decoded_b_avdd[0] comparator_0.vinn.t39 avdd.t507 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X784 a_10873_n2760# a_10873_n3956# dvdd.t277 dvdd.t276 sky130_fd_pr__pfet_01v8_hvt ad=0.2968 pd=2.77 as=0.1568 ps=1.4 w=1.12 l=0.15
X785 rstring_mux_0.vtrip0.t1 rstring_mux_0.otrip_decoded_b_avdd[0] vin avdd.t140 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=0.6
X786 a_n3085_6745# a_n3510_6789# dvss.t450 dvss.t449 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X787 dvss.t593 sky130_fd_sc_hd__inv_4_1.A sky130_fd_sc_hd__inv_4_1.Y dvss.t592 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X788 a_9203_n11914# a_8825_n19314# avss.t270 sky130_fd_pr__res_xhigh_po_1p41 l=35
X789 dvss.t179 a_n6007_n1230# a_n5907_n1142# dvss.t178 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X790 a_n5917_n11914# a_n5539_n19314# avss.t5 sky130_fd_pr__res_xhigh_po_1p41 l=35
X791 comparator_0.vnn comparator_0.vnn avdd.t187 avdd.t186 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X792 rstring_mux_0.vtrip7.t6 rstring_mux_0.vtrip_decoded_avdd[7] comparator_0.vinn.t25 avss.t266 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X793 a_n5907_n2876# a_n6007_n2964# dvss.t381 dvss.t380 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X794 avdd.t287 avdd.t285 avdd.t286 avdd.t230 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=8
X795 a_n5907_n2876# a_n6007_n2964# dvss.t379 dvss.t378 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X796 a_4653_n2876# a_4553_n2964# dvss.t274 dvss.t273 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X797 comparator_0.n0 comparator_0.ena_b avss.t110 avss.t109 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X798 avdd.t284 avdd.t283 avdd.t284 avdd.t240 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=8
X799 dvdd.t292 sky130_fd_sc_hd__inv_4_3.Y dcomp.t21 dvdd.t291 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X800 avdd.t592 a_2541_n2876# a_3748_n3212# avdd.t576 sky130_fd_pr__pfet_g5v0d10v5 ad=0.24375 pd=1.825 as=0.3975 ps=3.53 w=1.5 l=0.5
X801 avss.t297 rstring_mux_0.ena_b rstring_mux_0.vtop.t0 avss.t296 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X802 avdd.t70 comparator_1.vnn comparator_1.vpp avdd.t65 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X803 avss.t125 ibias_gen_0.vn1.t15 ibias_gen_0.vp1.t5 avss.t120 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=8
X804 a_n7326_n2256# a_n7751_n2212# dvss.t462 dvss.t461 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X805 avdd.t571 a_9570_n3990# a_8877_n2876# avdd.t570 sky130_fd_pr__pfet_g5v0d10v5 ad=0.2142 pd=1.99 as=0.2142 ps=1.99 w=0.42 l=1
X806 vin rstring_mux_0.otrip_decoded_avdd[3] rstring_mux_0.vtrip3.t6 avss.t252 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X807 rstring_mux_0.vtrip4.t8 rstring_mux_0.vtrip_decoded_b_avdd[4] comparator_0.vinn.t38 avdd.t496 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X808 comparator_1.vnn comparator_1.vpp avdd.t641 avdd.t73 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X809 comparator_1.vt vin comparator_1.vpp comparator_1.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X810 a_n8019_n1142# a_n8119_n1230# dvss.t616 dvss.t615 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X811 a_n1415_n3946# a_n1783_n2964# dvss.t349 dvss.t348 sky130_fd_pr__nfet_01v8 ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X812 comparator_0.vt comparator_0.vn avss.t391 avss.t109 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X813 dvss.t448 a_n3510_6789# a_n3085_6745# dvss.t447 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X814 ibias_gen_0.vstart.t4 vbg_1v2.t23 ibias_gen_0.vn0.t12 avss.t128 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=0.6
X815 dvss.t704 a_n8119_n2964# a_n8019_n2876# dvss.t703 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X816 comparator_0.vinn.t14 avss.t183 comparator_0.vinn.t14 avss.t184 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=0.6
X817 porb.t7 sky130_fd_sc_hd__inv_4_1.Y dvss.t505 dvss.t504 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X818 a_3911_n11914# a_3533_n19314# avss.t233 sky130_fd_pr__res_xhigh_po_1p41 l=35
X819 vin rstring_mux_0.otrip_decoded_avdd[6] rstring_mux_0.vtrip6.t8 avss.t309 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X820 a_1122_n2256# a_697_n2212# dvss.t209 dvss.t208 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X821 dvss.t260 a_10514_n3890# a_10873_n3956# dvss.t259 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.105 ps=1.03 w=0.75 l=0.5
X822 comparator_1.vnn comparator_1.vpp avdd.t640 avdd.t73 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X823 avss.t182 avss.t180 avss.t181 avss.t146 sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0 ps=0 w=5 l=8
X824 a_10874_n1026# a_10515_n1026# dvss.t122 dvss.t119 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.105 ps=1.03 w=0.75 l=0.5
X825 a_n8019_n2876# a_n8119_n2964# dvss.t702 dvss.t701 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X826 a_6765_n2876# a_6665_n2964# dvss.t393 dvss.t392 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X827 dvss.t336 force_pdnb.t0 a_8777_n2964# dvss.t335 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X828 comparator_0.ibias ibias_gen_0.vp.t10 avdd.t431 avdd.t430 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X829 dvss.t330 a_2809_n2212# a_3234_n2256# dvss.t329 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X830 a_n8019_n2876# a_n8119_n2964# dvss.t700 dvss.t699 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X831 rstring_mux_0.otrip_decoded_b_avdd[0] rstring_mux_0.otrip_decoded_avdd[0] avdd.t501 avdd.t500 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X832 dvdd.t201 por_unbuf.t7 sky130_fd_sc_hd__inv_4_1.A dvdd.t200 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X833 avdd.t624 a_4653_n2876# a_5860_n3212# avdd.t452 sky130_fd_pr__pfet_g5v0d10v5 ad=0.24375 pd=1.825 as=0.3975 ps=3.53 w=1.5 l=0.5
X834 dvss.t566 a_10514_n2760# a_10873_n2760# dvss.t565 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X835 rstring_mux_0.vtrip5.t9 rstring_mux_0.vtrip6.t9 avss.t405 sky130_fd_pr__res_xhigh_po_1p41 l=35
X836 osc_ck.t0 rc_osc_0.ena_b rc_osc_0.vr dvdd.t80 sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.1475 ps=1.295 w=1 l=0.18
X837 dvss.t116 dcomp3v3 a_10515_n1026# dvss.t115 sky130_fd_pr__nfet_g5v0d10v5 ad=0.178875 pd=1.26 as=0.1197 ps=1.41 w=0.42 l=0.5
X838 dvss.t207 a_697_n2212# a_1122_n2256# dvss.t206 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X839 a_n3527_n3946# a_n3895_n2964# dvss.t408 dvss.t407 sky130_fd_pr__nfet_01v8 ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X840 a_429_n2876# a_329_n2964# dvss.t96 dvss.t95 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X841 vin rstring_mux_0.otrip_decoded_avdd[7] rstring_mux_0.vtrip7.t3 avss.t99 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X842 dvss.t479 osc_ena.t2 rc_osc_0.ena_b dvss.t478 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.6
X843 a_n14243_9395# a_n13865_1995# avss.t69 sky130_fd_pr__res_xhigh_po_1p41 l=35
X844 porb.t6 sky130_fd_sc_hd__inv_4_1.Y dvss.t503 dvss.t502 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X845 comparator_0.vinn.t3 rstring_mux_0.vtrip_decoded_avdd[4] rstring_mux_0.vtrip4.t1 avss.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X846 avdd.t639 comparator_1.vpp comparator_1.vnn avdd.t80 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X847 por.t21 sky130_fd_sc_hd__inv_4_4.Y dvdd.t253 dvdd.t252 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X848 a_3234_n2256# a_2809_n2212# dvss.t328 dvss.t327 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X849 rstring_mux_0.vtrip7.t0 rstring_mux_0.vtrip6.t0 avss.t1 sky130_fd_pr__res_xhigh_po_1p41 l=35
X850 a_n9697_n11914# a_n9319_n19314# avss.t232 sky130_fd_pr__res_xhigh_po_1p41 l=35
X851 avdd.t282 avdd.t281 avdd.t282 avdd.t240 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=8
X852 comparator_0.vt vbg_1v2.t24 comparator_0.vpp comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X853 schmitt_trigger_0.out.t1 schmitt_trigger_0.m.t16 dvdd.t99 dvdd.t98 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X854 avdd.t13 a_n3795_n1142# a_n3102_n2256# avdd.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.1365 ps=1.49 w=0.42 l=1
X855 dvss.t444 a_2809_n3946# a_3234_n3990# dvss.t443 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X856 a_n10279_n23467# a_12321_n23845# dvss.t768 sky130_fd_pr__res_xhigh_po_1p41 l=111
X857 comparator_1.vn comparator_1.ena_b avss.t287 avss.t286 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X858 pwup_filt.t5 sky130_fd_sc_hd__inv_4_0.Y dvss.t68 dvss.t67 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X859 dvss.t94 a_329_n2964# a_429_n2876# dvss.t93 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X860 comparator_0.vt avss.t427 comparator_0.vnn comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=8
X861 comparator_0.vt vbg_1v2.t25 comparator_0.vpp comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X862 avdd.t605 comparator_0.vpp comparator_0.vnn avdd.t182 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X863 dvss.t662 sky130_fd_sc_hd__inv_4_4.Y por.t6 dvss.t661 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X864 rstring_mux_0.otrip_decoded_avdd[7] a_n476_n1478# dvss.t236 dvss.t175 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.121875 ps=1.075 w=0.75 l=0.5
X865 comparator_1.vnn vbg_1v2.t26 comparator_1.vt comparator_1.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X866 dvss.t221 a_4921_n2212# a_5346_n2256# dvss.t220 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X867 comparator_0.vinn.t24 rstring_mux_0.vtrip_decoded_avdd[7] rstring_mux_0.vtrip7.t5 avss.t265 sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=0.6
X868 avdd.t25 comparator_1.n1 dcomp3v3 avdd.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.6
X869 avss.t400 a_n27208_n10337# avss.t0 sky130_fd_pr__res_xhigh_po_1p41 l=35
X870 a_n5639_n3946# a_n6007_n2964# dvss.t377 dvss.t376 sky130_fd_pr__nfet_01v8 ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X871 porb_h.t23 sky130_fd_sc_hvl__inv_16_0.A avdd.t553 avdd.t552 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X872 sky130_fd_sc_hd__inv_4_0.Y schmitt_trigger_0.out.t10 dvss.t156 dvss.t155 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X873 dvdd.t149 sky130_fd_sc_hd__inv_4_1.Y porb.t20 dvdd.t148 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X874 rstring_mux_0.vtrip5.t3 rstring_mux_0.vtrip_decoded_avdd[5] comparator_0.vinn.t22 avss.t247 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X875 comparator_1.vt avss.t428 comparator_1.vnn comparator_1.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=8
X876 ibias_gen_0.ibias0 ibias_gen_0.vp.t11 avdd.t433 avdd.t432 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X877 rstring_mux_0.vtrip5.t2 rstring_mux_0.otrip_decoded_b_avdd[5] vin avdd.t158 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X878 a_5346_n2256# a_4921_n2212# dvss.t219 dvss.t218 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X879 rstring_mux_0.vtrip_decoded_b_avdd[3] rstring_mux_0.vtrip_decoded_avdd[3] avdd.t106 avdd.t105 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X880 a_n4405_n11914# a_n4783_n19314# avss.t238 sky130_fd_pr__res_xhigh_po_1p41 l=35
X881 avss.t49 comparator_0.n1 dcomp3v3uv avss.t48 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X882 comparator_0.vpp avss.t429 avdd.t166 avdd.t165 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X883 vin rstring_mux_0.otrip_decoded_avdd[5] rstring_mux_0.vtrip5.t7 avss.t395 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X884 avdd.t551 sky130_fd_sc_hvl__inv_16_0.A porb_h.t22 avdd.t550 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X885 avdd.t280 avdd.t278 avdd.t279 avdd.t230 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=8
X886 a_9570_n3990# a_9145_n3946# dvss.t646 dvss.t645 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X887 avdd.t638 comparator_1.vpp comparator_1.vnn avdd.t80 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X888 avss.t179 avss.t178 avss.t179 avss.t171 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=8
X889 avdd.t441 a_429_n1142# a_1122_n2256# avdd.t440 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.1365 ps=1.49 w=0.42 l=1
X890 avdd.t277 avdd.t276 avdd.t277 avdd.t240 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=8
X891 comparator_1.vnn avss.t430 comparator_1.vt comparator_1.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=8
X892 dvss.t231 a_7033_n2212# a_7458_n2256# dvss.t230 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X893 avdd.t54 comparator_0.n1 dcomp3v3uv avdd.t53 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.6
X894 a_n15479_n3901# ibias_gen_0.isrc_sel ibias_gen_0.vn1.t9 avss.t336 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X895 dcomp.t7 sky130_fd_sc_hd__inv_4_3.Y dvss.t742 dvss.t741 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X896 dvss.t361 a_2541_n1142# a_3748_n1478# dvss.t175 sky130_fd_pr__nfet_g5v0d10v5 ad=0.121875 pd=1.075 as=0.19875 ps=2.03 w=0.75 l=0.5
X897 por.t20 sky130_fd_sc_hd__inv_4_4.Y dvdd.t251 dvdd.t250 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X898 rstring_mux_0.otrip_decoded_avdd[2] a_n4700_n3212# dvss.t446 dvss.t445 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.121875 ps=1.075 w=0.75 l=0.5
X899 a_7458_n3990# a_7033_n3946# dvss.t714 dvss.t713 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X900 rstring_mux_0.vtrip_decoded_b_avdd[3] rstring_mux_0.vtrip_decoded_avdd[3] avss.t74 avss.t73 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X901 comparator_0.n0 comparator_0.vpp avdd.t604 avdd.t186 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X902 avdd.t23 comparator_1.n1 dcomp3v3 avdd.t22 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X903 schmitt_trigger_0.m.t2 schmitt_trigger_0.out.t11 dvdd.t63 dvdd.t62 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X904 dvdd.t179 rc_osc_0.n.t9 osc_ck.t4 dvdd.t178 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X905 rc_osc_0.m rc_osc_0.n.t10 dvss.t537 dvss.t536 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X906 dvss.t347 a_n1783_n2964# a_n1683_n2876# dvss.t346 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X907 avss.t177 avss.t176 avss.t177 avss.t109 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=8
X908 ibias_gen_0.vp0.t10 ibias_gen_0.vn0.t20 ibias_gen_0.vr.t3 avss.t67 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X909 sky130_fd_sc_hd__inv_4_1.A por_unbuf.t8 dvss.t545 dvss.t544 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X910 a_2809_n2212# a_2441_n1230# dvss.t46 dvss.t45 sky130_fd_pr__nfet_01v8 ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X911 avdd.t603 comparator_0.vpp comparator_0.vnn avdd.t182 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X912 pwup_filt.t22 sky130_fd_sc_hd__inv_4_0.Y dvdd.t23 dvdd.t22 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X913 dvss.t5 a_n3527_n2212# a_n3102_n2256# dvss.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X914 avdd.t92 a_n5214_n3990# a_n5907_n2876# avdd.t91 sky130_fd_pr__pfet_g5v0d10v5 ad=0.2142 pd=1.99 as=0.2142 ps=1.99 w=0.42 l=1
X915 porb.t5 sky130_fd_sc_hd__inv_4_1.Y dvss.t501 dvss.t500 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X916 a_n3102_n3990# a_n3527_n3946# dvss.t476 dvss.t475 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X917 a_2541_n2876# a_2441_n2964# dvss.t428 dvss.t427 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X918 dvss.t292 dvss.t290 a_4553_n2964# dvss.t291 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X919 rstring_mux_0.otrip_decoded_b_avdd[5] rstring_mux_0.otrip_decoded_avdd[5] avdd.t623 avdd.t622 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X920 avss.t351 sky130_fd_sc_hvl__inv_16_0.A porb_h.t4 avss.t350 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X921 avdd.t216 a_2541_n1142# a_3234_n2256# avdd.t215 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.1365 ps=1.49 w=0.42 l=1
X922 dvss.t27 a_9145_n2212# a_9570_n2256# dvss.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X923 rstring_mux_0.vtrip7.t2 rstring_mux_0.otrip_decoded_b_avdd[7] vin avdd.t5 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X924 dcomp3v3 comparator_1.n1 avss.t30 avss.t29 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X925 a_n8185_n11914# a_n7807_n19314# avss.t20 sky130_fd_pr__res_xhigh_po_1p41 l=35
X926 comparator_0.vinn.t43 rstring_mux_0.vtrip_decoded_avdd[2] rstring_mux_0.vtrip2.t6 avss.t380 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X927 a_n3102_n2256# a_n3527_n2212# dvss.t3 dvss.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X928 rstring_mux_0.otrip_decoded_avdd[0] a_n6812_n3212# dvss.t601 dvss.t600 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.121875 ps=1.075 w=0.75 l=0.5
X929 a_9570_n3990# a_9145_n3946# dvss.t644 dvss.t643 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X930 dvss.t474 a_n3527_n3946# a_n3102_n3990# dvss.t473 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X931 dvss.t21 a_n1415_n3946# a_n990_n3990# dvss.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X932 a_4921_n3946# a_4553_n2964# dvss.t272 dvss.t271 sky130_fd_pr__nfet_01v8 ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X933 comparator_1.vpp comparator_1.vpp avdd.t637 avdd.t63 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X934 sky130_fd_sc_hvl__inv_16_0.A sky130_fd_sc_hvl__inv_4_0.A avss.t87 avss.t86 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.21375 ps=2.07 w=0.75 l=0.5
X935 dvss.t406 a_n3895_n2964# a_n3795_n2876# dvss.t405 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X936 dvss.t564 a_10514_n2760# a_10873_n2760# dvss.t563 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.19875 ps=2.03 w=0.75 l=0.5
X937 rstring_mux_0.vtrip_decoded_b_avdd[2] rstring_mux_0.vtrip_decoded_avdd[2] avdd.t575 avdd.t574 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X938 a_n11209_n11914# a_n11587_n19314# avss.t68 sky130_fd_pr__res_xhigh_po_1p41 l=35
X939 comparator_0.vpp comparator_0.vnn avdd.t185 avdd.t177 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X940 comparator_0.vinn.t30 avdd.t274 comparator_0.vinn.t30 avdd.t275 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=0.6
X941 avdd.t273 avdd.t271 avdd.t272 avdd.t230 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=8
X942 schmitt_trigger_0.m.t3 schmitt_trigger_0.out.t12 dvss.t158 dvss.t157 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X943 comparator_0.ena_b avss.t173 avss.t175 avss.t174 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X944 a_7033_n2212# a_6665_n1230# dvss.t583 dvss.t582 sky130_fd_pr__nfet_01v8 ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X945 comparator_1.vt vin comparator_1.vpp comparator_1.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X946 dvss.t38 a_n5639_n2212# a_n5214_n2256# dvss.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X947 avdd.t589 a_n7326_n3990# a_n8019_n2876# avdd.t588 sky130_fd_pr__pfet_g5v0d10v5 ad=0.2142 pd=1.99 as=0.2142 ps=1.99 w=0.42 l=1
X948 dvss.t354 a_4553_n1230# a_4653_n1142# dvss.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X949 a_n5214_n3990# a_n5639_n3946# dvss.t150 dvss.t149 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X950 avss.t293 comparator_1.vn comparator_1.vt avss.t282 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X951 dvss.t338 otrip_decoded[7].t0 a_n1783_n1230# dvss.t337 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X952 dvss.t289 dvss.t287 a_6665_n2964# dvss.t288 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X953 comparator_0.vt avss.t431 comparator_0.vnn comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=8
X954 porb.t4 sky130_fd_sc_hd__inv_4_1.Y dvss.t499 dvss.t498 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X955 avdd.t411 a_4653_n1142# a_5346_n2256# avdd.t410 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.1365 ps=1.49 w=0.42 l=1
X956 a_4653_n2876# a_4553_n2964# dvss.t270 dvss.t269 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X957 a_n990_n3990# a_n1415_n3946# dvss.t19 dvss.t18 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X958 comparator_0.vnn avss.t432 comparator_0.vt comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=8
X959 vin rstring_mux_0.otrip_decoded_b_avdd[4] rstring_mux_0.vtrip4.t3 avdd.t109 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X960 por.t5 sky130_fd_sc_hd__inv_4_4.Y dvss.t660 dvss.t659 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X961 comparator_0.vt avss.t433 comparator_0.vnn comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=8
X962 porb_h.t21 sky130_fd_sc_hvl__inv_16_0.A avdd.t549 avdd.t548 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X963 comparator_0.vpp vbg_1v2.t27 comparator_0.vt comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X964 comparator_0.vinn.t4 rstring_mux_0.vtrip_decoded_b_avdd[6] rstring_mux_0.vtrip6.t2 avdd.t94 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X965 comparator_1.n0 comparator_1.vm avss.t281 avss.t280 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X966 dvdd.t203 por_unbuf.t9 sky130_fd_sc_hd__inv_4_4.Y dvdd.t202 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X967 a_n5214_n2256# a_n5639_n2212# dvss.t36 dvss.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X968 dvss.t391 a_6665_n2964# a_6765_n2876# dvss.t390 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X969 dvss.t148 a_n5639_n3946# a_n5214_n3990# dvss.t147 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X970 avdd.t602 comparator_0.vpp comparator_0.vnn avdd.t182 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X971 sky130_fd_sc_hd__inv_4_4.Y por_unbuf.t10 dvss.t547 dvss.t546 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X972 rstring_mux_0.otrip_decoded_b_avdd[7] rstring_mux_0.otrip_decoded_avdd[7] avdd.t126 avdd.t125 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X973 avdd.t270 avdd.t269 avdd.t270 avdd.t234 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=8
X974 comparator_1.vt avss.t434 comparator_1.vnn comparator_1.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=8
X975 pwup_filt.t4 sky130_fd_sc_hd__inv_4_0.Y dvss.t66 dvss.t65 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X976 a_1122_n2256# a_697_n2212# dvss.t205 dvss.t204 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X977 a_9145_n2212# a_8777_n1230# dvss.t198 dvss.t197 sky130_fd_pr__nfet_01v8 ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X978 comparator_0.vnn avss.t435 comparator_0.vt comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=8
X979 dvss.t460 a_n7751_n2212# a_n7326_n2256# dvss.t459 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X980 comparator_0.vnn comparator_0.vinn.t60 comparator_0.vt comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X981 comparator_1.vpp comparator_1.vpp avdd.t636 avdd.t63 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X982 dvss.t631 vl sky130_fd_sc_hd__inv_4_3.Y dvss.t630 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X983 a_n7326_n3990# a_n7751_n3946# dvss.t688 dvss.t687 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X984 comparator_0.vpp comparator_0.vnn avdd.t184 avdd.t177 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X985 dvss.t164 otrip_decoded[5].t0 a_n3895_n1230# dvss.t163 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X986 comparator_0.vpp vbg_1v2.t28 comparator_0.vt comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X987 por.t19 sky130_fd_sc_hd__inv_4_4.Y dvdd.t249 dvdd.t248 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X988 avdd.t503 a_6765_n1142# a_7458_n2256# avdd.t502 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.1365 ps=1.49 w=0.42 l=1
X989 a_6765_n2876# a_6665_n2964# dvss.t389 dvss.t388 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X990 comparator_1.vnn avss.t436 comparator_1.vt comparator_1.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=8
X991 por.t4 sky130_fd_sc_hd__inv_4_4.Y dvss.t658 dvss.t657 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X992 a_697_n2212# a_329_n1230# dvss.t418 dvss.t417 sky130_fd_pr__nfet_01v8 ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X993 avdd.t635 comparator_1.vpp comparator_1.vnn avdd.t80 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X994 comparator_1.vnn avss.t437 comparator_1.vt comparator_1.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=8
X995 a_1122_n3990# a_697_n3946# dvss.t487 dvss.t486 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X996 a_n26074_n2937# a_n25696_n10337# avss.t0 sky130_fd_pr__res_xhigh_po_1p41 l=35
X997 avdd.t268 avdd.t267 avdd.t268 avdd.t240 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=8
X998 dvdd.t65 schmitt_trigger_0.out.t13 sky130_fd_sc_hd__inv_4_0.Y dvdd.t64 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X999 dvss.t130 a_8777_n2964# a_8877_n2876# dvss.t129 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X1000 dvss.t686 a_n7751_n3946# a_n7326_n3990# dvss.t685 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X1001 sky130_fd_sc_hvl__inv_4_0.A sky130_fd_sc_hvl__inv_1_0.A avdd.t591 avdd.t590 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X1002 a_n11219_9395# a_n11597_1995# avss.t234 sky130_fd_pr__res_xhigh_po_1p41 l=35
X1003 dcomp.t6 sky130_fd_sc_hd__inv_4_3.Y dvss.t740 dvss.t739 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1004 avss.t28 comparator_1.n1 dcomp3v3 avss.t27 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X1005 rstring_mux_0.vtrip_decoded_b_avdd[7] rstring_mux_0.vtrip_decoded_avdd[7] avdd.t409 avdd.t408 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X1006 a_n12731_9395# a_n12353_1995# avss.t409 sky130_fd_pr__res_xhigh_po_1p41 l=35
X1007 a_429_n1142# a_329_n1230# dvss.t416 dvss.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X1008 a_3234_n2256# a_2809_n2212# dvss.t326 dvss.t325 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X1009 a_n25318_n2937# a_n24940_n10337# avss.t0 sky130_fd_pr__res_xhigh_po_1p41 l=35
X1010 avdd.t134 a_8877_n2876# a_10084_n3212# avdd.t133 sky130_fd_pr__pfet_g5v0d10v5 ad=0.24375 pd=1.825 as=0.3975 ps=3.53 w=1.5 l=0.5
X1011 avdd.t601 comparator_0.vpp comparator_0.vnn avdd.t182 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1012 avdd.t266 avdd.t265 avdd.t266 avdd.t234 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=8
X1013 rstring_mux_0.vtrip_decoded_avdd[6] a_7972_n3212# dvss.t629 dvss.t628 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.121875 ps=1.075 w=0.75 l=0.5
X1014 vin rstring_mux_0.otrip_decoded_b_avdd[5] rstring_mux_0.vtrip5.t1 avdd.t157 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X1015 sky130_fd_sc_hd__inv_4_1.A por_unbuf.t11 dvss.t549 dvss.t548 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1016 dvss.t1 otrip_decoded[3].t0 a_n6007_n1230# dvss.t0 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X1017 a_8877_n2876# a_8777_n2964# dvss.t128 dvss.t127 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X1018 osc_ck.t5 rc_osc_0.n.t11 dvdd.t181 dvdd.t180 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X1019 avss.t335 ibias_gen_0.isrc_sel ibias_gen_0.vn0.t4 avss.t334 sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=2
X1020 dvdd.t290 sky130_fd_sc_hd__inv_4_3.Y dcomp.t20 dvdd.t289 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1021 pwup_filt.t21 sky130_fd_sc_hd__inv_4_0.Y dvdd.t21 dvdd.t20 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1022 dvss.t217 a_4921_n2212# a_5346_n2256# dvss.t216 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X1023 avss.t333 ibias_gen_0.isrc_sel ibias_gen_0.isrc_sel_b avss.t332 sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=1
X1024 pwup_filt.t3 sky130_fd_sc_hd__inv_4_0.Y dvss.t64 dvss.t63 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1025 a_n1415_n3946# a_n1783_n2964# dvdd.t119 dvdd.t118 sky130_fd_pr__pfet_01v8_hvt ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X1026 a_3234_n3990# a_2809_n3946# dvss.t442 dvss.t441 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X1027 a_7691_n11914# a_7313_n19314# avss.t62 sky130_fd_pr__res_xhigh_po_1p41 l=35
X1028 avdd.t600 comparator_0.vpp comparator_0.vnn avdd.t182 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1029 comparator_1.vpp comparator_1.vpp avdd.t634 avdd.t63 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1030 a_n22294_n2937# a_n22672_n10337# avss.t0 sky130_fd_pr__res_xhigh_po_1p41 l=35
X1031 a_5346_n2256# a_4921_n2212# dvss.t215 dvss.t214 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X1032 comparator_1.vnn comparator_1.vpp avdd.t633 avdd.t73 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1033 ibias_gen_0.vp1.t10 ibias_gen_0.isrc_sel_b ibias_gen_0.vp.t2 avdd.t488 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X1034 avdd.t463 rstring_mux_0.ena_b rstring_mux_0.vtop.t5 avdd.t462 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X1035 dvss.t323 otrip_decoded[1].t0 a_n8119_n1230# dvss.t322 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X1036 comparator_1.vt vin comparator_1.vpp comparator_1.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1037 dvdd.t7 force_pdnb.t1 a_8777_n2964# dvdd.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X1038 dvss.t286 dvss.t284 rc_osc_0.m dvss.t285 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X1039 a_n24562_n2937# a_n24940_n10337# avss.t0 sky130_fd_pr__res_xhigh_po_1p41 l=35
X1040 a_n21538_n2937# a_n21916_n10337# avss.t0 sky130_fd_pr__res_xhigh_po_1p41 l=35
X1041 dvss.t229 a_7033_n2212# a_7458_n2256# dvss.t228 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X1042 dvdd.t183 rc_osc_0.n.t12 rc_osc_0.m dvdd.t182 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1043 comparator_1.vpp vin comparator_1.vt comparator_1.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1044 a_n3527_n3946# a_n3895_n2964# dvdd.t129 dvdd.t128 sky130_fd_pr__pfet_01v8_hvt ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X1045 comparator_0.vnn avss.t438 comparator_0.vt comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=8
X1046 ibias_gen_0.vstart.t3 vbg_1v2.t29 ibias_gen_0.vn0.t11 avss.t130 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X1047 avss.t399 ibias_gen_0.vn1.t0 ibias_gen_0.vn1.t1 avss.t120 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=8
X1048 rstring_mux_0.otrip_decoded_avdd[6] a_n476_n3212# dvss.t192 dvss.t191 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.121875 ps=1.075 w=0.75 l=0.5
X1049 avdd.t145 a_n1683_n2876# a_n990_n3990# avdd.t144 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.1365 ps=1.49 w=0.42 l=1
X1050 vin rstring_mux_0.otrip_decoded_b_avdd[7] rstring_mux_0.vtrip7.t1 avdd.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X1051 comparator_1.vpp vin comparator_1.vt comparator_1.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1052 por.t3 sky130_fd_sc_hd__inv_4_4.Y dvss.t656 dvss.t655 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1053 a_n10279_n24979# a_12321_n24601# dvss.t400 sky130_fd_pr__res_xhigh_po_1p41 l=111
X1054 avdd.t69 comparator_1.vnn comparator_1.vpp avdd.t65 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1055 avss.t172 avss.t170 avss.t172 avss.t171 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=8
X1056 a_n23806_n2937# a_n24184_n10337# avss.t0 sky130_fd_pr__res_xhigh_po_1p41 l=35
X1057 avss.t317 ibias_gen_0.ena_b ibias_gen_0.vn1.t8 avss.t316 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X1058 a_2809_n2212# a_2441_n1230# dvdd.t9 dvdd.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X1059 dvss.t345 a_n1783_n2964# a_n1683_n2876# dvss.t344 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X1060 comparator_0.vpp vbg_1v2.t30 comparator_0.vt comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1061 porb.t3 sky130_fd_sc_hd__inv_4_1.Y dvss.t497 dvss.t496 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1062 a_7458_n2256# a_7033_n2212# dvss.t227 dvss.t226 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X1063 rstring_mux_0.ena a_10084_n3212# avdd.t130 avdd.t129 sky130_fd_pr__pfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.24375 ps=1.825 w=1.5 l=0.5
X1064 rc_osc_0.vr a_12321_n22333# dvss.t34 sky130_fd_pr__res_xhigh_po_1p41 l=111
X1065 avdd.t461 rstring_mux_0.ena_b rstring_mux_0.vtop.t4 avdd.t460 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X1066 dcomp3v3 comparator_1.n1 avss.t26 avss.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X1067 dvdd.t205 por_unbuf.t12 sky130_fd_sc_hd__inv_4_1.A dvdd.t204 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1068 rstring_mux_0.vtrip_decoded_b_avdd[5] rstring_mux_0.vtrip_decoded_avdd[5] avss.t246 avss.t245 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X1069 comparator_1.vpp comparator_1.vpp avdd.t632 avdd.t63 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1070 sky130_fd_sc_hd__inv_4_4.Y por_unbuf.t13 dvss.t551 dvss.t550 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1071 vin rstring_mux_0.otrip_decoded_b_avdd[0] rstring_mux_0.vtrip0.t0 avdd.t139 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X1072 comparator_0.vm comparator_0.vm avss.t90 avss.t88 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1073 avss.t169 avss.t168 ibias_gen_0.ve.t1 sky130_fd_pr__pnp_05v5_W0p68L0p68
**devattr s=18496,544 d=4547244,10712
X1074 ibias_gen_0.isrc_sel a_10084_n1478# dvss.t340 dvss.t175 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.121875 ps=1.075 w=0.75 l=0.5
X1075 comparator_0.vt comparator_0.vinn.t61 comparator_0.vnn comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1076 comparator_1.vnn comparator_1.vpp avdd.t631 avdd.t73 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1077 avss.t167 avss.t166 avss.t167 avss.t136 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=8
X1078 dvss.t738 sky130_fd_sc_hd__inv_4_3.Y dcomp.t5 dvss.t737 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1079 dvdd.t77 schmitt_trigger_0.in.t9 schmitt_trigger_0.m.t8 dvdd.t76 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X1080 dvss.t25 a_9145_n2212# a_9570_n2256# dvss.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X1081 a_n1683_n2876# a_n1783_n2964# dvss.t343 dvss.t342 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X1082 avss.t349 sky130_fd_sc_hvl__inv_16_0.A porb_h.t3 avss.t348 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X1083 ibias_gen_0.ve.t0 avss.t164 avss.t165 avss.t67 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=4
X1084 schmitt_trigger_0.m.t7 schmitt_trigger_0.in.t10 dvdd.t79 dvdd.t78 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X1085 rstring_mux_0.otrip_decoded_avdd[3] a_n4700_n1478# avdd.t449 avdd.t438 sky130_fd_pr__pfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.24375 ps=1.825 w=1.5 l=0.5
X1086 a_n5639_n3946# a_n6007_n2964# dvdd.t125 dvdd.t124 sky130_fd_pr__pfet_01v8_hvt ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X1087 avdd.t52 comparator_0.n1 dcomp3v3uv avdd.t51 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X1088 dvss.t160 schmitt_trigger_0.out.t14 sky130_fd_sc_hd__inv_4_0.Y dvss.t159 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1089 a_9570_n3990# a_9145_n3946# dvss.t642 dvss.t641 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X1090 dvdd.t147 sky130_fd_sc_hd__inv_4_1.Y porb.t19 dvdd.t146 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1091 a_7033_n2212# a_6665_n1230# dvdd.t221 dvdd.t220 sky130_fd_pr__pfet_01v8_hvt ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X1092 dvss.t426 a_2441_n2964# a_2541_n2876# dvss.t425 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X1093 dvss.t17 a_n1415_n3946# a_n990_n3990# dvss.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X1094 a_n8185_n11914# a_n8563_n19314# avss.t235 sky130_fd_pr__res_xhigh_po_1p41 l=35
X1095 dvss.t404 a_n3895_n2964# a_n3795_n2876# dvss.t403 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X1096 rstring_mux_0.vtrip6.t1 rstring_mux_0.vtrip_decoded_b_avdd[6] comparator_0.vinn.t5 avdd.t93 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X1097 porb_h.t2 sky130_fd_sc_hvl__inv_16_0.A avss.t347 avss.t346 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X1098 ibias_gen_0.vp1.t6 ibias_gen_0.vn1.t16 avss.t126 avss.t117 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=8
X1099 sky130_fd_sc_hd__inv_4_1.Y sky130_fd_sc_hd__inv_4_1.A dvdd.t225 dvdd.t224 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1100 dvss.t56 a_n3795_n1142# a_n2588_n1478# dvss.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0.121875 pd=1.075 as=0.19875 ps=2.03 w=0.75 l=0.5
X1101 avss.t127 ibias_gen_0.vn1.t17 ibias_gen_0.vp1.t7 avss.t120 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=8
X1102 dvdd.t19 sky130_fd_sc_hd__inv_4_0.Y pwup_filt.t20 dvdd.t18 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1103 dvdd.t71 otrip_decoded[7].t1 a_n1783_n1230# dvdd.t70 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X1104 comparator_0.vnn comparator_0.vpp avdd.t599 avdd.t186 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1105 avdd.t183 comparator_0.vnn comparator_0.vnn avdd.t182 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1106 a_n3510_6789# a_n3878_7771# dvss.t525 dvss.t524 sky130_fd_pr__nfet_01v8 ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X1107 a_n20782_n2937# a_n20404_n10337# avss.t0 sky130_fd_pr__res_xhigh_po_1p41 l=35
X1108 dvss.t254 a_10515_n2156# a_10874_n2222# dvss.t252 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.105 ps=1.03 w=0.75 l=0.5
X1109 rc_osc_0.m rc_osc_0.in dvdd.t211 dvdd.t210 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.1475 ps=1.295 w=1 l=0.5
X1110 a_n5214_n3990# a_n5639_n3946# dvss.t146 dvss.t145 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X1111 avdd.t264 avdd.t263 avdd.t264 avdd.t234 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=8
X1112 a_n3102_n3990# a_n3527_n3946# dvss.t472 dvss.t471 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X1113 a_n990_n3990# a_n1415_n3946# dvss.t15 dvss.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X1114 comparator_0.vinn.t29 avdd.t261 comparator_0.vinn.t29 avdd.t262 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=0.6
X1115 avss.t85 sky130_fd_sc_hvl__inv_4_0.A sky130_fd_sc_hvl__inv_16_0.A avss.t84 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X1116 pwup_filt.t2 sky130_fd_sc_hd__inv_4_0.Y dvss.t62 dvss.t61 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1117 rstring_mux_0.vtrip1.t8 rstring_mux_0.otrip_decoded_avdd[1] vin avss.t298 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X1118 rstring_mux_0.otrip_decoded_avdd[1] a_n6812_n1478# avdd.t11 avdd.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.24375 ps=1.825 w=1.5 l=0.5
X1119 rstring_mux_0.vtrip1.t3 rstring_mux_0.vtrip0.t2 avss.t236 sky130_fd_pr__res_xhigh_po_1p41 l=35
X1120 porb_h.t20 sky130_fd_sc_hvl__inv_16_0.A avdd.t547 avdd.t546 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X1121 dcomp.t19 sky130_fd_sc_hd__inv_4_3.Y dvdd.t288 dvdd.t287 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1122 dvss.t121 a_10515_n1026# a_10874_n1026# dvss.t119 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X1123 a_n7326_n2256# a_n7751_n2212# dvss.t458 dvss.t457 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X1124 dvss.t225 a_n1683_n2876# a_n476_n3212# dvss.t224 sky130_fd_pr__nfet_g5v0d10v5 ad=0.121875 pd=1.075 as=0.19875 ps=2.03 w=0.75 l=0.5
X1125 por.t18 sky130_fd_sc_hd__inv_4_4.Y dvdd.t247 dvdd.t246 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1126 a_10874_n2222# a_10515_n2156# dvss.t253 dvss.t252 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.178875 ps=1.26 w=0.75 l=0.5
X1127 avdd.t260 avdd.t257 avdd.t259 avdd.t258 sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.58 as=0 ps=0 w=5 l=4
X1128 a_9145_n2212# a_8777_n1230# dvdd.t84 dvdd.t83 sky130_fd_pr__pfet_01v8_hvt ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X1129 dvss.t375 a_n6007_n2964# a_n5907_n2876# dvss.t374 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X1130 a_n3649_n11914# rstring_mux_0.vtrip0.t3 avss.t275 sky130_fd_pr__res_xhigh_po_1p41 l=35
X1131 avdd.t459 rstring_mux_0.ena_b rstring_mux_0.vtop.t3 avdd.t458 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X1132 sky130_fd_sc_hd__inv_4_3.Y vl dvdd.t237 dvdd.t236 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1133 dvdd.t5 otrip_decoded[5].t1 a_n3895_n1230# dvdd.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X1134 avdd.t545 sky130_fd_sc_hvl__inv_16_0.A porb_h.t19 avdd.t544 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X1135 comparator_1.vt comparator_1.vn avss.t292 avss.t280 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1136 a_10874_n1026# a_10515_n1026# dvss.t120 dvss.t119 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.178875 ps=1.26 w=0.75 l=0.5
X1137 a_n7326_n3990# a_n7751_n3946# dvss.t684 dvss.t683 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X1138 avdd.t256 avdd.t254 avdd.t255 avdd.t221 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=8
X1139 a_697_n2212# a_329_n1230# dvdd.t131 dvdd.t130 sky130_fd_pr__pfet_01v8_hvt ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X1140 a_n8019_n2876# a_n8119_n2964# dvss.t698 dvss.t697 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X1141 dvdd.t103 dvss.t776 a_4553_n2964# dvdd.t102 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X1142 avdd.t435 ibias_gen_0.vp.t12 comparator_0.ibias avdd.t434 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X1143 porb.t2 sky130_fd_sc_hd__inv_4_1.Y dvss.t495 dvss.t494 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1144 comparator_0.vnn comparator_0.vpp avdd.t598 avdd.t186 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1145 avdd.t597 comparator_0.vpp comparator_0.vpp avdd.t179 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1146 comparator_1.vnn vbg_1v2.t31 comparator_1.vt comparator_1.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1147 dcomp.t18 sky130_fd_sc_hd__inv_4_3.Y dvdd.t286 dvdd.t285 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1148 a_1122_n3990# a_697_n3946# dvss.t485 dvss.t484 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X1149 comparator_0.vinn.t1 rstring_mux_0.vtrip_decoded_avdd[1] rstring_mux_0.vtrip1.t0 avss.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X1150 ibg_200n rstring_mux_0.ena a_n15479_n3901# avss.t324 sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=0.6
X1151 avdd.t132 a_8877_n2876# a_9570_n3990# avdd.t131 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.1365 ps=1.49 w=0.42 l=1
X1152 a_4921_n3946# a_4553_n2964# dvdd.t89 dvdd.t88 sky130_fd_pr__pfet_01v8_hvt ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X1153 dcomp3v3uv comparator_0.n1 avss.t47 avss.t46 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X1154 avdd.t457 rstring_mux_0.ena_b rstring_mux_0.vtop.t2 avdd.t456 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X1155 avdd.t68 comparator_1.vnn comparator_1.vpp avdd.t65 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1156 comparator_1.vpp vin comparator_1.vt comparator_1.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1157 a_n16775_n2223# ibias_gen_0.ena_b ibias_gen_0.vstart.t0 avdd.t506 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=0.6
X1158 comparator_0.vinn.t21 rstring_mux_0.vtrip_decoded_b_avdd[1] rstring_mux_0.vtrip1.t5 avdd.t176 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X1159 avdd.t405 ibias_gen_0.vp0.t12 ibias_gen_0.vn0.t1 avdd.t404 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X1160 dvss.t440 a_2809_n3946# a_3234_n3990# dvss.t439 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X1161 comparator_1.vpp comparator_1.vnn avdd.t67 avdd.t63 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1162 avdd.t21 comparator_1.n1 dcomp3v3 avdd.t20 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X1163 dvss.t493 sky130_fd_sc_hd__inv_4_1.Y porb.t1 dvss.t492 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1164 dvdd.t3 otrip_decoded[3].t1 a_n6007_n1230# dvdd.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X1165 dvss.t483 a_697_n3946# a_1122_n3990# dvss.t482 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X1166 ibias_gen_0.ve.t3 ibias_gen_0.vn0.t7 ibias_gen_0.vn0.t8 avss.t67 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X1167 dvdd.t101 dvss.t777 a_6665_n2964# dvdd.t100 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X1168 rstring_mux_0.vtrip3.t4 rstring_mux_0.otrip_decoded_b_avdd[3] vin avdd.t172 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X1169 a_2399_n11914# a_2021_n19314# avss.t61 sky130_fd_pr__res_xhigh_po_1p41 l=35
X1170 a_n6673_n11914# a_n7051_n19314# avss.t240 sky130_fd_pr__res_xhigh_po_1p41 l=35
X1171 avdd.t66 comparator_1.vnn comparator_1.vpp avdd.t65 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1172 avss.t345 sky130_fd_sc_hvl__inv_16_0.A porb_h.t1 avss.t344 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X1173 comparator_0.vinn.t42 rstring_mux_0.vtrip_decoded_avdd[0] rstring_mux_0.vtrip0.t8 avss.t374 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X1174 comparator_1.vnn comparator_1.vpp avdd.t630 avdd.t73 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1175 por.t2 sky130_fd_sc_hd__inv_4_4.Y dvss.t654 dvss.t653 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1176 a_n7429_n11914# a_n7051_n19314# avss.t11 sky130_fd_pr__res_xhigh_po_1p41 l=35
X1177 a_n10453_n11914# a_n10075_n19314# avss.t12 sky130_fd_pr__res_xhigh_po_1p41 l=35
X1178 a_3234_n3990# a_2809_n3946# dvss.t438 dvss.t437 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X1179 dvss.t736 sky130_fd_sc_hd__inv_4_3.Y dcomp.t4 dvss.t735 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1180 rc_osc_0.in dvss.t572 sky130_fd_pr__cap_mim_m3_2 l=30 w=30
X1181 avdd.t253 avdd.t251 avdd.t252 avdd.t221 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=8
X1182 ibias_gen_0.vn0.t10 vbg_1v2.t32 ibias_gen_0.vstart.t2 avss.t131 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X1183 rc_osc_0.n.t0 rc_osc_0.m dvss.t112 dvss.t111 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X1184 avdd.t629 comparator_1.vpp comparator_1.n0 avdd.t80 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1185 rstring_mux_0.vtrip_decoded_avdd[7] a_7972_n1478# avdd.t102 avdd.t101 sky130_fd_pr__pfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.24375 ps=1.825 w=1.5 l=0.5
X1186 dvdd.t1 otrip_decoded[1].t1 a_n8119_n1230# dvdd.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X1187 dvss.t106 a_4921_n3946# a_5346_n3990# dvss.t105 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X1188 comparator_0.vnn avss.t439 comparator_0.vt comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=8
X1189 a_n12731_9395# a_n13109_1995# avss.t401 sky130_fd_pr__res_xhigh_po_1p41 l=35
X1190 avdd.t596 comparator_0.vpp comparator_0.vpp avdd.t179 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1191 avdd.t543 sky130_fd_sc_hvl__inv_16_0.A porb_h.t18 avdd.t542 sky130_fd_pr__pfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X1192 dvdd.t145 sky130_fd_sc_hd__inv_4_1.Y porb.t18 dvdd.t144 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1193 avdd.t250 avdd.t249 avdd.t250 avdd.t240 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=8
X1194 dvdd.t207 por_unbuf.t14 sky130_fd_sc_hd__inv_4_4.Y dvdd.t206 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1195 schmitt_trigger_0.in.t11 dvss.t171 sky130_fd_pr__cap_mim_m3_2 l=30 w=30
X1196 comparator_0.vpp vbg_1v2.t33 comparator_0.vt comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1197 dvdd.t17 sky130_fd_sc_hd__inv_4_0.Y pwup_filt.t19 dvdd.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1198 sky130_fd_sc_hd__inv_4_1.Y sky130_fd_sc_hd__inv_4_1.A dvdd.t223 dvdd.t222 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1199 rstring_mux_0.vtrip6.t7 rstring_mux_0.otrip_decoded_avdd[6] vin avss.t308 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X1200 avdd.t455 rstring_mux_0.ena_b rstring_mux_0.vtop.t1 avdd.t454 sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=0.6
X1201 dvdd.t67 a_10874_n1026# a_10874_n2222# dvdd.t66 sky130_fd_pr__pfet_01v8_hvt ad=0.2968 pd=2.77 as=0.2968 ps=2.77 w=1.12 l=0.15
X1202 porb_h.t17 sky130_fd_sc_hvl__inv_16_0.A avdd.t541 avdd.t540 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X1203 dvss.t560 a_429_n1142# a_1636_n1478# dvss.t175 sky130_fd_pr__nfet_g5v0d10v5 ad=0.121875 pd=1.075 as=0.19875 ps=2.03 w=0.75 l=0.5
X1204 avdd.t1 a_n5907_n2876# a_n5214_n3990# avdd.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.1365 ps=1.49 w=0.42 l=1
X1205 vin avdd.t247 vin avdd.t248 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=0.6
X1206 dvss.t553 por_unbuf.t15 a_n3878_7771# dvss.t552 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X1207 rstring_mux_0.otrip_decoded_avdd[4] a_n2588_n3212# dvss.t767 dvss.t766 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.121875 ps=1.075 w=0.75 l=0.5
X1208 a_5346_n3990# a_4921_n3946# dvss.t104 dvss.t103 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X1209 dvss.t562 a_10514_n2760# a_10514_n3890# dvss.t561 sky130_fd_pr__nfet_g5v0d10v5 ad=0.178875 pd=1.26 as=0.1197 ps=1.41 w=0.42 l=0.5
X1210 rstring_mux_0.otrip_decoded_b_avdd[3] rstring_mux_0.otrip_decoded_avdd[3] avdd.t219 avdd.t218 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X1211 rstring_mux_0.vtrip_decoded_b_avdd[0] rstring_mux_0.vtrip_decoded_avdd[0] avdd.t573 avdd.t572 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X1212 dvdd.t209 rc_osc_0.in rc_osc_0.m dvdd.t208 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X1213 dvss.t734 sky130_fd_sc_hd__inv_4_3.Y dcomp.t3 dvss.t733 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1214 ibias_gen_0.vn1.t6 ibias_gen_0.isrc_sel_b avss.t304 avss.t303 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=2
X1215 avss.t163 avss.t162 avss.t163 avss.t136 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=8
X1216 dcomp.t17 sky130_fd_sc_hd__inv_4_3.Y dvdd.t284 dvdd.t283 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1217 dvss.t118 a_10515_n1026# a_10874_n1026# dvss.t117 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.19875 ps=2.03 w=0.75 l=0.5
X1218 avdd.t514 rstring_mux_0.ena rstring_mux_0.ena_b avdd.t513 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X1219 osc_ck.t6 rc_osc_0.n.t13 dvdd.t185 dvdd.t184 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X1220 vin avss.t160 vin avss.t161 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=0.6
X1221 por.t17 sky130_fd_sc_hd__inv_4_4.Y dvdd.t245 dvdd.t244 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1222 por.t1 sky130_fd_sc_hd__inv_4_4.Y dvss.t652 dvss.t651 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1223 dvss.t712 a_7033_n3946# a_7458_n3990# dvss.t711 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X1224 a_6179_n11914# a_5801_n19314# avss.t404 sky130_fd_pr__res_xhigh_po_1p41 l=35
X1225 a_n13477_n11914# a_n13855_n19314# avss.t259 sky130_fd_pr__res_xhigh_po_1p41 l=35
X1226 rstring_mux_0.otrip_decoded_avdd[1] a_n6812_n1478# dvss.t54 dvss.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.121875 ps=1.075 w=0.75 l=0.5
X1227 avdd.t246 avdd.t244 avdd.t245 avdd.t221 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=8
X1228 comparator_0.vinn.t28 avdd.t242 comparator_0.vinn.t28 avdd.t243 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=0.6
X1229 a_n8195_9395# a_n8573_1995# avss.t406 sky130_fd_pr__res_xhigh_po_1p41 l=35
X1230 dvss.t555 por_unbuf.t16 sky130_fd_sc_hd__inv_4_1.A dvss.t554 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1231 rstring_mux_0.vtrip_decoded_b_avdd[4] rstring_mux_0.vtrip_decoded_avdd[4] avdd.t17 avdd.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X1232 comparator_0.vm comparator_0.ena_b avss.t108 avss.t88 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X1233 comparator_0.vinn.t12 avss.t158 vin avss.t159 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X1234 sky130_fd_sc_hd__inv_4_3.Y vl dvdd.t235 dvdd.t234 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1235 dvdd.t15 sky130_fd_sc_hd__inv_4_0.Y pwup_filt.t18 dvdd.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1236 avdd.t595 comparator_0.vpp comparator_0.vpp avdd.t179 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1237 rstring_mux_0.otrip_decoded_avdd[7] a_n476_n1478# avdd.t148 avdd.t147 sky130_fd_pr__pfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.24375 ps=1.825 w=1.5 l=0.5
X1238 comparator_0.vt vbg_1v2.t34 comparator_0.vpp comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1239 comparator_0.n0 comparator_0.vm avss.t89 avss.t88 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1240 avdd.t241 avdd.t239 avdd.t241 avdd.t240 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=8
X1241 vin avss.t156 vin avss.t157 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=0.6
X1242 comparator_1.vnn vbg_1v2.t35 comparator_1.vt comparator_1.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1243 avdd.t657 a_n8019_n2876# a_n7326_n3990# avdd.t656 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.1365 ps=1.49 w=0.42 l=1
X1244 pwup_filt.t1 sky130_fd_sc_hd__inv_4_0.Y dvss.t60 dvss.t59 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1245 a_2809_n3946# a_2441_n2964# dvss.t424 dvss.t423 sky130_fd_pr__nfet_01v8 ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X1246 avss.t155 avss.t153 avss.t154 avss.t109 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=8
X1247 dvss.t732 sky130_fd_sc_hd__inv_4_3.Y dcomp.t2 dvss.t731 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1248 dvss.t470 a_n3527_n3946# a_n3102_n3990# dvss.t469 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X1249 avss.t272 comparator_0.n0 comparator_0.n1 avss.t271 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X1250 vin avss.t151 vin avss.t152 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=0.6
X1251 sky130_fd_sc_hvl__inv_16_0.A sky130_fd_sc_hvl__inv_4_0.A avss.t83 avss.t82 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X1252 comparator_1.vnn vbg_1v2.t36 comparator_1.vt comparator_1.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1253 a_n3778_7859# a_n3878_7771# dvss.t523 dvss.t522 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X1254 avss.t390 comparator_0.vn comparator_0.vn avss.t109 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1255 ibg_200n ibias_gen_0.ena_b a_n15529_n2223# avdd.t505 sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=0.6
X1256 porb_h.t0 sky130_fd_sc_hvl__inv_16_0.A avss.t343 avss.t342 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X1257 dvss.t640 a_9145_n3946# a_9570_n3990# dvss.t639 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X1258 a_887_n11914# a_1265_n19314# avss.t262 sky130_fd_pr__res_xhigh_po_1p41 l=35
X1259 avdd.t50 comparator_0.n1 dcomp3v3uv avdd.t49 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X1260 comparator_1.vt avss.t440 comparator_1.vnn comparator_1.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=8
X1261 a_n3102_n3990# a_n3527_n3946# dvss.t468 dvss.t467 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X1262 a_n10279_n23467# a_12321_n23089# dvss.t769 sky130_fd_pr__res_xhigh_po_1p41 l=111
X1263 avss.t81 sky130_fd_sc_hvl__inv_4_0.A sky130_fd_sc_hvl__inv_16_0.A avss.t80 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.105 ps=1.03 w=0.75 l=0.5
X1264 dvdd.t13 sky130_fd_sc_hd__inv_4_0.Y pwup_filt.t17 dvdd.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1265 rstring_mux_0.vtrip3.t1 rstring_mux_0.vtrip_decoded_avdd[3] comparator_0.vinn.t6 avss.t72 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X1266 dvss.t491 sky130_fd_sc_hd__inv_4_1.Y porb.t0 dvss.t490 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1267 avdd.t238 avdd.t236 avdd.t237 avdd.t230 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=8
X1268 dvss.t248 a_n3795_n2876# a_n2588_n3212# dvss.t247 sky130_fd_pr__nfet_g5v0d10v5 ad=0.121875 pd=1.075 as=0.19875 ps=2.03 w=0.75 l=0.5
X1269 a_7033_n3946# a_6665_n2964# dvss.t387 dvss.t386 sky130_fd_pr__nfet_01v8 ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X1270 dvss.t144 a_n5639_n3946# a_n5214_n3990# dvss.t143 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X1271 schmitt_trigger_0.in.t12 dvss.t172 sky130_fd_pr__cap_mim_m3_2 l=30 w=30
X1272 sky130_fd_sc_hvl__inv_1_0.A a_n2571_7523# avdd.t581 avdd.t163 sky130_fd_pr__pfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.24375 ps=1.825 w=1.5 l=0.5
X1273 dvss.t268 a_4553_n2964# a_4653_n2876# dvss.t267 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X1274 rstring_mux_0.vtrip6.t3 rstring_mux_0.vtrip_decoded_avdd[6] comparator_0.vinn.t8 avss.t93 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X1275 dvss.t152 otrip_decoded[6].t1 a_n1783_n2964# dvss.t151 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X1276 comparator_1.vt vbg_1v2.t37 comparator_1.vnn comparator_1.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1277 comparator_0.vnn avss.t441 comparator_0.vt comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=8
X1278 avdd.t539 sky130_fd_sc_hvl__inv_16_0.A porb_h.t16 avdd.t538 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X1279 comparator_1.vt vbg_1v2.t38 comparator_1.vnn comparator_1.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1280 dvss.t557 por_unbuf.t17 sky130_fd_sc_hd__inv_4_4.Y dvss.t556 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1281 comparator_0.vnn comparator_0.vinn.t62 comparator_0.vt comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1282 rstring_mux_0.vtrip1.t4 rstring_mux_0.vtrip_decoded_b_avdd[1] comparator_0.vinn.t20 avdd.t175 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X1283 comparator_1.vpp comparator_1.vnn avdd.t64 avdd.t63 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1284 dcomp3v3uv comparator_0.n1 avss.t45 avss.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X1285 comparator_0.vpp comparator_0.vnn avdd.t181 avdd.t177 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1286 comparator_1.vpp vin comparator_1.vt comparator_1.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1287 a_n5214_n3990# a_n5639_n3946# dvss.t142 dvss.t141 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X1288 schmitt_trigger_0.in.t13 dvss.t173 sky130_fd_pr__cap_mim_m3_2 l=30 w=30
X1289 comparator_0.vpp vbg_1v2.t39 comparator_0.vt comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1290 comparator_0.vnn avss.t442 comparator_0.vt comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=8
X1291 avdd.t510 a_n1683_n1142# a_n476_n1478# avdd.t147 sky130_fd_pr__pfet_g5v0d10v5 ad=0.24375 pd=1.825 as=0.3975 ps=3.53 w=1.5 l=0.5
X1292 rstring_mux_0.vtrip_decoded_b_avdd[2] rstring_mux_0.vtrip_decoded_avdd[2] avss.t379 avss.t378 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X1293 comparator_0.vpp vbg_1v2.t40 comparator_0.vt comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1294 dvdd.t243 sky130_fd_sc_hd__inv_4_4.Y por.t16 dvdd.t242 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1295 dvdd.t143 sky130_fd_sc_hd__inv_4_1.Y porb.t17 dvdd.t142 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1296 dvss.t13 a_n5907_n2876# a_n4700_n3212# dvss.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0.121875 pd=1.075 as=0.19875 ps=2.03 w=0.75 l=0.5
X1297 vin rstring_mux_0.otrip_decoded_b_avdd[3] rstring_mux_0.vtrip3.t3 avdd.t171 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X1298 a_4667_n11914# a_4289_n19314# avss.t237 sky130_fd_pr__res_xhigh_po_1p41 l=35
X1299 dvss.t283 dvss.t281 rc_osc_0.n.t4 dvss.t282 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X1300 a_1122_n3990# a_697_n3946# dvss.t481 dvss.t480 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X1301 a_9145_n3946# a_8777_n2964# dvss.t126 dvss.t125 sky130_fd_pr__nfet_01v8 ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X1302 a_n8941_n11914# a_n9319_n19314# avss.t239 sky130_fd_pr__res_xhigh_po_1p41 l=35
X1303 a_n11965_n11914# a_n12343_n19314# avss.t4 sky130_fd_pr__res_xhigh_po_1p41 l=35
X1304 comparator_1.n1 comparator_1.n0 avdd.t583 avdd.t582 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.6
X1305 avdd.t235 avdd.t233 avdd.t235 avdd.t234 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=8
X1306 avdd.t150 a_n990_n2256# a_n1683_n1142# avdd.t149 sky130_fd_pr__pfet_g5v0d10v5 ad=0.2142 pd=1.99 as=0.2142 ps=1.99 w=0.42 l=1
X1307 dvss.t682 a_n7751_n3946# a_n7326_n3990# dvss.t681 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X1308 comparator_0.vinn.t13 avss.t149 comparator_0.vinn.t13 avss.t150 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=0.6
X1309 avdd.t232 avdd.t229 avdd.t231 avdd.t230 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=8
X1310 avss.t279 comparator_1.vm comparator_1.vm avss.t278 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1311 ibias_gen_0.vn0.t2 ibias_gen_0.vp0.t13 avdd.t407 avdd.t406 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X1312 avss.t148 avss.t145 avss.t147 avss.t146 sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0 ps=0 w=5 l=8
X1313 a_4667_n11914# a_5045_n19314# avss.t257 sky130_fd_pr__res_xhigh_po_1p41 l=35
X1314 comparator_0.vnn comparator_0.vinn.t63 comparator_0.vt comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1315 por.t0 sky130_fd_sc_hd__inv_4_4.Y dvss.t650 dvss.t649 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1316 dvss.t762 otrip_decoded[4].t1 a_n3895_n2964# dvss.t761 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X1317 schmitt_trigger_0.in.t14 dvss.t174 sky130_fd_pr__cap_mim_m3_2 l=30 w=30
X1318 a_n12721_n11914# a_n12343_n19314# avss.t276 sky130_fd_pr__res_xhigh_po_1p41 l=35
X1319 ibias_gen_0.vr.t1 avss.t144 ibias_gen_0.ve.t2 avss.t67 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X1320 dvss.t730 sky130_fd_sc_hd__inv_4_3.Y dcomp.t1 dvss.t729 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1321 a_697_n3946# a_329_n2964# dvss.t92 dvss.t91 sky130_fd_pr__nfet_01v8 ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X1322 vin avss.t142 vin avss.t143 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=0.6
X1323 ibias_gen_0.vp0.t0 avss.t140 ibias_gen_0.vn0.t0 avss.t141 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X1324 rstring_mux_0.vtrip_decoded_avdd[4] a_5860_n3212# dvss.t590 dvss.t589 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.121875 ps=1.075 w=0.75 l=0.5
X1325 ibias_gen_0.vn1.t5 avdd.t227 ibias_gen_0.vp1.t9 avdd.t228 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X1326 dvss.t162 schmitt_trigger_0.out.t15 sky130_fd_sc_hd__inv_4_0.Y dvss.t161 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1327 dcomp3v3uv comparator_0.n1 avdd.t48 avdd.t47 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X1328 vin avss.t138 vin avss.t139 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=0.6
X1329 comparator_1.vt vin comparator_1.vpp comparator_1.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1330 avdd.t226 avdd.t224 avdd.t226 avdd.t225 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=4
X1331 avss.t137 avss.t135 avss.t137 avss.t136 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=8
X1332 dvdd.t141 sky130_fd_sc_hd__inv_4_1.Y porb.t16 dvdd.t140 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1333 dvss.t764 a_n8019_n2876# a_n6812_n3212# dvss.t763 sky130_fd_pr__nfet_g5v0d10v5 ad=0.121875 pd=1.075 as=0.19875 ps=2.03 w=0.75 l=0.5
X1334 avdd.t154 a_n3795_n2876# a_n3102_n3990# avdd.t153 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.1365 ps=1.49 w=0.42 l=1
X1335 a_10514_n2760# dcomp3v3uv avdd.t46 avdd.t45 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.1197 ps=1.41 w=0.42 l=0.5
X1336 avss.t134 avss.t133 avss.t134 avss.t88 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=8
X1337 avdd.t223 avdd.t220 avdd.t222 avdd.t221 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=8
X1338 dcomp3v3 comparator_1.n1 avdd.t19 avdd.t18 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X1339 dcomp.t16 sky130_fd_sc_hd__inv_4_3.Y dvdd.t282 dvdd.t281 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1340 dvdd.t11 sky130_fd_sc_hd__inv_4_0.Y pwup_filt.t16 dvdd.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1341 a_429_n2876# a_329_n2964# dvss.t90 dvss.t89 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X1342 a_3234_n3990# a_2809_n3946# dvss.t436 dvss.t435 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X1343 comparator_0.vt avss.t443 comparator_0.vnn comparator_0.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=8
X1344 avdd.t180 comparator_0.vnn comparator_0.vm avdd.t179 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1345 a_10874_n1026# a_10874_n2222# dvdd.t86 dvdd.t85 sky130_fd_pr__pfet_01v8_hvt ad=0.2968 pd=2.77 as=0.1568 ps=1.4 w=1.12 l=0.15
X1346 dvss.t140 otrip_decoded[2].t1 a_n6007_n2964# dvss.t139 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X1347 rstring_mux_0.otrip_decoded_b_avdd[6] rstring_mux_0.otrip_decoded_avdd[6] avss.t307 avss.t306 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X1348 ibias_gen_0.vstart.t1 vbg_1v2.t41 ibias_gen_0.vn0.t9 avss.t128 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X1349 pwup_filt.t0 sky130_fd_sc_hd__inv_4_0.Y dvss.t58 dvss.t57 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1350 dvdd.t139 osc_ena.t3 rc_osc_0.in dvdd.t138 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X1351 comparator_0.vpp comparator_0.vnn avdd.t178 avdd.t177 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1352 dvss.t728 sky130_fd_sc_hd__inv_4_3.Y dcomp.t0 dvss.t727 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1353 dvss.t102 a_4921_n3946# a_5346_n3990# dvss.t101 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X1354 schmitt_trigger_0.out.t0 schmitt_trigger_0.m.t17 dvss.t280 dvss.t279 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X1355 comparator_1.vt avss.t444 comparator_1.vnn comparator_1.vt sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=8
X1356 dvss.t399 a_429_n2876# a_1636_n3212# dvss.t398 sky130_fd_pr__nfet_g5v0d10v5 ad=0.121875 pd=1.075 as=0.19875 ps=2.03 w=0.75 l=0.5
R0 dvss.n995 dvss.n853 198880
R1 dvss.n837 dvss.n836 198880
R2 dvss.t255 dvss.n836 192115
R3 dvss.n995 dvss.t261 192115
R4 dvss.n4289 dvss.n4288 82533.9
R5 dvss.n2519 dvss.n2111 79031.1
R6 dvss.n4286 dvss.n4264 78608.8
R7 dvss.n4265 dvss.n4264 78608.8
R8 dvss.n4286 dvss.n4270 78608.8
R9 dvss.n4270 dvss.n4265 78608.8
R10 dvss.n2491 dvss.n2490 37915.2
R11 dvss.n2179 dvss.n2111 29969.5
R12 dvss.n2520 dvss.n103 22284.8
R13 dvss.n2180 dvss.n2179 16469.1
R14 dvss.n4267 dvss.n4249 12828.2
R15 dvss.n4290 dvss.n4249 12828.2
R16 dvss.n4267 dvss.n4263 12822.4
R17 dvss.n4290 dvss.n4263 12822.4
R18 dvss.n2574 dvss.n2573 12752.5
R19 dvss dvss.n2443 12161.8
R20 dvss.n4310 dvss.n58 8941.81
R21 dvss.n2442 dvss.n2308 8034.33
R22 dvss.n687 dvss.t717 8003.11
R23 dvss.n4187 dvss.t687 8003.11
R24 dvss.n4152 dvss.t149 8003.11
R25 dvss.t475 dvss.n3238 8003.11
R26 dvss.t22 dvss.n351 8003.11
R27 dvss.t480 dvss.n1946 8003.11
R28 dvss.n1681 dvss.t435 8003.11
R29 dvss.t109 dvss.n1389 8003.11
R30 dvss.n1162 dvss.t641 8003.11
R31 dvss.t713 dvss.t711 7626.67
R32 dvss.t719 dvss.t717 7626.67
R33 dvss.t683 dvss.t681 7626.67
R34 dvss.t685 dvss.t687 7626.67
R35 dvss.t145 dvss.t143 7626.67
R36 dvss.t147 dvss.t149 7626.67
R37 dvss.t471 dvss.t469 7626.67
R38 dvss.t475 dvss.t473 7626.67
R39 dvss.t18 dvss.t16 7626.67
R40 dvss.t22 dvss.t20 7626.67
R41 dvss.t484 dvss.t488 7626.67
R42 dvss.t480 dvss.t482 7626.67
R43 dvss.t437 dvss.t439 7626.67
R44 dvss.t443 dvss.t435 7626.67
R45 dvss.t103 dvss.t105 7626.67
R46 dvss.t109 dvss.t101 7626.67
R47 dvss.t643 dvss.t639 7626.67
R48 dvss.t647 dvss.t641 7626.67
R49 dvss.n1012 dvss.n1011 6912.63
R50 dvss.n3977 dvss.n3976 6332.05
R51 dvss.n3893 dvss.n249 6332.05
R52 dvss.n1989 dvss.n1924 6332.05
R53 dvss.n1964 dvss.n1930 6332.05
R54 dvss.n1936 dvss.n1935 6332.05
R55 dvss.n1762 dvss.n495 6332.05
R56 dvss.n1379 dvss.n1378 6332.05
R57 dvss.n1279 dvss.n615 6332.05
R58 dvss.n1460 dvss.t47 6153.5
R59 dvss.n3409 dvss.t47 6153.5
R60 dvss.n2222 dvss.t522 6153.5
R61 dvss.n4226 dvss.t619 6153.5
R62 dvss.n4066 dvss.t184 6153.5
R63 dvss.t47 dvss.n389 6153.5
R64 dvss.n1749 dvss.t47 6153.5
R65 dvss.n1266 dvss.t47 6153.5
R66 dvss.n2488 dvss.n2365 5792.85
R67 dvss.n4312 dvss.n4311 5772.37
R68 dvss.n4311 dvss.n4310 5605.26
R69 dvss.n2443 dvss.n2442 5502.51
R70 dvss.n1012 dvss.n838 5116.78
R71 dvss.n4285 dvss.n4271 5107.58
R72 dvss.n4283 dvss.n4271 5107.58
R73 dvss.n4285 dvss.n4284 5107.58
R74 dvss.n4284 dvss.n4283 5107.58
R75 dvss.n4226 dvss.n80 5082
R76 dvss.n4066 dvss.n4065 5082
R77 dvss.n3880 dvss.n259 5082
R78 dvss.n3881 dvss.n3880 5082
R79 dvss.n3185 dvss.n327 5082
R80 dvss.n1986 dvss.n327 5082
R81 dvss.n1961 dvss.n389 5082
R82 dvss.n3409 dvss.n3408 5082
R83 dvss.n1750 dvss.n1749 5082
R84 dvss.n1460 dvss.n1459 5082
R85 dvss.n1267 dvss.n1266 5082
R86 dvss.n2489 dvss.n2488 4826.37
R87 dvss.n2487 dvss.t516 4465.22
R88 dvss.n837 dvss.t257 4455
R89 dvss.t263 dvss.n853 4455
R90 dvss.n2369 dvss.n2366 4160.18
R91 dvss.n2440 dvss.n2366 4160.18
R92 dvss.n2369 dvss.n2367 4160.18
R93 dvss.n2440 dvss.n2367 4160.18
R94 dvss.n2234 dvss.n2233 4092
R95 dvss.n2491 dvss.n2308 3708.43
R96 dvss.n2574 dvss.n2111 3423.01
R97 dvss.n2488 dvss.n2487 3328.76
R98 dvss.n2575 dvss.n2574 3297.36
R99 dvss.n2180 dvss.t695 3216.06
R100 dvss.n2520 dvss.n2519 3196.46
R101 dvss.n2490 dvss.n2489 2962.09
R102 dvss dvss.n2308 2800
R103 dvss dvss.n2491 2763.24
R104 dvss.t257 dvss.t255 2310
R105 dvss.t261 dvss.t263 2310
R106 dvss.n1103 dvss.t252 2079.65
R107 dvss.n4289 dvss.t478 2014.07
R108 dvss.n2519 dvss.n2518 1808.4
R109 dvss.n2487 dvss.t85 1808.05
R110 dvss.t528 dvss.t526 1778.24
R111 dvss.t621 dvss.t615 1778.24
R112 dvss.t186 dvss.t178 1778.24
R113 dvss dvss.t159 1681.61
R114 dvss.n2234 dvss.t526 1652.85
R115 dvss.n4187 dvss.t621 1652.85
R116 dvss.t178 dvss.n4152 1652.85
R117 dvss.n4268 dvss.t534 1589.55
R118 dvss.n2489 dvss.t735 1395.12
R119 dvss.n2490 dvss.t673 1376.81
R120 dvss dvss.t632 1297.56
R121 dvss dvss.t556 1280.53
R122 dvss.n2442 dvss.n2441 1258.81
R123 dvss.t279 dvss.n2365 1124.77
R124 dvss.n2441 dvss.t165 1124.77
R125 dvss.t65 dvss.t85 1062.07
R126 dvss.t87 dvss.t65 1062.07
R127 dvss.t67 dvss.t87 1062.07
R128 dvss.t79 dvss.t67 1062.07
R129 dvss.t71 dvss.t79 1062.07
R130 dvss.t73 dvss.t71 1062.07
R131 dvss.t61 dvss.t73 1062.07
R132 dvss.t83 dvss.t61 1062.07
R133 dvss.t57 dvss.t83 1062.07
R134 dvss.t75 dvss.t57 1062.07
R135 dvss.t59 dvss.t77 1062.07
R136 dvss.t77 dvss.t69 1062.07
R137 dvss.t69 dvss.t81 1062.07
R138 dvss.t81 dvss.t63 1062.07
R139 dvss.t159 dvss.t155 1062.07
R140 dvss.t155 dvss.t161 1062.07
R141 dvss.t161 dvss.t153 1062.07
R142 dvss.t63 dvss 986.207
R143 dvss.t153 dvss 948.277
R144 dvss.t297 dvss.t279 920.795
R145 dvss.t157 dvss.t297 920.795
R146 dvss.t157 dvss.t167 920.795
R147 dvss.t167 dvss.t165 920.795
R148 dvss.n1052 dvss.t252 867.946
R149 dvss.n1091 dvss.t565 867.946
R150 dvss.n2443 dvss 847.126
R151 dvss.n4292 dvss.n4291 833.506
R152 dvss.n4292 dvss.n4248 833.506
R153 dvss.n4291 dvss.n4262 833.13
R154 dvss.n4262 dvss.n4248 833.13
R155 dvss.t735 dvss.t747 819.513
R156 dvss.t747 dvss.t737 819.513
R157 dvss.t737 dvss.t749 819.513
R158 dvss.t749 dvss.t729 819.513
R159 dvss.t729 dvss.t753 819.513
R160 dvss.t753 dvss.t755 819.513
R161 dvss.t755 dvss.t743 819.513
R162 dvss.t743 dvss.t733 819.513
R163 dvss.t733 dvss.t739 819.513
R164 dvss.t739 dvss.t757 819.513
R165 dvss.t741 dvss.t727 819.513
R166 dvss.t727 dvss.t751 819.513
R167 dvss.t751 dvss.t731 819.513
R168 dvss.t731 dvss.t745 819.513
R169 dvss.t632 dvss.t634 819.513
R170 dvss.t634 dvss.t630 819.513
R171 dvss.t630 dvss.t636 819.513
R172 dvss.t673 dvss.t653 808.754
R173 dvss.t653 dvss.t675 808.754
R174 dvss.t675 dvss.t655 808.754
R175 dvss.t655 dvss.t667 808.754
R176 dvss.t667 dvss.t659 808.754
R177 dvss.t659 dvss.t661 808.754
R178 dvss.t661 dvss.t649 808.754
R179 dvss.t649 dvss.t671 808.754
R180 dvss.t671 dvss.t677 808.754
R181 dvss.t677 dvss.t663 808.754
R182 dvss.t679 dvss.t665 808.754
R183 dvss.t665 dvss.t657 808.754
R184 dvss.t657 dvss.t669 808.754
R185 dvss.t669 dvss.t651 808.754
R186 dvss.t556 dvss.t550 808.754
R187 dvss.t550 dvss.t542 808.754
R188 dvss.t542 dvss.t546 808.754
R189 dvss.n2181 dvss.n2175 769.572
R190 dvss.n3142 dvss.n3141 769.572
R191 dvss.n4303 dvss.n58 769.572
R192 dvss.n4187 dvss.t465 761.905
R193 dvss.n4152 dvss.t43 761.905
R194 dvss.n3238 dvss.t10 761.905
R195 dvss.t245 dvss.n351 761.905
R196 dvss.n1946 dvss.t204 761.905
R197 dvss.n1681 dvss.t325 761.905
R198 dvss.n1389 dvss.t214 761.905
R199 dvss.n687 dvss.t226 761.905
R200 dvss.n1162 dvss.t28 761.905
R201 dvss.t745 dvss 760.976
R202 dvss.t651 dvss 750.986
R203 dvss.n4072 dvss.n179 747.437
R204 dvss.n3817 dvss.n3816 747.437
R205 dvss.n3665 dvss.n324 747.437
R206 dvss.n3562 dvss.n382 747.437
R207 dvss.n3442 dvss.n444 747.437
R208 dvss.n1656 dvss.n1644 747.437
R209 dvss.n1491 dvss.n563 747.437
R210 dvss.n1258 dvss.n1257 747.437
R211 dvss.t563 dvss.t565 745.433
R212 dvss.t636 dvss 731.707
R213 dvss.t546 dvss 722.101
R214 dvss.n2411 dvss.t59 682.76
R215 dvss.n836 dvss.t250 610.777
R216 dvss.n4156 dvss.n4155 607.51
R217 dvss.n4180 dvss.n50 607.51
R218 dvss.n4153 dvss.t186 604.145
R219 dvss.n2249 dvss.n2150 593.402
R220 dvss.n4154 dvss.n101 592.001
R221 dvss.n4181 dvss.n49 592.001
R222 dvss.n3982 dvss.n3981 590.068
R223 dvss.n3907 dvss.n3906 590.068
R224 dvss.n1993 dvss.n1992 590.068
R225 dvss.n1968 dvss.n1967 590.068
R226 dvss.n1941 dvss.n1940 590.068
R227 dvss.n1776 dvss.n1775 590.068
R228 dvss.n1384 dvss.n1383 590.068
R229 dvss.n1293 dvss.n1292 590.068
R230 dvss.n897 dvss.n890 590.068
R231 dvss.n4182 dvss.n4179 588.516
R232 dvss.n2250 dvss.n2161 587.614
R233 dvss.n3985 dvss.n3972 587.271
R234 dvss.n3920 dvss.n240 587.271
R235 dvss.n1996 dvss.n1919 587.271
R236 dvss.n1971 dvss.n1925 587.271
R237 dvss.n1944 dvss.n1931 587.271
R238 dvss.n1789 dvss.n486 587.271
R239 dvss.n1387 dvss.n1374 587.271
R240 dvss.n1306 dvss.n606 587.271
R241 dvss.n962 dvss.n961 587.271
R242 dvss.n2252 dvss.n2251 586.313
R243 dvss.n2183 dvss.n2182 585
R244 dvss.n2177 dvss.n2176 585
R245 dvss.n2178 dvss.n2177 585
R246 dvss.n2173 dvss.n2172 585
R247 dvss.n2172 dvss.n2171 585
R248 dvss.n2194 dvss.n2193 585
R249 dvss.n2195 dvss.n2194 585
R250 dvss.n2170 dvss.n2169 585
R251 dvss.n2196 dvss.n2170 585
R252 dvss.n2199 dvss.n2198 585
R253 dvss.n2198 dvss.n2197 585
R254 dvss.n2168 dvss.n2167 585
R255 dvss.n2167 dvss.n2166 585
R256 dvss.n2205 dvss.n2204 585
R257 dvss.n2206 dvss.n2205 585
R258 dvss.n2165 dvss.n2164 585
R259 dvss.n2207 dvss.n2165 585
R260 dvss.n2238 dvss.n2237 585
R261 dvss.n2237 dvss.n2236 585
R262 dvss.n2163 dvss.n2162 585
R263 dvss.n2235 dvss.n2162 585
R264 dvss.n2246 dvss.n2245 585
R265 dvss.n2247 dvss.n2246 585
R266 dvss.n2160 dvss.n2156 585
R267 dvss.n2248 dvss.n2160 585
R268 dvss.n2253 dvss.n2252 585
R269 dvss.n2161 dvss.n2159 585
R270 dvss.n2151 dvss.n2150 585
R271 dvss.n2264 dvss.n2263 585
R272 dvss.n2265 dvss.n2264 585
R273 dvss.n2149 dvss.n2148 585
R274 dvss.n2266 dvss.n2149 585
R275 dvss.n2269 dvss.n2268 585
R276 dvss.n2268 dvss.n2267 585
R277 dvss.n2147 dvss.n2146 585
R278 dvss.n2146 dvss.n2145 585
R279 dvss.n2517 dvss.n2516 585
R280 dvss.n2518 dvss.n2517 585
R281 dvss.n2091 dvss.n2090 585
R282 dvss.n2090 dvss.n2089 585
R283 dvss.n3195 dvss.n3194 585
R284 dvss.n3196 dvss.n3195 585
R285 dvss.n2088 dvss.n2087 585
R286 dvss.n3197 dvss.n2088 585
R287 dvss.n3201 dvss.n3200 585
R288 dvss.n3200 dvss.n3199 585
R289 dvss.n2085 dvss.n2084 585
R290 dvss.n3198 dvss.n2084 585
R291 dvss.n3211 dvss.n3210 585
R292 dvss.n3212 dvss.n3211 585
R293 dvss.n2083 dvss.n2082 585
R294 dvss.n3213 dvss.n2083 585
R295 dvss.n3216 dvss.n3215 585
R296 dvss.n3215 dvss.n3214 585
R297 dvss.n2081 dvss.n2080 585
R298 dvss.n2080 dvss.n2079 585
R299 dvss.n3222 dvss.n3221 585
R300 dvss.n3223 dvss.n3222 585
R301 dvss.n2078 dvss.n2077 585
R302 dvss.n3224 dvss.n2078 585
R303 dvss.n3228 dvss.n3227 585
R304 dvss.n3227 dvss.n3226 585
R305 dvss.n2000 dvss.n1998 585
R306 dvss.n3225 dvss.n1998 585
R307 dvss.n3236 dvss.n3235 585
R308 dvss.n3237 dvss.n3236 585
R309 dvss.n2001 dvss.n1999 585
R310 dvss.n2012 dvss.n1999 585
R311 dvss.n2015 dvss.n2014 585
R312 dvss.n2014 dvss.n2013 585
R313 dvss.n2009 dvss.n2008 585
R314 dvss.n2008 dvss.n2007 585
R315 dvss.n2024 dvss.n2023 585
R316 dvss.n2025 dvss.n2024 585
R317 dvss.n2010 dvss.n2006 585
R318 dvss.n2026 dvss.n2006 585
R319 dvss.n2028 dvss.n2005 585
R320 dvss.n2028 dvss.n2027 585
R321 dvss.n2071 dvss.n2029 585
R322 dvss.n2039 dvss.n2029 585
R323 dvss.n2070 dvss.n2030 585
R324 dvss.n2040 dvss.n2030 585
R325 dvss.n2041 dvss.n2031 585
R326 dvss.n2042 dvss.n2041 585
R327 dvss.n2066 dvss.n2032 585
R328 dvss.n2043 dvss.n2032 585
R329 dvss.n2065 dvss.n2033 585
R330 dvss.n2044 dvss.n2033 585
R331 dvss.n2037 dvss.n2034 585
R332 dvss.n2045 dvss.n2037 585
R333 dvss.n2058 dvss.n2057 585
R334 dvss.n2057 dvss.n2056 585
R335 dvss.n2038 dvss.n10 585
R336 dvss.n2055 dvss.n2038 585
R337 dvss.n4387 dvss.n11 585
R338 dvss.n2054 dvss.n11 585
R339 dvss.n4386 dvss.n12 585
R340 dvss.n2053 dvss.n12 585
R341 dvss.n2051 dvss.n13 585
R342 dvss.n2052 dvss.n2051 585
R343 dvss.n4382 dvss.n14 585
R344 dvss.n2050 dvss.n14 585
R345 dvss.n4381 dvss.n15 585
R346 dvss.n2049 dvss.n15 585
R347 dvss.n2047 dvss.n16 585
R348 dvss.n2048 dvss.n2047 585
R349 dvss.n4377 dvss.n17 585
R350 dvss.n2046 dvss.n17 585
R351 dvss.n4376 dvss.n18 585
R352 dvss.n106 dvss.n18 585
R353 dvss.n120 dvss.n19 585
R354 dvss.n121 dvss.n120 585
R355 dvss.n119 dvss.n118 585
R356 dvss.n119 dvss.n104 585
R357 dvss.n108 dvss.n107 585
R358 dvss.n107 dvss.n105 585
R359 dvss.n112 dvss.n101 585
R360 dvss.n4156 dvss.n102 585
R361 dvss.n4157 dvss.n23 585
R362 dvss.n4158 dvss.n4157 585
R363 dvss.n4366 dvss.n24 585
R364 dvss.n4159 dvss.n24 585
R365 dvss.n4365 dvss.n25 585
R366 dvss.n4160 dvss.n25 585
R367 dvss.n4161 dvss.n26 585
R368 dvss.n4162 dvss.n4161 585
R369 dvss.n4361 dvss.n27 585
R370 dvss.n4163 dvss.n27 585
R371 dvss.n4360 dvss.n28 585
R372 dvss.n4164 dvss.n28 585
R373 dvss.n4166 dvss.n29 585
R374 dvss.n4166 dvss.n4165 585
R375 dvss.n4167 dvss.n33 585
R376 dvss.n4168 dvss.n4167 585
R377 dvss.n4353 dvss.n34 585
R378 dvss.n4169 dvss.n34 585
R379 dvss.n4352 dvss.n35 585
R380 dvss.n4170 dvss.n35 585
R381 dvss.n4171 dvss.n36 585
R382 dvss.n4172 dvss.n4171 585
R383 dvss.n4348 dvss.n37 585
R384 dvss.n4173 dvss.n37 585
R385 dvss.n4347 dvss.n38 585
R386 dvss.n4174 dvss.n38 585
R387 dvss.n4175 dvss.n39 585
R388 dvss.n4176 dvss.n4175 585
R389 dvss.n4343 dvss.n40 585
R390 dvss.n4177 dvss.n40 585
R391 dvss.n4342 dvss.n41 585
R392 dvss.n4178 dvss.n41 585
R393 dvss.n4183 dvss.n42 585
R394 dvss.n4184 dvss.n4183 585
R395 dvss.n4335 dvss.n45 585
R396 dvss.n4186 dvss.n45 585
R397 dvss.n4334 dvss.n46 585
R398 dvss.n4185 dvss.n46 585
R399 dvss.n4179 dvss.n47 585
R400 dvss.n4327 dvss.n49 585
R401 dvss.n4326 dvss.n50 585
R402 dvss.n78 dvss.n51 585
R403 dvss.n79 dvss.n78 585
R404 dvss.n4319 dvss.n52 585
R405 dvss.n77 dvss.n52 585
R406 dvss.n4318 dvss.n53 585
R407 dvss.n76 dvss.n53 585
R408 dvss.n55 dvss.n54 585
R409 dvss.n56 dvss.n55 585
R410 dvss.n4314 dvss.n4313 585
R411 dvss.n4313 dvss.n4312 585
R412 dvss.n3152 dvss.n3151 585
R413 dvss.n3153 dvss.n3152 585
R414 dvss.n2110 dvss.n2109 585
R415 dvss.n3154 dvss.n2110 585
R416 dvss.n3157 dvss.n3156 585
R417 dvss.n3156 dvss.n3155 585
R418 dvss.n2108 dvss.n2107 585
R419 dvss.n2107 dvss.n2106 585
R420 dvss.n3165 dvss.n3164 585
R421 dvss.n3166 dvss.n3165 585
R422 dvss.n2104 dvss.n2100 585
R423 dvss.n3167 dvss.n2104 585
R424 dvss.n3172 dvss.n3171 585
R425 dvss.n3171 dvss.n3170 585
R426 dvss.n2105 dvss.n2103 585
R427 dvss.n3169 dvss.n2105 585
R428 dvss.n2095 dvss.n2094 585
R429 dvss.n3168 dvss.n2094 585
R430 dvss.n3183 dvss.n3182 585
R431 dvss.n3184 dvss.n3183 585
R432 dvss.n2093 dvss.n2092 585
R433 dvss.n3186 dvss.n2093 585
R434 dvss.n3189 dvss.n3188 585
R435 dvss.n3188 dvss.n3187 585
R436 dvss.n1487 dvss.n567 585
R437 dvss.n567 dvss.n563 585
R438 dvss.n1478 dvss.n570 585
R439 dvss.n1481 dvss.n1480 585
R440 dvss.n1477 dvss.n559 585
R441 dvss.n1477 dvss.n563 585
R442 dvss.n557 dvss.n556 585
R443 dvss.n1492 dvss.n556 585
R444 dvss.n1504 dvss.n1503 585
R445 dvss.n1505 dvss.n1504 585
R446 dvss.n553 dvss.n552 585
R447 dvss.n1506 dvss.n552 585
R448 dvss.n1517 dvss.n1516 585
R449 dvss.n1517 dvss.n550 585
R450 dvss.n1518 dvss.n545 585
R451 dvss.n1519 dvss.n1518 585
R452 dvss.n1531 dvss.n546 585
R453 dvss.n551 dvss.n546 585
R454 dvss.n1532 dvss.n541 585
R455 dvss.n1537 dvss.n541 585
R456 dvss.n1541 dvss.n542 585
R457 dvss.n1541 dvss.n1540 585
R458 dvss.n1542 dvss.n536 585
R459 dvss.n1543 dvss.n1542 585
R460 dvss.n1552 dvss.n537 585
R461 dvss.n1388 dvss.n537 585
R462 dvss.n1553 dvss.n531 585
R463 dvss.n533 dvss.n531 585
R464 dvss.n1566 dvss.n532 585
R465 dvss.n1566 dvss.n1565 585
R466 dvss.n1567 dvss.n524 585
R467 dvss.n1568 dvss.n1567 585
R468 dvss.n530 dvss.n529 585
R469 dvss.n1569 dvss.n530 585
R470 dvss.n1573 dvss.n1572 585
R471 dvss.n1572 dvss.n1571 585
R472 dvss.n510 dvss.n508 585
R473 dvss.n508 dvss.n505 585
R474 dvss.n1747 dvss.n1746 585
R475 dvss.n1748 dvss.n1747 585
R476 dvss.n511 dvss.n509 585
R477 dvss.n509 dvss.n507 585
R478 dvss.n1654 dvss.n1588 585
R479 dvss.n1653 dvss.n1589 585
R480 dvss.n1652 dvss.n1593 585
R481 dvss.n1658 dvss.n1594 585
R482 dvss.n1660 dvss.n1659 585
R483 dvss.n1661 dvss.n1660 585
R484 dvss.n1643 dvss.n1598 585
R485 dvss.n1662 dvss.n1643 585
R486 dvss.n1664 dvss.n1603 585
R487 dvss.n1664 dvss.n1663 585
R488 dvss.n1666 dvss.n1665 585
R489 dvss.n1665 dvss.n1640 585
R490 dvss.n1670 dvss.n1669 585
R491 dvss.n1671 dvss.n1670 585
R492 dvss.n1639 dvss.n1609 585
R493 dvss.n1672 dvss.n1639 585
R494 dvss.n1675 dvss.n1614 585
R495 dvss.n1675 dvss.n1674 585
R496 dvss.n1676 dvss.n1615 585
R497 dvss.n1677 dvss.n1676 585
R498 dvss.n1637 dvss.n1636 585
R499 dvss.n1680 dvss.n1637 585
R500 dvss.n1683 dvss.n1618 585
R501 dvss.n1683 dvss.n1682 585
R502 dvss.n1684 dvss.n1626 585
R503 dvss.n1685 dvss.n1684 585
R504 dvss.n1634 dvss.n1627 585
R505 dvss.n1686 dvss.n1634 585
R506 dvss.n1690 dvss.n1635 585
R507 dvss.n1690 dvss.n1689 585
R508 dvss.n1691 dvss.n1631 585
R509 dvss.n1692 dvss.n1691 585
R510 dvss.n460 dvss.n459 585
R511 dvss.n1693 dvss.n460 585
R512 dvss.n3412 dvss.n3411 585
R513 dvss.n3411 dvss.n3410 585
R514 dvss.n449 dvss.n447 585
R515 dvss.n447 dvss.n445 585
R516 dvss.n3440 dvss.n3439 585
R517 dvss.n3441 dvss.n3440 585
R518 dvss.n450 dvss.n448 585
R519 dvss.n3428 dvss.n3426 585
R520 dvss.n3432 dvss.n3431 585
R521 dvss.n3429 dvss.n440 585
R522 dvss.n438 dvss.n437 585
R523 dvss.n3443 dvss.n437 585
R524 dvss.n3455 dvss.n3454 585
R525 dvss.n3456 dvss.n3455 585
R526 dvss.n434 dvss.n433 585
R527 dvss.n3457 dvss.n433 585
R528 dvss.n3468 dvss.n3467 585
R529 dvss.n3468 dvss.n431 585
R530 dvss.n3469 dvss.n426 585
R531 dvss.n3470 dvss.n3469 585
R532 dvss.n3482 dvss.n427 585
R533 dvss.n432 dvss.n427 585
R534 dvss.n3483 dvss.n422 585
R535 dvss.n3488 dvss.n422 585
R536 dvss.n3492 dvss.n423 585
R537 dvss.n3492 dvss.n3491 585
R538 dvss.n3493 dvss.n417 585
R539 dvss.n3494 dvss.n3493 585
R540 dvss.n3503 dvss.n418 585
R541 dvss.n1945 dvss.n418 585
R542 dvss.n3504 dvss.n412 585
R543 dvss.n414 dvss.n412 585
R544 dvss.n3517 dvss.n413 585
R545 dvss.n3517 dvss.n3516 585
R546 dvss.n3518 dvss.n405 585
R547 dvss.n3519 dvss.n3518 585
R548 dvss.n411 dvss.n410 585
R549 dvss.n3520 dvss.n411 585
R550 dvss.n3525 dvss.n3524 585
R551 dvss.n3524 dvss.n3523 585
R552 dvss.n391 dvss.n390 585
R553 dvss.n3522 dvss.n390 585
R554 dvss.n3541 dvss.n3540 585
R555 dvss.n3542 dvss.n3541 585
R556 dvss.n385 dvss.n384 585
R557 dvss.n3543 dvss.n384 585
R558 dvss.n3560 dvss.n3559 585
R559 dvss.n386 dvss.n383 585
R560 dvss.n380 dvss.n379 585
R561 dvss.n3565 dvss.n3564 585
R562 dvss.n374 dvss.n373 585
R563 dvss.n381 dvss.n373 585
R564 dvss.n3577 dvss.n3576 585
R565 dvss.n3578 dvss.n3577 585
R566 dvss.n370 dvss.n369 585
R567 dvss.n3579 dvss.n370 585
R568 dvss.n3585 dvss.n3584 585
R569 dvss.n3584 dvss.n3583 585
R570 dvss.n364 dvss.n363 585
R571 dvss.n3582 dvss.n363 585
R572 dvss.n3603 dvss.n3602 585
R573 dvss.n3604 dvss.n3603 585
R574 dvss.n358 dvss.n357 585
R575 dvss.n360 dvss.n358 585
R576 dvss.n3609 dvss.n3608 585
R577 dvss.n3608 dvss.n3607 585
R578 dvss.n353 dvss.n352 585
R579 dvss.n359 dvss.n352 585
R580 dvss.n3620 dvss.n3619 585
R581 dvss.n3621 dvss.n3620 585
R582 dvss.n348 dvss.n347 585
R583 dvss.n347 dvss.n345 585
R584 dvss.n3634 dvss.n3633 585
R585 dvss.n3635 dvss.n3634 585
R586 dvss.n343 dvss.n337 585
R587 dvss.n3636 dvss.n343 585
R588 dvss.n3642 dvss.n3641 585
R589 dvss.n3641 dvss.n3640 585
R590 dvss.n344 dvss.n331 585
R591 dvss.n3639 dvss.n344 585
R592 dvss.n3654 dvss.n332 585
R593 dvss.n3638 dvss.n332 585
R594 dvss.n3655 dvss.n325 585
R595 dvss.n3660 dvss.n325 585
R596 dvss.n3662 dvss.n326 585
R597 dvss.n3662 dvss.n3661 585
R598 dvss.n3663 dvss.n319 585
R599 dvss.n321 dvss.n320 585
R600 dvss.n3668 dvss.n3667 585
R601 dvss.n322 dvss.n310 585
R602 dvss.n3686 dvss.n311 585
R603 dvss.n323 dvss.n311 585
R604 dvss.n3687 dvss.n306 585
R605 dvss.n3697 dvss.n306 585
R606 dvss.n3699 dvss.n307 585
R607 dvss.n3699 dvss.n3698 585
R608 dvss.n3700 dvss.n301 585
R609 dvss.n3701 dvss.n3700 585
R610 dvss.n296 dvss.n295 585
R611 dvss.n305 dvss.n295 585
R612 dvss.n3719 dvss.n3718 585
R613 dvss.n3720 dvss.n3719 585
R614 dvss.n297 dvss.n291 585
R615 dvss.n293 dvss.n291 585
R616 dvss.n3724 dvss.n292 585
R617 dvss.n3724 dvss.n3723 585
R618 dvss.n3725 dvss.n286 585
R619 dvss.n3726 dvss.n3725 585
R620 dvss.n3735 dvss.n287 585
R621 dvss.n1997 dvss.n287 585
R622 dvss.n3736 dvss.n281 585
R623 dvss.n283 dvss.n281 585
R624 dvss.n3749 dvss.n282 585
R625 dvss.n3749 dvss.n3748 585
R626 dvss.n3750 dvss.n274 585
R627 dvss.n3751 dvss.n3750 585
R628 dvss.n280 dvss.n279 585
R629 dvss.n3752 dvss.n280 585
R630 dvss.n3756 dvss.n3755 585
R631 dvss.n3755 dvss.n3754 585
R632 dvss.n265 dvss.n263 585
R633 dvss.n263 dvss.n260 585
R634 dvss.n3878 dvss.n3877 585
R635 dvss.n3879 dvss.n3878 585
R636 dvss.n266 dvss.n264 585
R637 dvss.n264 dvss.n262 585
R638 dvss.n3814 dvss.n3771 585
R639 dvss.n3813 dvss.n3772 585
R640 dvss.n3812 dvss.n3776 585
R641 dvss.n3810 dvss.n3777 585
R642 dvss.n3809 dvss.n3808 585
R643 dvss.n3825 dvss.n3809 585
R644 dvss.n3827 dvss.n3781 585
R645 dvss.n3827 dvss.n3826 585
R646 dvss.n3828 dvss.n3786 585
R647 dvss.n3829 dvss.n3828 585
R648 dvss.n3804 dvss.n3803 585
R649 dvss.n3830 dvss.n3803 585
R650 dvss.n3834 dvss.n3807 585
R651 dvss.n3834 dvss.n3833 585
R652 dvss.n3835 dvss.n3792 585
R653 dvss.n3836 dvss.n3835 585
R654 dvss.n3798 dvss.n3797 585
R655 dvss.n3802 dvss.n3798 585
R656 dvss.n3841 dvss.n3840 585
R657 dvss.n3840 dvss.n3839 585
R658 dvss.n125 dvss.n123 585
R659 dvss.n3799 dvss.n123 585
R660 dvss.n4150 dvss.n4149 585
R661 dvss.n4151 dvss.n4150 585
R662 dvss.n126 dvss.n124 585
R663 dvss.n196 dvss.n124 585
R664 dvss.n195 dvss.n130 585
R665 dvss.n197 dvss.n195 585
R666 dvss.n203 dvss.n202 585
R667 dvss.n202 dvss.n201 585
R668 dvss.n206 dvss.n205 585
R669 dvss.n207 dvss.n206 585
R670 dvss.n192 dvss.n191 585
R671 dvss.n208 dvss.n191 585
R672 dvss.n214 dvss.n213 585
R673 dvss.n215 dvss.n214 585
R674 dvss.n189 dvss.n139 585
R675 dvss.n4067 dvss.n189 585
R676 dvss.n4069 dvss.n144 585
R677 dvss.n4069 dvss.n4068 585
R678 dvss.n4070 dvss.n145 585
R679 dvss.n188 dvss.n146 585
R680 dvss.n187 dvss.n150 585
R681 dvss.n4074 dvss.n151 585
R682 dvss.n4076 dvss.n4075 585
R683 dvss.n4077 dvss.n4076 585
R684 dvss.n178 dvss.n155 585
R685 dvss.n4078 dvss.n178 585
R686 dvss.n4080 dvss.n160 585
R687 dvss.n4080 dvss.n4079 585
R688 dvss.n4082 dvss.n4081 585
R689 dvss.n4081 dvss.n175 585
R690 dvss.n4086 dvss.n4085 585
R691 dvss.n4087 dvss.n4086 585
R692 dvss.n174 dvss.n166 585
R693 dvss.n4088 dvss.n174 585
R694 dvss.n4091 dvss.n171 585
R695 dvss.n4091 dvss.n4090 585
R696 dvss.n4092 dvss.n172 585
R697 dvss.n4093 dvss.n4092 585
R698 dvss.n100 dvss.n99 585
R699 dvss.n4095 dvss.n100 585
R700 dvss.n4190 dvss.n4189 585
R701 dvss.n4189 dvss.n4188 585
R702 dvss.n94 dvss.n93 585
R703 dvss.n96 dvss.n94 585
R704 dvss.n4201 dvss.n4200 585
R705 dvss.n4200 dvss.n4199 585
R706 dvss.n95 dvss.n89 585
R707 dvss.n4198 dvss.n95 585
R708 dvss.n84 dvss.n83 585
R709 dvss.n4197 dvss.n83 585
R710 dvss.n4221 dvss.n4220 585
R711 dvss.n4222 dvss.n4221 585
R712 dvss.n75 dvss.n74 585
R713 dvss.n4225 dvss.n75 585
R714 dvss.n4229 dvss.n4228 585
R715 dvss.n4228 dvss.n4227 585
R716 dvss.n70 dvss.n68 585
R717 dvss.n68 dvss.n67 585
R718 dvss.n4236 dvss.n4235 585
R719 dvss.n4237 dvss.n4236 585
R720 dvss.n69 dvss.n64 585
R721 dvss.n69 dvss.n57 585
R722 dvss.n1261 dvss.n1260 585
R723 dvss.n635 dvss.n634 585
R724 dvss.n1209 dvss.n1208 585
R725 dvss.n641 dvss.n639 585
R726 dvss.n1255 dvss.n1254 585
R727 dvss.n1256 dvss.n1255 585
R728 dvss.n1253 dvss.n640 585
R729 dvss.n1219 dvss.n640 585
R730 dvss.n1252 dvss.n1251 585
R731 dvss.n1251 dvss.n1250 585
R732 dvss.n646 dvss.n645 585
R733 dvss.n1249 dvss.n646 585
R734 dvss.n1247 dvss.n1246 585
R735 dvss.n1248 dvss.n1247 585
R736 dvss.n1245 dvss.n650 585
R737 dvss.n657 dvss.n650 585
R738 dvss.n1244 dvss.n1243 585
R739 dvss.n1243 dvss.n1242 585
R740 dvss.n655 dvss.n654 585
R741 dvss.n683 dvss.n655 585
R742 dvss.n682 dvss.n681 585
R743 dvss.n686 dvss.n682 585
R744 dvss.n689 dvss.n664 585
R745 dvss.n689 dvss.n688 585
R746 dvss.n690 dvss.n671 585
R747 dvss.n691 dvss.n690 585
R748 dvss.n679 dvss.n672 585
R749 dvss.n692 dvss.n679 585
R750 dvss.n696 dvss.n680 585
R751 dvss.n696 dvss.n695 585
R752 dvss.n697 dvss.n676 585
R753 dvss.n698 dvss.n697 585
R754 dvss.n580 dvss.n579 585
R755 dvss.n699 dvss.n580 585
R756 dvss.n1463 dvss.n1462 585
R757 dvss.n1462 dvss.n1461 585
R758 dvss.n568 dvss.n566 585
R759 dvss.n566 dvss.n564 585
R760 dvss.n1489 dvss.n1488 585
R761 dvss.n1490 dvss.n1489 585
R762 dvss.n1289 dvss.n1288 585
R763 dvss.n1290 dvss.n1289 585
R764 dvss.n614 dvss.n613 585
R765 dvss.n1291 dvss.n614 585
R766 dvss.n1294 dvss.n1293 585
R767 dvss.n609 dvss.n608 585
R768 dvss.n608 dvss.n607 585
R769 dvss.n1304 dvss.n1303 585
R770 dvss.n1305 dvss.n1304 585
R771 dvss.n606 dvss.n605 585
R772 dvss.n1310 dvss.n1309 585
R773 dvss.n1309 dvss.n1308 585
R774 dvss.n599 dvss.n598 585
R775 dvss.n1307 dvss.n598 585
R776 dvss.n1319 dvss.n1318 585
R777 dvss.n1320 dvss.n1319 585
R778 dvss.n597 dvss.n596 585
R779 dvss.n1321 dvss.n597 585
R780 dvss.n1325 dvss.n1324 585
R781 dvss.n1324 dvss.n1323 585
R782 dvss.n591 dvss.n590 585
R783 dvss.n1322 dvss.n590 585
R784 dvss.n1334 dvss.n1333 585
R785 dvss.n1335 dvss.n1334 585
R786 dvss.n589 dvss.n588 585
R787 dvss.n1336 dvss.n589 585
R788 dvss.n1339 dvss.n1338 585
R789 dvss.n1338 dvss.n1337 585
R790 dvss.n586 dvss.n584 585
R791 dvss.n584 dvss.n582 585
R792 dvss.n1457 dvss.n1456 585
R793 dvss.n1458 dvss.n1457 585
R794 dvss.n587 dvss.n585 585
R795 dvss.n585 dvss.n583 585
R796 dvss.n1452 dvss.n1347 585
R797 dvss.n1451 dvss.n1348 585
R798 dvss.n1375 dvss.n1349 585
R799 dvss.n1447 dvss.n1350 585
R800 dvss.n1446 dvss.n1351 585
R801 dvss.n1380 dvss.n1351 585
R802 dvss.n1382 dvss.n1352 585
R803 dvss.n1382 dvss.n1381 585
R804 dvss.n1383 dvss.n1355 585
R805 dvss.n1438 dvss.n1356 585
R806 dvss.n1385 dvss.n1356 585
R807 dvss.n1437 dvss.n1357 585
R808 dvss.n1386 dvss.n1357 585
R809 dvss.n1374 dvss.n1358 585
R810 dvss.n1429 dvss.n1362 585
R811 dvss.n1390 dvss.n1362 585
R812 dvss.n1428 dvss.n1363 585
R813 dvss.n1391 dvss.n1363 585
R814 dvss.n1392 dvss.n1364 585
R815 dvss.n1393 dvss.n1392 585
R816 dvss.n1421 dvss.n1366 585
R817 dvss.n1394 dvss.n1366 585
R818 dvss.n1420 dvss.n1367 585
R819 dvss.n1395 dvss.n1367 585
R820 dvss.n1397 dvss.n1368 585
R821 dvss.n1397 dvss.n1396 585
R822 dvss.n1398 dvss.n1372 585
R823 dvss.n1399 dvss.n1398 585
R824 dvss.n1411 dvss.n1373 585
R825 dvss.n1400 dvss.n1373 585
R826 dvss.n1410 dvss.n1402 585
R827 dvss.n1402 dvss.n1401 585
R828 dvss.n503 dvss.n502 585
R829 dvss.n504 dvss.n503 585
R830 dvss.n1754 dvss.n1753 585
R831 dvss.n1753 dvss.n1752 585
R832 dvss.n501 dvss.n500 585
R833 dvss.n1751 dvss.n500 585
R834 dvss.n1760 dvss.n1759 585
R835 dvss.n499 dvss.n498 585
R836 dvss.n1765 dvss.n1764 585
R837 dvss.n497 dvss.n496 585
R838 dvss.n1772 dvss.n1771 585
R839 dvss.n1773 dvss.n1772 585
R840 dvss.n494 dvss.n493 585
R841 dvss.n1774 dvss.n494 585
R842 dvss.n1777 dvss.n1776 585
R843 dvss.n489 dvss.n488 585
R844 dvss.n488 dvss.n487 585
R845 dvss.n1787 dvss.n1786 585
R846 dvss.n1788 dvss.n1787 585
R847 dvss.n486 dvss.n485 585
R848 dvss.n1793 dvss.n1792 585
R849 dvss.n1792 dvss.n1791 585
R850 dvss.n479 dvss.n478 585
R851 dvss.n1790 dvss.n478 585
R852 dvss.n1802 dvss.n1801 585
R853 dvss.n1803 dvss.n1802 585
R854 dvss.n477 dvss.n476 585
R855 dvss.n1804 dvss.n477 585
R856 dvss.n1808 dvss.n1807 585
R857 dvss.n1807 dvss.n1806 585
R858 dvss.n471 dvss.n470 585
R859 dvss.n1805 dvss.n470 585
R860 dvss.n1817 dvss.n1816 585
R861 dvss.n1818 dvss.n1817 585
R862 dvss.n469 dvss.n468 585
R863 dvss.n1819 dvss.n469 585
R864 dvss.n1822 dvss.n1821 585
R865 dvss.n1821 dvss.n1820 585
R866 dvss.n466 dvss.n464 585
R867 dvss.n464 dvss.n462 585
R868 dvss.n3406 dvss.n3405 585
R869 dvss.n3407 dvss.n3406 585
R870 dvss.n467 dvss.n465 585
R871 dvss.n465 dvss.n463 585
R872 dvss.n3401 dvss.n1830 585
R873 dvss.n3400 dvss.n1831 585
R874 dvss.n1932 dvss.n1832 585
R875 dvss.n3396 dvss.n1833 585
R876 dvss.n3395 dvss.n1834 585
R877 dvss.n1937 dvss.n1834 585
R878 dvss.n1939 dvss.n1835 585
R879 dvss.n1939 dvss.n1938 585
R880 dvss.n1940 dvss.n1838 585
R881 dvss.n3387 dvss.n1839 585
R882 dvss.n1942 dvss.n1839 585
R883 dvss.n3386 dvss.n1840 585
R884 dvss.n1943 dvss.n1840 585
R885 dvss.n1931 dvss.n1841 585
R886 dvss.n3378 dvss.n1845 585
R887 dvss.n1947 dvss.n1845 585
R888 dvss.n3377 dvss.n1846 585
R889 dvss.n1948 dvss.n1846 585
R890 dvss.n1949 dvss.n1847 585
R891 dvss.n1950 dvss.n1949 585
R892 dvss.n3370 dvss.n1849 585
R893 dvss.n1951 dvss.n1849 585
R894 dvss.n3369 dvss.n1850 585
R895 dvss.n1952 dvss.n1850 585
R896 dvss.n1954 dvss.n1851 585
R897 dvss.n1954 dvss.n1953 585
R898 dvss.n1955 dvss.n1855 585
R899 dvss.n1956 dvss.n1955 585
R900 dvss.n3360 dvss.n1856 585
R901 dvss.n1957 dvss.n1856 585
R902 dvss.n3359 dvss.n1857 585
R903 dvss.n1958 dvss.n1857 585
R904 dvss.n1959 dvss.n1858 585
R905 dvss.n1960 dvss.n1959 585
R906 dvss.n3350 dvss.n1859 585
R907 dvss.n1962 dvss.n1859 585
R908 dvss.n3349 dvss.n1860 585
R909 dvss.n1963 dvss.n1860 585
R910 dvss.n1928 dvss.n1861 585
R911 dvss.n3345 dvss.n1862 585
R912 dvss.n3344 dvss.n1863 585
R913 dvss.n1926 dvss.n1864 585
R914 dvss.n3340 dvss.n1865 585
R915 dvss.n1965 dvss.n1865 585
R916 dvss.n3339 dvss.n1866 585
R917 dvss.n1966 dvss.n1866 585
R918 dvss.n1967 dvss.n1867 585
R919 dvss.n3332 dvss.n1870 585
R920 dvss.n1969 dvss.n1870 585
R921 dvss.n3331 dvss.n1871 585
R922 dvss.n1970 dvss.n1871 585
R923 dvss.n1925 dvss.n1872 585
R924 dvss.n3323 dvss.n1876 585
R925 dvss.n1972 dvss.n1876 585
R926 dvss.n3322 dvss.n1877 585
R927 dvss.n1973 dvss.n1877 585
R928 dvss.n1974 dvss.n1878 585
R929 dvss.n1975 dvss.n1974 585
R930 dvss.n3315 dvss.n1880 585
R931 dvss.n1976 dvss.n1880 585
R932 dvss.n3314 dvss.n1881 585
R933 dvss.n1977 dvss.n1881 585
R934 dvss.n1979 dvss.n1882 585
R935 dvss.n1979 dvss.n1978 585
R936 dvss.n1980 dvss.n1886 585
R937 dvss.n1981 dvss.n1980 585
R938 dvss.n3305 dvss.n1887 585
R939 dvss.n1982 dvss.n1887 585
R940 dvss.n3304 dvss.n1888 585
R941 dvss.n1983 dvss.n1888 585
R942 dvss.n1984 dvss.n1889 585
R943 dvss.n1985 dvss.n1984 585
R944 dvss.n3300 dvss.n1890 585
R945 dvss.n1987 dvss.n1890 585
R946 dvss.n3299 dvss.n1891 585
R947 dvss.n1988 dvss.n1891 585
R948 dvss.n1922 dvss.n1892 585
R949 dvss.n3295 dvss.n1893 585
R950 dvss.n3294 dvss.n1894 585
R951 dvss.n1920 dvss.n1895 585
R952 dvss.n3290 dvss.n1896 585
R953 dvss.n1990 dvss.n1896 585
R954 dvss.n3289 dvss.n1897 585
R955 dvss.n1991 dvss.n1897 585
R956 dvss.n1992 dvss.n1898 585
R957 dvss.n3282 dvss.n1901 585
R958 dvss.n1994 dvss.n1901 585
R959 dvss.n3281 dvss.n1902 585
R960 dvss.n1995 dvss.n1902 585
R961 dvss.n1919 dvss.n1903 585
R962 dvss.n3273 dvss.n1907 585
R963 dvss.n3239 dvss.n1907 585
R964 dvss.n3272 dvss.n1908 585
R965 dvss.n3240 dvss.n1908 585
R966 dvss.n3241 dvss.n1909 585
R967 dvss.n3242 dvss.n3241 585
R968 dvss.n3265 dvss.n1911 585
R969 dvss.n3243 dvss.n1911 585
R970 dvss.n3264 dvss.n1912 585
R971 dvss.n3244 dvss.n1912 585
R972 dvss.n3246 dvss.n1913 585
R973 dvss.n3246 dvss.n3245 585
R974 dvss.n3247 dvss.n1917 585
R975 dvss.n3248 dvss.n3247 585
R976 dvss.n3255 dvss.n1918 585
R977 dvss.n3249 dvss.n1918 585
R978 dvss.n3254 dvss.n3251 585
R979 dvss.n3251 dvss.n3250 585
R980 dvss.n257 dvss.n256 585
R981 dvss.n258 dvss.n257 585
R982 dvss.n3885 dvss.n3884 585
R983 dvss.n3884 dvss.n3883 585
R984 dvss.n255 dvss.n254 585
R985 dvss.n3882 dvss.n254 585
R986 dvss.n3891 dvss.n3890 585
R987 dvss.n253 dvss.n252 585
R988 dvss.n3896 dvss.n3895 585
R989 dvss.n251 dvss.n250 585
R990 dvss.n3903 dvss.n3902 585
R991 dvss.n3904 dvss.n3903 585
R992 dvss.n248 dvss.n247 585
R993 dvss.n3905 dvss.n248 585
R994 dvss.n3908 dvss.n3907 585
R995 dvss.n243 dvss.n242 585
R996 dvss.n242 dvss.n241 585
R997 dvss.n3918 dvss.n3917 585
R998 dvss.n3919 dvss.n3918 585
R999 dvss.n240 dvss.n239 585
R1000 dvss.n3924 dvss.n3923 585
R1001 dvss.n3923 dvss.n3922 585
R1002 dvss.n233 dvss.n232 585
R1003 dvss.n3921 dvss.n232 585
R1004 dvss.n3933 dvss.n3932 585
R1005 dvss.n3934 dvss.n3933 585
R1006 dvss.n231 dvss.n230 585
R1007 dvss.n3935 dvss.n231 585
R1008 dvss.n3939 dvss.n3938 585
R1009 dvss.n3938 dvss.n3937 585
R1010 dvss.n225 dvss.n224 585
R1011 dvss.n3936 dvss.n224 585
R1012 dvss.n3948 dvss.n3947 585
R1013 dvss.n3949 dvss.n3948 585
R1014 dvss.n223 dvss.n222 585
R1015 dvss.n3950 dvss.n223 585
R1016 dvss.n3953 dvss.n3952 585
R1017 dvss.n3952 dvss.n3951 585
R1018 dvss.n220 dvss.n218 585
R1019 dvss.n218 dvss.n216 585
R1020 dvss.n4063 dvss.n4062 585
R1021 dvss.n4064 dvss.n4063 585
R1022 dvss.n221 dvss.n219 585
R1023 dvss.n219 dvss.n217 585
R1024 dvss.n4058 dvss.n3956 585
R1025 dvss.n4057 dvss.n3957 585
R1026 dvss.n3973 dvss.n3958 585
R1027 dvss.n4053 dvss.n3959 585
R1028 dvss.n4052 dvss.n3960 585
R1029 dvss.n3978 dvss.n3960 585
R1030 dvss.n3980 dvss.n3961 585
R1031 dvss.n3980 dvss.n3979 585
R1032 dvss.n3981 dvss.n3964 585
R1033 dvss.n4044 dvss.n3965 585
R1034 dvss.n3983 dvss.n3965 585
R1035 dvss.n4043 dvss.n3966 585
R1036 dvss.n3984 dvss.n3966 585
R1037 dvss.n3972 dvss.n3967 585
R1038 dvss.n4035 dvss.n3971 585
R1039 dvss.n3986 dvss.n3971 585
R1040 dvss.n4034 dvss.n3988 585
R1041 dvss.n3988 dvss.n3987 585
R1042 dvss.n4000 dvss.n3989 585
R1043 dvss.n4001 dvss.n4000 585
R1044 dvss.n4027 dvss.n3991 585
R1045 dvss.n4002 dvss.n3991 585
R1046 dvss.n4026 dvss.n3992 585
R1047 dvss.n4003 dvss.n3992 585
R1048 dvss.n4005 dvss.n3993 585
R1049 dvss.n4005 dvss.n4004 585
R1050 dvss.n4006 dvss.n3997 585
R1051 dvss.n4007 dvss.n4006 585
R1052 dvss.n4017 dvss.n3998 585
R1053 dvss.n4008 dvss.n3998 585
R1054 dvss.n4016 dvss.n3999 585
R1055 dvss.n4009 dvss.n3999 585
R1056 dvss.n4012 dvss.n4011 585
R1057 dvss.n4011 dvss.n4010 585
R1058 dvss.n62 dvss.n60 585
R1059 dvss.n60 dvss.n59 585
R1060 dvss.n4308 dvss.n4307 585
R1061 dvss.n4309 dvss.n4308 585
R1062 dvss.n63 dvss.n61 585
R1063 dvss.n1277 dvss.n1276 585
R1064 dvss.n619 dvss.n618 585
R1065 dvss.n1282 dvss.n1281 585
R1066 dvss.n617 dvss.n616 585
R1067 dvss.n889 dvss.n888 585
R1068 dvss.n971 dvss.n889 585
R1069 dvss.n969 dvss.n968 585
R1070 dvss.n970 dvss.n969 585
R1071 dvss.n967 dvss.n890 585
R1072 dvss.n966 dvss.n965 585
R1073 dvss.n965 dvss.n964 585
R1074 dvss.n896 dvss.n895 585
R1075 dvss.n963 dvss.n896 585
R1076 dvss.n961 dvss.n960 585
R1077 dvss.n959 dvss.n898 585
R1078 dvss.n955 dvss.n898 585
R1079 dvss.n958 dvss.n957 585
R1080 dvss.n957 dvss.n956 585
R1081 dvss.n954 dvss.n902 585
R1082 dvss.n954 dvss.n953 585
R1083 dvss.n906 dvss.n903 585
R1084 dvss.n952 dvss.n903 585
R1085 dvss.n950 dvss.n949 585
R1086 dvss.n951 dvss.n950 585
R1087 dvss.n948 dvss.n905 585
R1088 dvss.n905 dvss.n904 585
R1089 dvss.n947 dvss.n946 585
R1090 dvss.n946 dvss.n945 585
R1091 dvss.n930 dvss.n929 585
R1092 dvss.n944 dvss.n930 585
R1093 dvss.n942 dvss.n941 585
R1094 dvss.n943 dvss.n942 585
R1095 dvss.n623 dvss.n622 585
R1096 dvss.n624 dvss.n623 585
R1097 dvss.n1271 dvss.n1270 585
R1098 dvss.n1270 dvss.n1269 585
R1099 dvss.n621 dvss.n620 585
R1100 dvss.n1268 dvss.n620 585
R1101 dvss.n1146 dvss.n1143 585
R1102 dvss.n1146 dvss.n1145 585
R1103 dvss.n750 dvss.n747 585
R1104 dvss.n1161 dvss.n750 585
R1105 dvss.n1165 dvss.n1164 585
R1106 dvss.n1164 dvss.n1163 585
R1107 dvss.n1166 dvss.n742 585
R1108 dvss.n744 dvss.n742 585
R1109 dvss.n1179 dvss.n743 585
R1110 dvss.n1179 dvss.n1178 585
R1111 dvss.n1180 dvss.n735 585
R1112 dvss.n1181 dvss.n1180 585
R1113 dvss.n741 dvss.n740 585
R1114 dvss.n1182 dvss.n741 585
R1115 dvss.n1186 dvss.n1185 585
R1116 dvss.n1185 dvss.n1184 585
R1117 dvss.n630 dvss.n628 585
R1118 dvss.n628 dvss.n625 585
R1119 dvss.n1264 dvss.n1263 585
R1120 dvss.n1265 dvss.n1264 585
R1121 dvss.n1262 dvss.n629 585
R1122 dvss.n629 dvss.n627 585
R1123 dvss.n1119 dvss.n1118 585
R1124 dvss.n1118 dvss.n1117 585
R1125 dvss.n1120 dvss.n770 585
R1126 dvss.n777 dvss.n770 585
R1127 dvss.n1127 dvss.n769 585
R1128 dvss.n1127 dvss.n1126 585
R1129 dvss.n1129 dvss.n1128 585
R1130 dvss.n1128 dvss.n762 585
R1131 dvss.n765 dvss.n760 585
R1132 dvss.n1139 dvss.n760 585
R1133 dvss.n1141 dvss.n761 585
R1134 dvss.n1141 dvss.n1140 585
R1135 dvss.n1147 dvss.n756 585
R1136 dvss.n1148 dvss.n1147 585
R1137 dvss.n1116 dvss.n1115 585
R1138 dvss.n1117 dvss.n1116 585
R1139 dvss.n772 dvss.n771 585
R1140 dvss.n777 dvss.n771 585
R1141 dvss.n1125 dvss.n1124 585
R1142 dvss.n1126 dvss.n1125 585
R1143 dvss.n764 dvss.n763 585
R1144 dvss.n763 dvss.n762 585
R1145 dvss.n1138 dvss.n1137 585
R1146 dvss.n1139 dvss.n1138 585
R1147 dvss.n758 dvss.n757 585
R1148 dvss.n1140 dvss.n758 585
R1149 dvss.n1150 dvss.n1149 585
R1150 dvss.n1149 dvss.n1148 585
R1151 dvss.n752 dvss.n751 585
R1152 dvss.n1145 dvss.n751 585
R1153 dvss.n1160 dvss.n1159 585
R1154 dvss.n1161 dvss.n1160 585
R1155 dvss.n746 dvss.n745 585
R1156 dvss.n1163 dvss.n745 585
R1157 dvss.n1176 dvss.n1175 585
R1158 dvss.n1176 dvss.n744 585
R1159 dvss.n1177 dvss.n737 585
R1160 dvss.n1178 dvss.n1177 585
R1161 dvss.n1190 dvss.n738 585
R1162 dvss.n1181 dvss.n738 585
R1163 dvss.n1189 dvss.n739 585
R1164 dvss.n1182 dvss.n739 585
R1165 dvss.n1183 dvss.n729 585
R1166 dvss.n1184 dvss.n1183 585
R1167 dvss.n1199 dvss.n730 585
R1168 dvss.n730 dvss.n625 585
R1169 dvss.n1200 dvss.n626 585
R1170 dvss.n1265 dvss.n626 585
R1171 dvss.n1202 dvss.n1201 585
R1172 dvss.n1202 dvss.n627 585
R1173 dvss.n1203 dvss.n725 585
R1174 dvss.n1206 dvss.n1205 585
R1175 dvss.n726 dvss.n723 585
R1176 dvss.n1217 dvss.n724 585
R1177 dvss.n1218 dvss.n638 585
R1178 dvss.n1256 dvss.n638 585
R1179 dvss.n1221 dvss.n1220 585
R1180 dvss.n1220 dvss.n1219 585
R1181 dvss.n1222 dvss.n647 585
R1182 dvss.n1250 dvss.n647 585
R1183 dvss.n1224 dvss.n648 585
R1184 dvss.n1249 dvss.n648 585
R1185 dvss.n1223 dvss.n649 585
R1186 dvss.n1248 dvss.n649 585
R1187 dvss.n660 dvss.n658 585
R1188 dvss.n658 dvss.n657 585
R1189 dvss.n1241 dvss.n1240 585
R1190 dvss.n1242 dvss.n1241 585
R1191 dvss.n1239 dvss.n659 585
R1192 dvss.n683 dvss.n659 585
R1193 dvss.n685 dvss.n661 585
R1194 dvss.n686 dvss.n685 585
R1195 dvss.n717 dvss.n665 585
R1196 dvss.n688 dvss.n665 585
R1197 dvss.n716 dvss.n666 585
R1198 dvss.n691 dvss.n666 585
R1199 dvss.n693 dvss.n667 585
R1200 dvss.n693 dvss.n692 585
R1201 dvss.n694 dvss.n677 585
R1202 dvss.n695 dvss.n694 585
R1203 dvss.n703 dvss.n678 585
R1204 dvss.n698 dvss.n678 585
R1205 dvss.n702 dvss.n700 585
R1206 dvss.n700 dvss.n699 585
R1207 dvss.n581 dvss.n571 585
R1208 dvss.n1461 dvss.n581 585
R1209 dvss.n1469 dvss.n572 585
R1210 dvss.n572 dvss.n564 585
R1211 dvss.n1470 dvss.n565 585
R1212 dvss.n1490 dvss.n565 585
R1213 dvss.n1485 dvss.n1471 585
R1214 dvss.n1484 dvss.n1476 585
R1215 dvss.n1472 dvss.n560 585
R1216 dvss.n1495 dvss.n561 585
R1217 dvss.n1494 dvss.n1493 585
R1218 dvss.n1493 dvss.n1492 585
R1219 dvss.n555 dvss.n554 585
R1220 dvss.n1505 dvss.n555 585
R1221 dvss.n1508 dvss.n1507 585
R1222 dvss.n1507 dvss.n1506 585
R1223 dvss.n549 dvss.n548 585
R1224 dvss.n550 dvss.n549 585
R1225 dvss.n1521 dvss.n1520 585
R1226 dvss.n1520 dvss.n1519 585
R1227 dvss.n544 dvss.n543 585
R1228 dvss.n551 dvss.n543 585
R1229 dvss.n1536 dvss.n1535 585
R1230 dvss.n1537 dvss.n1536 585
R1231 dvss.n540 dvss.n539 585
R1232 dvss.n1540 dvss.n540 585
R1233 dvss.n1545 dvss.n1544 585
R1234 dvss.n1544 dvss.n1543 585
R1235 dvss.n535 dvss.n534 585
R1236 dvss.n1388 dvss.n534 585
R1237 dvss.n1563 dvss.n1562 585
R1238 dvss.n1563 dvss.n533 585
R1239 dvss.n1564 dvss.n526 585
R1240 dvss.n1565 dvss.n1564 585
R1241 dvss.n1577 dvss.n527 585
R1242 dvss.n1568 dvss.n527 585
R1243 dvss.n1576 dvss.n528 585
R1244 dvss.n1569 dvss.n528 585
R1245 dvss.n1570 dvss.n513 585
R1246 dvss.n1571 dvss.n1570 585
R1247 dvss.n1585 dvss.n514 585
R1248 dvss.n514 dvss.n505 585
R1249 dvss.n1744 dvss.n506 585
R1250 dvss.n1748 dvss.n506 585
R1251 dvss.n1743 dvss.n1586 585
R1252 dvss.n1586 dvss.n507 585
R1253 dvss.n1646 dvss.n1587 585
R1254 dvss.n1739 dvss.n1590 585
R1255 dvss.n1738 dvss.n1591 585
R1256 dvss.n1650 dvss.n1592 585
R1257 dvss.n1651 dvss.n1599 585
R1258 dvss.n1661 dvss.n1651 585
R1259 dvss.n1731 dvss.n1600 585
R1260 dvss.n1662 dvss.n1600 585
R1261 dvss.n1730 dvss.n1601 585
R1262 dvss.n1663 dvss.n1601 585
R1263 dvss.n1641 dvss.n1602 585
R1264 dvss.n1641 dvss.n1640 585
R1265 dvss.n1642 dvss.n1610 585
R1266 dvss.n1671 dvss.n1642 585
R1267 dvss.n1722 dvss.n1611 585
R1268 dvss.n1672 dvss.n1611 585
R1269 dvss.n1721 dvss.n1612 585
R1270 dvss.n1674 dvss.n1612 585
R1271 dvss.n1678 dvss.n1613 585
R1272 dvss.n1678 dvss.n1677 585
R1273 dvss.n1679 dvss.n1619 585
R1274 dvss.n1680 dvss.n1679 585
R1275 dvss.n1711 dvss.n1620 585
R1276 dvss.n1682 dvss.n1620 585
R1277 dvss.n1710 dvss.n1621 585
R1278 dvss.n1685 dvss.n1621 585
R1279 dvss.n1687 dvss.n1622 585
R1280 dvss.n1687 dvss.n1686 585
R1281 dvss.n1688 dvss.n1632 585
R1282 dvss.n1689 dvss.n1688 585
R1283 dvss.n1697 dvss.n1633 585
R1284 dvss.n1692 dvss.n1633 585
R1285 dvss.n1696 dvss.n1694 585
R1286 dvss.n1694 dvss.n1693 585
R1287 dvss.n461 dvss.n451 585
R1288 dvss.n3410 dvss.n461 585
R1289 dvss.n3418 dvss.n452 585
R1290 dvss.n452 dvss.n445 585
R1291 dvss.n3437 dvss.n446 585
R1292 dvss.n3441 dvss.n446 585
R1293 dvss.n3436 dvss.n3419 585
R1294 dvss.n3425 dvss.n3424 585
R1295 dvss.n3420 dvss.n441 585
R1296 dvss.n3446 dvss.n442 585
R1297 dvss.n3445 dvss.n3444 585
R1298 dvss.n3444 dvss.n3443 585
R1299 dvss.n436 dvss.n435 585
R1300 dvss.n3456 dvss.n436 585
R1301 dvss.n3459 dvss.n3458 585
R1302 dvss.n3458 dvss.n3457 585
R1303 dvss.n430 dvss.n429 585
R1304 dvss.n431 dvss.n430 585
R1305 dvss.n3472 dvss.n3471 585
R1306 dvss.n3471 dvss.n3470 585
R1307 dvss.n425 dvss.n424 585
R1308 dvss.n432 dvss.n424 585
R1309 dvss.n3487 dvss.n3486 585
R1310 dvss.n3488 dvss.n3487 585
R1311 dvss.n421 dvss.n420 585
R1312 dvss.n3491 dvss.n421 585
R1313 dvss.n3496 dvss.n3495 585
R1314 dvss.n3495 dvss.n3494 585
R1315 dvss.n416 dvss.n415 585
R1316 dvss.n1945 dvss.n415 585
R1317 dvss.n3514 dvss.n3513 585
R1318 dvss.n3514 dvss.n414 585
R1319 dvss.n3515 dvss.n407 585
R1320 dvss.n3516 dvss.n3515 585
R1321 dvss.n3529 dvss.n408 585
R1322 dvss.n3519 dvss.n408 585
R1323 dvss.n3528 dvss.n409 585
R1324 dvss.n3520 dvss.n409 585
R1325 dvss.n3521 dvss.n394 585
R1326 dvss.n3523 dvss.n3521 585
R1327 dvss.n3537 dvss.n395 585
R1328 dvss.n3522 dvss.n395 585
R1329 dvss.n3538 dvss.n388 585
R1330 dvss.n3542 dvss.n388 585
R1331 dvss.n3544 dvss.n387 585
R1332 dvss.n3544 dvss.n3543 585
R1333 dvss.n3557 dvss.n3545 585
R1334 dvss.n3556 dvss.n3546 585
R1335 dvss.n3553 dvss.n3552 585
R1336 dvss.n3547 dvss.n377 585
R1337 dvss.n3573 dvss.n378 585
R1338 dvss.n381 dvss.n378 585
R1339 dvss.n3574 dvss.n371 585
R1340 dvss.n3578 dvss.n371 585
R1341 dvss.n3580 dvss.n372 585
R1342 dvss.n3580 dvss.n3579 585
R1343 dvss.n3581 dvss.n365 585
R1344 dvss.n3583 dvss.n3581 585
R1345 dvss.n3599 dvss.n366 585
R1346 dvss.n3582 dvss.n366 585
R1347 dvss.n3600 dvss.n362 585
R1348 dvss.n3604 dvss.n362 585
R1349 dvss.n361 dvss.n355 585
R1350 dvss.n361 dvss.n360 585
R1351 dvss.n3611 dvss.n356 585
R1352 dvss.n3607 dvss.n356 585
R1353 dvss.n3612 dvss.n350 585
R1354 dvss.n359 dvss.n350 585
R1355 dvss.n3622 dvss.n349 585
R1356 dvss.n3622 dvss.n3621 585
R1357 dvss.n3624 dvss.n3623 585
R1358 dvss.n3623 dvss.n345 585
R1359 dvss.n346 dvss.n339 585
R1360 dvss.n3635 dvss.n346 585
R1361 dvss.n3646 dvss.n340 585
R1362 dvss.n3636 dvss.n340 585
R1363 dvss.n3645 dvss.n341 585
R1364 dvss.n3640 dvss.n341 585
R1365 dvss.n3637 dvss.n342 585
R1366 dvss.n3639 dvss.n3637 585
R1367 dvss.n329 dvss.n328 585
R1368 dvss.n3638 dvss.n328 585
R1369 dvss.n3659 dvss.n3658 585
R1370 dvss.n3660 dvss.n3659 585
R1371 dvss.n317 dvss.n316 585
R1372 dvss.n3661 dvss.n316 585
R1373 dvss.n3673 dvss.n3672 585
R1374 dvss.n318 dvss.n315 585
R1375 dvss.n313 dvss.n312 585
R1376 dvss.n3678 dvss.n3677 585
R1377 dvss.n309 dvss.n308 585
R1378 dvss.n323 dvss.n308 585
R1379 dvss.n3696 dvss.n3695 585
R1380 dvss.n3697 dvss.n3696 585
R1381 dvss.n303 dvss.n302 585
R1382 dvss.n3698 dvss.n303 585
R1383 dvss.n3703 dvss.n3702 585
R1384 dvss.n3702 dvss.n3701 585
R1385 dvss.n304 dvss.n298 585
R1386 dvss.n305 dvss.n304 585
R1387 dvss.n3716 dvss.n294 585
R1388 dvss.n3720 dvss.n294 585
R1389 dvss.n3715 dvss.n299 585
R1390 dvss.n299 dvss.n293 585
R1391 dvss.n290 dvss.n289 585
R1392 dvss.n3723 dvss.n290 585
R1393 dvss.n3728 dvss.n3727 585
R1394 dvss.n3727 dvss.n3726 585
R1395 dvss.n285 dvss.n284 585
R1396 dvss.n1997 dvss.n284 585
R1397 dvss.n3746 dvss.n3745 585
R1398 dvss.n3746 dvss.n283 585
R1399 dvss.n3747 dvss.n276 585
R1400 dvss.n3748 dvss.n3747 585
R1401 dvss.n3760 dvss.n277 585
R1402 dvss.n3751 dvss.n277 585
R1403 dvss.n3759 dvss.n278 585
R1404 dvss.n3752 dvss.n278 585
R1405 dvss.n3753 dvss.n268 585
R1406 dvss.n3754 dvss.n3753 585
R1407 dvss.n3768 dvss.n269 585
R1408 dvss.n269 dvss.n260 585
R1409 dvss.n3875 dvss.n261 585
R1410 dvss.n3879 dvss.n261 585
R1411 dvss.n3874 dvss.n3769 585
R1412 dvss.n3769 dvss.n262 585
R1413 dvss.n3819 dvss.n3770 585
R1414 dvss.n3870 dvss.n3773 585
R1415 dvss.n3869 dvss.n3774 585
R1416 dvss.n3823 dvss.n3775 585
R1417 dvss.n3824 dvss.n3782 585
R1418 dvss.n3825 dvss.n3824 585
R1419 dvss.n3862 dvss.n3783 585
R1420 dvss.n3826 dvss.n3783 585
R1421 dvss.n3861 dvss.n3784 585
R1422 dvss.n3829 dvss.n3784 585
R1423 dvss.n3831 dvss.n3785 585
R1424 dvss.n3831 dvss.n3830 585
R1425 dvss.n3832 dvss.n3793 585
R1426 dvss.n3833 dvss.n3832 585
R1427 dvss.n3853 dvss.n3794 585
R1428 dvss.n3836 dvss.n3794 585
R1429 dvss.n3852 dvss.n3795 585
R1430 dvss.n3802 dvss.n3795 585
R1431 dvss.n3801 dvss.n3796 585
R1432 dvss.n3839 dvss.n3801 585
R1433 dvss.n3800 dvss.n127 585
R1434 dvss.n3800 dvss.n3799 585
R1435 dvss.n4147 dvss.n122 585
R1436 dvss.n4151 dvss.n122 585
R1437 dvss.n4146 dvss.n128 585
R1438 dvss.n196 dvss.n128 585
R1439 dvss.n198 dvss.n129 585
R1440 dvss.n198 dvss.n197 585
R1441 dvss.n200 dvss.n199 585
R1442 dvss.n201 dvss.n200 585
R1443 dvss.n194 dvss.n193 585
R1444 dvss.n207 dvss.n194 585
R1445 dvss.n210 dvss.n209 585
R1446 dvss.n209 dvss.n208 585
R1447 dvss.n190 dvss.n140 585
R1448 dvss.n215 dvss.n190 585
R1449 dvss.n4131 dvss.n141 585
R1450 dvss.n4067 dvss.n141 585
R1451 dvss.n4130 dvss.n142 585
R1452 dvss.n4068 dvss.n142 585
R1453 dvss.n181 dvss.n143 585
R1454 dvss.n4126 dvss.n147 585
R1455 dvss.n4125 dvss.n148 585
R1456 dvss.n185 dvss.n149 585
R1457 dvss.n186 dvss.n156 585
R1458 dvss.n4077 dvss.n186 585
R1459 dvss.n4118 dvss.n157 585
R1460 dvss.n4078 dvss.n157 585
R1461 dvss.n4117 dvss.n158 585
R1462 dvss.n4079 dvss.n158 585
R1463 dvss.n176 dvss.n159 585
R1464 dvss.n176 dvss.n175 585
R1465 dvss.n177 dvss.n167 585
R1466 dvss.n4087 dvss.n177 585
R1467 dvss.n4109 dvss.n168 585
R1468 dvss.n4088 dvss.n168 585
R1469 dvss.n4108 dvss.n169 585
R1470 dvss.n4090 dvss.n169 585
R1471 dvss.n4094 dvss.n170 585
R1472 dvss.n4094 dvss.n4093 585
R1473 dvss.n4097 dvss.n4096 585
R1474 dvss.n4096 dvss.n4095 585
R1475 dvss.n98 dvss.n97 585
R1476 dvss.n4188 dvss.n97 585
R1477 dvss.n4195 dvss.n4194 585
R1478 dvss.n4195 dvss.n96 585
R1479 dvss.n4196 dvss.n91 585
R1480 dvss.n4199 dvss.n4196 585
R1481 dvss.n4211 dvss.n92 585
R1482 dvss.n4198 dvss.n92 585
R1483 dvss.n4210 dvss.n81 585
R1484 dvss.n4197 dvss.n81 585
R1485 dvss.n4223 dvss.n82 585
R1486 dvss.n4223 dvss.n4222 585
R1487 dvss.n4224 dvss.n71 585
R1488 dvss.n4225 dvss.n4224 585
R1489 dvss.n4231 dvss.n72 585
R1490 dvss.n4227 dvss.n72 585
R1491 dvss.n4232 dvss.n66 585
R1492 dvss.n67 dvss.n66 585
R1493 dvss.n4238 dvss.n65 585
R1494 dvss.n4238 dvss.n4237 585
R1495 dvss.n4240 dvss.n4239 585
R1496 dvss.n4239 dvss.n57 585
R1497 dvss.n1019 dvss.n1018 585
R1498 dvss.n1018 dvss.n1017 585
R1499 dvss.n804 dvss.n803 585
R1500 dvss.n1015 dvss.n803 585
R1501 dvss.n1013 dvss.n835 585
R1502 dvss.n1014 dvss.n1013 585
R1503 dvss.n834 dvss.n833 585
R1504 dvss.n1016 dvss.n833 585
R1505 dvss.n1093 dvss.n786 585
R1506 dvss.n1096 dvss.n1095 585
R1507 dvss.n790 dvss.n789 585
R1508 dvss.n793 dvss.n790 585
R1509 dvss.n791 dvss.n779 585
R1510 dvss.n1114 dvss.n778 585
R1511 dvss.n1101 dvss.n1100 585
R1512 dvss.n1099 dvss.n782 585
R1513 dvss.n781 dvss.n780 585
R1514 dvss.n1103 dvss.n781 585
R1515 dvss.n1106 dvss.n1105 585
R1516 dvss.n775 dvss.n773 585
R1517 dvss.n1089 dvss.n1088 585
R1518 dvss.n1087 dvss.n802 585
R1519 dvss.n1086 dvss.n801 585
R1520 dvss.n1091 dvss.n801 585
R1521 dvss.n1085 dvss.n1084 585
R1522 dvss.n1083 dvss.n1082 585
R1523 dvss.n1081 dvss.n1080 585
R1524 dvss.n1079 dvss.n1078 585
R1525 dvss.n1077 dvss.n1076 585
R1526 dvss.n1075 dvss.n1074 585
R1527 dvss.n1073 dvss.n1072 585
R1528 dvss.n1071 dvss.n794 585
R1529 dvss.n1092 dvss.n795 585
R1530 dvss.n1092 dvss.n1091 585
R1531 dvss.n1050 dvss.n1049 585
R1532 dvss.n1048 dvss.n832 585
R1533 dvss.n1047 dvss.n831 585
R1534 dvss.n1052 dvss.n831 585
R1535 dvss.n1046 dvss.n1045 585
R1536 dvss.n1044 dvss.n1043 585
R1537 dvss.n1042 dvss.n1041 585
R1538 dvss.n1040 dvss.n1039 585
R1539 dvss.n1038 dvss.n1037 585
R1540 dvss.n1036 dvss.n1035 585
R1541 dvss.n827 dvss.n826 585
R1542 dvss.n1055 dvss.n1054 585
R1543 dvss.n784 dvss.n783 585
R1544 dvss.n1052 dvss.n783 585
R1545 dvss.n1010 dvss.n1009 585
R1546 dvss.n1011 dvss.n1010 585
R1547 dvss.n1008 dvss.n840 585
R1548 dvss.n840 dvss.n839 585
R1549 dvss.n1007 dvss.n1006 585
R1550 dvss.n1006 dvss.n1005 585
R1551 dvss.n844 dvss.n843 585
R1552 dvss.n1004 dvss.n844 585
R1553 dvss.n1002 dvss.n1001 585
R1554 dvss.n1003 dvss.n1002 585
R1555 dvss.n1000 dvss.n846 585
R1556 dvss.n846 dvss.n845 585
R1557 dvss.n999 dvss.n998 585
R1558 dvss.n998 dvss.n997 585
R1559 dvss.n852 dvss.n851 585
R1560 dvss.n996 dvss.n852 585
R1561 dvss.n993 dvss.n992 585
R1562 dvss.n994 dvss.n993 585
R1563 dvss.n991 dvss.n854 585
R1564 dvss.n864 dvss.n854 585
R1565 dvss.n990 dvss.n989 585
R1566 dvss.n989 dvss.n988 585
R1567 dvss.n863 dvss.n862 585
R1568 dvss.n987 dvss.n863 585
R1569 dvss.n985 dvss.n984 585
R1570 dvss.n986 dvss.n985 585
R1571 dvss.n983 dvss.n865 585
R1572 dvss.n877 dvss.n865 585
R1573 dvss.n982 dvss.n981 585
R1574 dvss.n981 dvss.n980 585
R1575 dvss.n876 dvss.n875 585
R1576 dvss.n979 dvss.n876 585
R1577 dvss.n977 dvss.n976 585
R1578 dvss.n978 dvss.n977 585
R1579 dvss.n975 dvss.n879 585
R1580 dvss.n879 dvss.n878 585
R1581 dvss.n974 dvss.n973 585
R1582 dvss.n973 dvss.n972 585
R1583 dvss.n3140 dvss.n2646 585
R1584 dvss.n3139 dvss.n2645 585
R1585 dvss.n3143 dvss.n2645 585
R1586 dvss.n3138 dvss.n3137 585
R1587 dvss.n3136 dvss.n3135 585
R1588 dvss.n3134 dvss.n3133 585
R1589 dvss.n3132 dvss.n3131 585
R1590 dvss.n3130 dvss.n3129 585
R1591 dvss.n3128 dvss.n3127 585
R1592 dvss.n3126 dvss.n3125 585
R1593 dvss.n3124 dvss.n3123 585
R1594 dvss.n3122 dvss.n3121 585
R1595 dvss.n3120 dvss.n3119 585
R1596 dvss.n3118 dvss.n3117 585
R1597 dvss.n3116 dvss.n3115 585
R1598 dvss.n3114 dvss.n3113 585
R1599 dvss.n3112 dvss.n3111 585
R1600 dvss.n3110 dvss.n3109 585
R1601 dvss.n3108 dvss.n3107 585
R1602 dvss.n3106 dvss.n3105 585
R1603 dvss.n3104 dvss.n3103 585
R1604 dvss.n3102 dvss.n3101 585
R1605 dvss.n3100 dvss.n3099 585
R1606 dvss.n3098 dvss.n3097 585
R1607 dvss.n3096 dvss.n3095 585
R1608 dvss.n3094 dvss.n3093 585
R1609 dvss.n3092 dvss.n3091 585
R1610 dvss.n3090 dvss.n3089 585
R1611 dvss.n3088 dvss.n3087 585
R1612 dvss.n3086 dvss.n3085 585
R1613 dvss.n3084 dvss.n3083 585
R1614 dvss.n3082 dvss.n3081 585
R1615 dvss.n3080 dvss.n3079 585
R1616 dvss.n3078 dvss.n3077 585
R1617 dvss.n3076 dvss.n3075 585
R1618 dvss.n3074 dvss.n3073 585
R1619 dvss.n3072 dvss.n3071 585
R1620 dvss.n3070 dvss.n3069 585
R1621 dvss.n3068 dvss.n3067 585
R1622 dvss.n3066 dvss.n3065 585
R1623 dvss.n3064 dvss.n3063 585
R1624 dvss.n3062 dvss.n3061 585
R1625 dvss.n3060 dvss.n3059 585
R1626 dvss.n3058 dvss.n3057 585
R1627 dvss.n3056 dvss.n3055 585
R1628 dvss.n3054 dvss.n3053 585
R1629 dvss.n3052 dvss.n3051 585
R1630 dvss.n3050 dvss.n3049 585
R1631 dvss.n3048 dvss.n3047 585
R1632 dvss.n3046 dvss.n3045 585
R1633 dvss.n3044 dvss.n3043 585
R1634 dvss.n3042 dvss.n3041 585
R1635 dvss.n3040 dvss.n3039 585
R1636 dvss.n3038 dvss.n3037 585
R1637 dvss.n3036 dvss.n3035 585
R1638 dvss.n3034 dvss.n3033 585
R1639 dvss.n3032 dvss.n3031 585
R1640 dvss.n3030 dvss.n3029 585
R1641 dvss.n3028 dvss.n3027 585
R1642 dvss.n3026 dvss.n3025 585
R1643 dvss.n3024 dvss.n3023 585
R1644 dvss.n3022 dvss.n3021 585
R1645 dvss.n3020 dvss.n3019 585
R1646 dvss.n3018 dvss.n3017 585
R1647 dvss.n3016 dvss.n3015 585
R1648 dvss.n3014 dvss.n3013 585
R1649 dvss.n3012 dvss.n3011 585
R1650 dvss.n3010 dvss.n3009 585
R1651 dvss.n3008 dvss.n3007 585
R1652 dvss.n3006 dvss.n3005 585
R1653 dvss.n3004 dvss.n3003 585
R1654 dvss.n3002 dvss.n3001 585
R1655 dvss.n3000 dvss.n2999 585
R1656 dvss.n2998 dvss.n2997 585
R1657 dvss.n2996 dvss.n2995 585
R1658 dvss.n2994 dvss.n2993 585
R1659 dvss.n2992 dvss.n2991 585
R1660 dvss.n2990 dvss.n2989 585
R1661 dvss.n2988 dvss.n2987 585
R1662 dvss.n2986 dvss.n2985 585
R1663 dvss.n2984 dvss.n2983 585
R1664 dvss.n2982 dvss.n2981 585
R1665 dvss.n2980 dvss.n2979 585
R1666 dvss.n2978 dvss.n2977 585
R1667 dvss.n2976 dvss.n2975 585
R1668 dvss.n2974 dvss.n2973 585
R1669 dvss.n2972 dvss.n2971 585
R1670 dvss.n2970 dvss.n2969 585
R1671 dvss.n2968 dvss.n2967 585
R1672 dvss.n2966 dvss.n2965 585
R1673 dvss.n2964 dvss.n2963 585
R1674 dvss.n2962 dvss.n2961 585
R1675 dvss.n2960 dvss.n2959 585
R1676 dvss.n2958 dvss.n2957 585
R1677 dvss.n2956 dvss.n2955 585
R1678 dvss.n2954 dvss.n2953 585
R1679 dvss.n2952 dvss.n2951 585
R1680 dvss.n2950 dvss.n2949 585
R1681 dvss.n2948 dvss.n2947 585
R1682 dvss.n2946 dvss.n2945 585
R1683 dvss.n2944 dvss.n2943 585
R1684 dvss.n2942 dvss.n2941 585
R1685 dvss.n2940 dvss.n2939 585
R1686 dvss.n2938 dvss.n2937 585
R1687 dvss.n2936 dvss.n2935 585
R1688 dvss.n2934 dvss.n2933 585
R1689 dvss.n2932 dvss.n2931 585
R1690 dvss.n2930 dvss.n2929 585
R1691 dvss.n2928 dvss.n2927 585
R1692 dvss.n2926 dvss.n2925 585
R1693 dvss.n2924 dvss.n2923 585
R1694 dvss.n2922 dvss.n2921 585
R1695 dvss.n2920 dvss.n2919 585
R1696 dvss.n2918 dvss.n2917 585
R1697 dvss.n2916 dvss.n2915 585
R1698 dvss.n2914 dvss.n2913 585
R1699 dvss.n2912 dvss.n2911 585
R1700 dvss.n2910 dvss.n2909 585
R1701 dvss.n2908 dvss.n2907 585
R1702 dvss.n2906 dvss.n2905 585
R1703 dvss.n2904 dvss.n2903 585
R1704 dvss.n2902 dvss.n2901 585
R1705 dvss.n2900 dvss.n2899 585
R1706 dvss.n2898 dvss.n2897 585
R1707 dvss.n2896 dvss.n2895 585
R1708 dvss.n2894 dvss.n2893 585
R1709 dvss.n2892 dvss.n2891 585
R1710 dvss.n2890 dvss.n2889 585
R1711 dvss.n2888 dvss.n2887 585
R1712 dvss.n2886 dvss.n2885 585
R1713 dvss.n2884 dvss.n2883 585
R1714 dvss.n2882 dvss.n2881 585
R1715 dvss.n2579 dvss.n2578 585
R1716 dvss.n3146 dvss.n3145 585
R1717 dvss.n2577 dvss.n2576 585
R1718 dvss.n2572 dvss.n2571 585
R1719 dvss.n2573 dvss.n2572 585
R1720 dvss.n2114 dvss.n2113 585
R1721 dvss.n2113 dvss.n2112 585
R1722 dvss.n2568 dvss.n2115 585
R1723 dvss.n2208 dvss.n2115 585
R1724 dvss.n2567 dvss.n2116 585
R1725 dvss.n2209 dvss.n2116 585
R1726 dvss.n2210 dvss.n2117 585
R1727 dvss.n2211 dvss.n2210 585
R1728 dvss.n2560 dvss.n2120 585
R1729 dvss.n2212 dvss.n2120 585
R1730 dvss.n2559 dvss.n2121 585
R1731 dvss.n2213 dvss.n2121 585
R1732 dvss.n2214 dvss.n2122 585
R1733 dvss.n2215 dvss.n2214 585
R1734 dvss.n2551 dvss.n2126 585
R1735 dvss.n2216 dvss.n2126 585
R1736 dvss.n2550 dvss.n2127 585
R1737 dvss.n2217 dvss.n2127 585
R1738 dvss.n2218 dvss.n2128 585
R1739 dvss.n2219 dvss.n2218 585
R1740 dvss.n2543 dvss.n2130 585
R1741 dvss.n2232 dvss.n2130 585
R1742 dvss.n2542 dvss.n2131 585
R1743 dvss.n2231 dvss.n2131 585
R1744 dvss.n2229 dvss.n2132 585
R1745 dvss.n2230 dvss.n2229 585
R1746 dvss.n2228 dvss.n2136 585
R1747 dvss.n2228 dvss.n2227 585
R1748 dvss.n2533 dvss.n2137 585
R1749 dvss.n2226 dvss.n2137 585
R1750 dvss.n2532 dvss.n2138 585
R1751 dvss.n2225 dvss.n2138 585
R1752 dvss.n2223 dvss.n2139 585
R1753 dvss.n2224 dvss.n2223 585
R1754 dvss.n2528 dvss.n2140 585
R1755 dvss.n2221 dvss.n2140 585
R1756 dvss.n2527 dvss.n2141 585
R1757 dvss.n2220 dvss.n2141 585
R1758 dvss.n2143 dvss.n2142 585
R1759 dvss.n2144 dvss.n2143 585
R1760 dvss.n2523 dvss.n2522 585
R1761 dvss.n2522 dvss.n2521 585
R1762 dvss.n4311 dvss.n57 583.256
R1763 dvss.n1014 dvss.n1012 578.14
R1764 dvss.n2364 dvss.t741 575.611
R1765 dvss.n2492 dvss.t679 568.053
R1766 dvss.n183 dvss.n180 564.282
R1767 dvss.n3821 dvss.n3818 564.282
R1768 dvss.n3675 dvss.n314 564.282
R1769 dvss.n3550 dvss.n3548 564.282
R1770 dvss.n3422 dvss.n443 564.282
R1771 dvss.n1648 dvss.n1645 564.282
R1772 dvss.n1474 dvss.n562 564.282
R1773 dvss.n728 dvss.n637 564.282
R1774 dvss.n2182 dvss.n2177 539.294
R1775 dvss.n2177 dvss.n2172 539.294
R1776 dvss.n2194 dvss.n2172 539.294
R1777 dvss.n2194 dvss.n2170 539.294
R1778 dvss.n2198 dvss.n2170 539.294
R1779 dvss.n2198 dvss.n2167 539.294
R1780 dvss.n2205 dvss.n2167 539.294
R1781 dvss.n2205 dvss.n2165 539.294
R1782 dvss.n2237 dvss.n2165 539.294
R1783 dvss.n2237 dvss.n2162 539.294
R1784 dvss.n2246 dvss.n2162 539.294
R1785 dvss.n2246 dvss.n2160 539.294
R1786 dvss.n2252 dvss.n2160 539.294
R1787 dvss.n2252 dvss.n2161 539.294
R1788 dvss.n2161 dvss.n2150 539.294
R1789 dvss.n2264 dvss.n2150 539.294
R1790 dvss.n2264 dvss.n2149 539.294
R1791 dvss.n2268 dvss.n2149 539.294
R1792 dvss.n2268 dvss.n2146 539.294
R1793 dvss.n2517 dvss.n2146 539.294
R1794 dvss.n2646 dvss.n2645 539.294
R1795 dvss.n3137 dvss.n2645 539.294
R1796 dvss.n3135 dvss.n3134 539.294
R1797 dvss.n3131 dvss.n3130 539.294
R1798 dvss.n3127 dvss.n3126 539.294
R1799 dvss.n3123 dvss.n3122 539.294
R1800 dvss.n3119 dvss.n3118 539.294
R1801 dvss.n3115 dvss.n3114 539.294
R1802 dvss.n3111 dvss.n3110 539.294
R1803 dvss.n3107 dvss.n3106 539.294
R1804 dvss.n3103 dvss.n3102 539.294
R1805 dvss.n3099 dvss.n3098 539.294
R1806 dvss.n3095 dvss.n3094 539.294
R1807 dvss.n3091 dvss.n3090 539.294
R1808 dvss.n3087 dvss.n3086 539.294
R1809 dvss.n3083 dvss.n3082 539.294
R1810 dvss.n3079 dvss.n3078 539.294
R1811 dvss.n3075 dvss.n3074 539.294
R1812 dvss.n3071 dvss.n3070 539.294
R1813 dvss.n3067 dvss.n3066 539.294
R1814 dvss.n3063 dvss.n3062 539.294
R1815 dvss.n3059 dvss.n3058 539.294
R1816 dvss.n3055 dvss.n3054 539.294
R1817 dvss.n3051 dvss.n3050 539.294
R1818 dvss.n3047 dvss.n3046 539.294
R1819 dvss.n3043 dvss.n3042 539.294
R1820 dvss.n3039 dvss.n3038 539.294
R1821 dvss.n3035 dvss.n3034 539.294
R1822 dvss.n3031 dvss.n3030 539.294
R1823 dvss.n3027 dvss.n3026 539.294
R1824 dvss.n3023 dvss.n3022 539.294
R1825 dvss.n3019 dvss.n3018 539.294
R1826 dvss.n3015 dvss.n3014 539.294
R1827 dvss.n3011 dvss.n3010 539.294
R1828 dvss.n3007 dvss.n3006 539.294
R1829 dvss.n3003 dvss.n3002 539.294
R1830 dvss.n2999 dvss.n2998 539.294
R1831 dvss.n2995 dvss.n2994 539.294
R1832 dvss.n2991 dvss.n2990 539.294
R1833 dvss.n2987 dvss.n2986 539.294
R1834 dvss.n2983 dvss.n2982 539.294
R1835 dvss.n2979 dvss.n2978 539.294
R1836 dvss.n2975 dvss.n2974 539.294
R1837 dvss.n2971 dvss.n2970 539.294
R1838 dvss.n2967 dvss.n2966 539.294
R1839 dvss.n2963 dvss.n2962 539.294
R1840 dvss.n2959 dvss.n2958 539.294
R1841 dvss.n2955 dvss.n2954 539.294
R1842 dvss.n2951 dvss.n2950 539.294
R1843 dvss.n2947 dvss.n2946 539.294
R1844 dvss.n2943 dvss.n2942 539.294
R1845 dvss.n2939 dvss.n2938 539.294
R1846 dvss.n2935 dvss.n2934 539.294
R1847 dvss.n2931 dvss.n2930 539.294
R1848 dvss.n2927 dvss.n2926 539.294
R1849 dvss.n2923 dvss.n2922 539.294
R1850 dvss.n2919 dvss.n2918 539.294
R1851 dvss.n2915 dvss.n2914 539.294
R1852 dvss.n2911 dvss.n2910 539.294
R1853 dvss.n2907 dvss.n2906 539.294
R1854 dvss.n2903 dvss.n2902 539.294
R1855 dvss.n2899 dvss.n2898 539.294
R1856 dvss.n2895 dvss.n2894 539.294
R1857 dvss.n2891 dvss.n2890 539.294
R1858 dvss.n2887 dvss.n2886 539.294
R1859 dvss.n2883 dvss.n2882 539.294
R1860 dvss.n3145 dvss.n2579 539.294
R1861 dvss.n3152 dvss.n2576 539.294
R1862 dvss.n3152 dvss.n2110 539.294
R1863 dvss.n3156 dvss.n2110 539.294
R1864 dvss.n3156 dvss.n2107 539.294
R1865 dvss.n3165 dvss.n2107 539.294
R1866 dvss.n3165 dvss.n2104 539.294
R1867 dvss.n3171 dvss.n2104 539.294
R1868 dvss.n3171 dvss.n2105 539.294
R1869 dvss.n2105 dvss.n2094 539.294
R1870 dvss.n3183 dvss.n2094 539.294
R1871 dvss.n3183 dvss.n2093 539.294
R1872 dvss.n3188 dvss.n2093 539.294
R1873 dvss.n3188 dvss.n2090 539.294
R1874 dvss.n3195 dvss.n2090 539.294
R1875 dvss.n3195 dvss.n2088 539.294
R1876 dvss.n3200 dvss.n2088 539.294
R1877 dvss.n3200 dvss.n2084 539.294
R1878 dvss.n3211 dvss.n2084 539.294
R1879 dvss.n3211 dvss.n2083 539.294
R1880 dvss.n3215 dvss.n2083 539.294
R1881 dvss.n3215 dvss.n2080 539.294
R1882 dvss.n3222 dvss.n2080 539.294
R1883 dvss.n3222 dvss.n2078 539.294
R1884 dvss.n3227 dvss.n2078 539.294
R1885 dvss.n3227 dvss.n1998 539.294
R1886 dvss.n3236 dvss.n1998 539.294
R1887 dvss.n3236 dvss.n1999 539.294
R1888 dvss.n2014 dvss.n1999 539.294
R1889 dvss.n2014 dvss.n2008 539.294
R1890 dvss.n2024 dvss.n2008 539.294
R1891 dvss.n2024 dvss.n2006 539.294
R1892 dvss.n2028 dvss.n2006 539.294
R1893 dvss.n2029 dvss.n2028 539.294
R1894 dvss.n2030 dvss.n2029 539.294
R1895 dvss.n2041 dvss.n2030 539.294
R1896 dvss.n2041 dvss.n2032 539.294
R1897 dvss.n2033 dvss.n2032 539.294
R1898 dvss.n2037 dvss.n2033 539.294
R1899 dvss.n2057 dvss.n2037 539.294
R1900 dvss.n2057 dvss.n2038 539.294
R1901 dvss.n2038 dvss.n11 539.294
R1902 dvss.n12 dvss.n11 539.294
R1903 dvss.n2051 dvss.n12 539.294
R1904 dvss.n2051 dvss.n14 539.294
R1905 dvss.n15 dvss.n14 539.294
R1906 dvss.n2047 dvss.n15 539.294
R1907 dvss.n2047 dvss.n17 539.294
R1908 dvss.n18 dvss.n17 539.294
R1909 dvss.n120 dvss.n18 539.294
R1910 dvss.n120 dvss.n119 539.294
R1911 dvss.n119 dvss.n107 539.294
R1912 dvss.n107 dvss.n101 539.294
R1913 dvss.n4156 dvss.n101 539.294
R1914 dvss.n4157 dvss.n4156 539.294
R1915 dvss.n4157 dvss.n24 539.294
R1916 dvss.n25 dvss.n24 539.294
R1917 dvss.n4161 dvss.n25 539.294
R1918 dvss.n4161 dvss.n27 539.294
R1919 dvss.n28 dvss.n27 539.294
R1920 dvss.n4166 dvss.n28 539.294
R1921 dvss.n4167 dvss.n4166 539.294
R1922 dvss.n4167 dvss.n34 539.294
R1923 dvss.n35 dvss.n34 539.294
R1924 dvss.n4171 dvss.n35 539.294
R1925 dvss.n4171 dvss.n37 539.294
R1926 dvss.n38 dvss.n37 539.294
R1927 dvss.n4175 dvss.n38 539.294
R1928 dvss.n4175 dvss.n40 539.294
R1929 dvss.n41 dvss.n40 539.294
R1930 dvss.n4183 dvss.n41 539.294
R1931 dvss.n4183 dvss.n45 539.294
R1932 dvss.n46 dvss.n45 539.294
R1933 dvss.n4179 dvss.n46 539.294
R1934 dvss.n4179 dvss.n49 539.294
R1935 dvss.n50 dvss.n49 539.294
R1936 dvss.n78 dvss.n50 539.294
R1937 dvss.n78 dvss.n52 539.294
R1938 dvss.n53 dvss.n52 539.294
R1939 dvss.n55 dvss.n53 539.294
R1940 dvss.n4313 dvss.n55 539.294
R1941 dvss.n1013 dvss.n833 539.294
R1942 dvss.n1050 dvss.n833 539.294
R1943 dvss.n832 dvss.n831 539.294
R1944 dvss.n1045 dvss.n831 539.294
R1945 dvss.n1043 dvss.n1042 539.294
R1946 dvss.n1039 dvss.n1038 539.294
R1947 dvss.n1035 dvss.n827 539.294
R1948 dvss.n1054 dvss.n783 539.294
R1949 dvss.n1101 dvss.n783 539.294
R1950 dvss.n782 dvss.n781 539.294
R1951 dvss.n1105 dvss.n781 539.294
R1952 dvss.n1118 dvss.n775 539.294
R1953 dvss.n1118 dvss.n770 539.294
R1954 dvss.n1127 dvss.n770 539.294
R1955 dvss.n1128 dvss.n1127 539.294
R1956 dvss.n1128 dvss.n760 539.294
R1957 dvss.n1141 dvss.n760 539.294
R1958 dvss.n1147 dvss.n1141 539.294
R1959 dvss.n1147 dvss.n1146 539.294
R1960 dvss.n1146 dvss.n750 539.294
R1961 dvss.n1164 dvss.n750 539.294
R1962 dvss.n1164 dvss.n742 539.294
R1963 dvss.n1179 dvss.n742 539.294
R1964 dvss.n1180 dvss.n1179 539.294
R1965 dvss.n1180 dvss.n741 539.294
R1966 dvss.n1185 dvss.n741 539.294
R1967 dvss.n1185 dvss.n628 539.294
R1968 dvss.n1264 dvss.n628 539.294
R1969 dvss.n1264 dvss.n629 539.294
R1970 dvss.n1260 dvss.n629 539.294
R1971 dvss.n1208 dvss.n635 539.294
R1972 dvss.n1255 dvss.n639 539.294
R1973 dvss.n1255 dvss.n640 539.294
R1974 dvss.n1251 dvss.n640 539.294
R1975 dvss.n1251 dvss.n646 539.294
R1976 dvss.n1247 dvss.n646 539.294
R1977 dvss.n1247 dvss.n650 539.294
R1978 dvss.n1243 dvss.n650 539.294
R1979 dvss.n1243 dvss.n655 539.294
R1980 dvss.n682 dvss.n655 539.294
R1981 dvss.n689 dvss.n682 539.294
R1982 dvss.n690 dvss.n689 539.294
R1983 dvss.n690 dvss.n679 539.294
R1984 dvss.n696 dvss.n679 539.294
R1985 dvss.n697 dvss.n696 539.294
R1986 dvss.n697 dvss.n580 539.294
R1987 dvss.n1462 dvss.n580 539.294
R1988 dvss.n1462 dvss.n566 539.294
R1989 dvss.n1489 dvss.n566 539.294
R1990 dvss.n1489 dvss.n567 539.294
R1991 dvss.n1478 dvss.n567 539.294
R1992 dvss.n1480 dvss.n1477 539.294
R1993 dvss.n1477 dvss.n556 539.294
R1994 dvss.n1504 dvss.n556 539.294
R1995 dvss.n1504 dvss.n552 539.294
R1996 dvss.n1517 dvss.n552 539.294
R1997 dvss.n1518 dvss.n1517 539.294
R1998 dvss.n1518 dvss.n546 539.294
R1999 dvss.n546 dvss.n541 539.294
R2000 dvss.n1541 dvss.n541 539.294
R2001 dvss.n1542 dvss.n1541 539.294
R2002 dvss.n1542 dvss.n537 539.294
R2003 dvss.n537 dvss.n531 539.294
R2004 dvss.n1566 dvss.n531 539.294
R2005 dvss.n1567 dvss.n1566 539.294
R2006 dvss.n1567 dvss.n530 539.294
R2007 dvss.n1572 dvss.n530 539.294
R2008 dvss.n1572 dvss.n508 539.294
R2009 dvss.n1747 dvss.n508 539.294
R2010 dvss.n1747 dvss.n509 539.294
R2011 dvss.n1654 dvss.n509 539.294
R2012 dvss.n1653 dvss.n1652 539.294
R2013 dvss.n1660 dvss.n1658 539.294
R2014 dvss.n1660 dvss.n1643 539.294
R2015 dvss.n1664 dvss.n1643 539.294
R2016 dvss.n1665 dvss.n1664 539.294
R2017 dvss.n1670 dvss.n1665 539.294
R2018 dvss.n1670 dvss.n1639 539.294
R2019 dvss.n1675 dvss.n1639 539.294
R2020 dvss.n1676 dvss.n1675 539.294
R2021 dvss.n1676 dvss.n1637 539.294
R2022 dvss.n1683 dvss.n1637 539.294
R2023 dvss.n1684 dvss.n1683 539.294
R2024 dvss.n1684 dvss.n1634 539.294
R2025 dvss.n1690 dvss.n1634 539.294
R2026 dvss.n1691 dvss.n1690 539.294
R2027 dvss.n1691 dvss.n460 539.294
R2028 dvss.n3411 dvss.n460 539.294
R2029 dvss.n3411 dvss.n447 539.294
R2030 dvss.n3440 dvss.n447 539.294
R2031 dvss.n3440 dvss.n448 539.294
R2032 dvss.n3431 dvss.n3428 539.294
R2033 dvss.n3429 dvss.n437 539.294
R2034 dvss.n3455 dvss.n437 539.294
R2035 dvss.n3455 dvss.n433 539.294
R2036 dvss.n3468 dvss.n433 539.294
R2037 dvss.n3469 dvss.n3468 539.294
R2038 dvss.n3469 dvss.n427 539.294
R2039 dvss.n427 dvss.n422 539.294
R2040 dvss.n3492 dvss.n422 539.294
R2041 dvss.n3493 dvss.n3492 539.294
R2042 dvss.n3493 dvss.n418 539.294
R2043 dvss.n418 dvss.n412 539.294
R2044 dvss.n3517 dvss.n412 539.294
R2045 dvss.n3518 dvss.n3517 539.294
R2046 dvss.n3518 dvss.n411 539.294
R2047 dvss.n3524 dvss.n411 539.294
R2048 dvss.n3524 dvss.n390 539.294
R2049 dvss.n3541 dvss.n390 539.294
R2050 dvss.n3541 dvss.n384 539.294
R2051 dvss.n3560 dvss.n384 539.294
R2052 dvss.n383 dvss.n380 539.294
R2053 dvss.n3564 dvss.n373 539.294
R2054 dvss.n3577 dvss.n373 539.294
R2055 dvss.n3577 dvss.n370 539.294
R2056 dvss.n3584 dvss.n370 539.294
R2057 dvss.n3584 dvss.n363 539.294
R2058 dvss.n3603 dvss.n363 539.294
R2059 dvss.n3603 dvss.n358 539.294
R2060 dvss.n3608 dvss.n358 539.294
R2061 dvss.n3608 dvss.n352 539.294
R2062 dvss.n3620 dvss.n352 539.294
R2063 dvss.n3620 dvss.n347 539.294
R2064 dvss.n3634 dvss.n347 539.294
R2065 dvss.n3634 dvss.n343 539.294
R2066 dvss.n3641 dvss.n343 539.294
R2067 dvss.n3641 dvss.n344 539.294
R2068 dvss.n344 dvss.n332 539.294
R2069 dvss.n332 dvss.n325 539.294
R2070 dvss.n3662 dvss.n325 539.294
R2071 dvss.n3663 dvss.n3662 539.294
R2072 dvss.n3667 dvss.n321 539.294
R2073 dvss.n322 dvss.n311 539.294
R2074 dvss.n311 dvss.n306 539.294
R2075 dvss.n3699 dvss.n306 539.294
R2076 dvss.n3700 dvss.n3699 539.294
R2077 dvss.n3700 dvss.n295 539.294
R2078 dvss.n3719 dvss.n295 539.294
R2079 dvss.n3719 dvss.n291 539.294
R2080 dvss.n3724 dvss.n291 539.294
R2081 dvss.n3725 dvss.n3724 539.294
R2082 dvss.n3725 dvss.n287 539.294
R2083 dvss.n287 dvss.n281 539.294
R2084 dvss.n3749 dvss.n281 539.294
R2085 dvss.n3750 dvss.n3749 539.294
R2086 dvss.n3750 dvss.n280 539.294
R2087 dvss.n3755 dvss.n280 539.294
R2088 dvss.n3755 dvss.n263 539.294
R2089 dvss.n3878 dvss.n263 539.294
R2090 dvss.n3878 dvss.n264 539.294
R2091 dvss.n3814 dvss.n264 539.294
R2092 dvss.n3813 dvss.n3812 539.294
R2093 dvss.n3810 dvss.n3809 539.294
R2094 dvss.n3827 dvss.n3809 539.294
R2095 dvss.n3828 dvss.n3827 539.294
R2096 dvss.n3828 dvss.n3803 539.294
R2097 dvss.n3834 dvss.n3803 539.294
R2098 dvss.n3835 dvss.n3834 539.294
R2099 dvss.n3835 dvss.n3798 539.294
R2100 dvss.n3840 dvss.n3798 539.294
R2101 dvss.n3840 dvss.n123 539.294
R2102 dvss.n4150 dvss.n123 539.294
R2103 dvss.n4150 dvss.n124 539.294
R2104 dvss.n195 dvss.n124 539.294
R2105 dvss.n202 dvss.n195 539.294
R2106 dvss.n206 dvss.n202 539.294
R2107 dvss.n206 dvss.n191 539.294
R2108 dvss.n214 dvss.n191 539.294
R2109 dvss.n214 dvss.n189 539.294
R2110 dvss.n4069 dvss.n189 539.294
R2111 dvss.n4070 dvss.n4069 539.294
R2112 dvss.n188 dvss.n187 539.294
R2113 dvss.n4076 dvss.n4074 539.294
R2114 dvss.n4076 dvss.n178 539.294
R2115 dvss.n4080 dvss.n178 539.294
R2116 dvss.n4081 dvss.n4080 539.294
R2117 dvss.n4086 dvss.n4081 539.294
R2118 dvss.n4086 dvss.n174 539.294
R2119 dvss.n4091 dvss.n174 539.294
R2120 dvss.n4092 dvss.n4091 539.294
R2121 dvss.n4092 dvss.n100 539.294
R2122 dvss.n4189 dvss.n100 539.294
R2123 dvss.n4189 dvss.n94 539.294
R2124 dvss.n4200 dvss.n94 539.294
R2125 dvss.n4200 dvss.n95 539.294
R2126 dvss.n95 dvss.n83 539.294
R2127 dvss.n4221 dvss.n83 539.294
R2128 dvss.n4221 dvss.n75 539.294
R2129 dvss.n4228 dvss.n75 539.294
R2130 dvss.n4228 dvss.n68 539.294
R2131 dvss.n4236 dvss.n68 539.294
R2132 dvss.n4236 dvss.n69 539.294
R2133 dvss.n1010 dvss.n840 539.294
R2134 dvss.n1006 dvss.n840 539.294
R2135 dvss.n1006 dvss.n844 539.294
R2136 dvss.n1002 dvss.n844 539.294
R2137 dvss.n1002 dvss.n846 539.294
R2138 dvss.n998 dvss.n846 539.294
R2139 dvss.n998 dvss.n852 539.294
R2140 dvss.n993 dvss.n852 539.294
R2141 dvss.n993 dvss.n854 539.294
R2142 dvss.n989 dvss.n854 539.294
R2143 dvss.n989 dvss.n863 539.294
R2144 dvss.n985 dvss.n863 539.294
R2145 dvss.n985 dvss.n865 539.294
R2146 dvss.n981 dvss.n865 539.294
R2147 dvss.n981 dvss.n876 539.294
R2148 dvss.n977 dvss.n876 539.294
R2149 dvss.n973 dvss.n879 539.294
R2150 dvss.n973 dvss.n889 539.294
R2151 dvss.n969 dvss.n889 539.294
R2152 dvss.n969 dvss.n890 539.294
R2153 dvss.n965 dvss.n890 539.294
R2154 dvss.n965 dvss.n896 539.294
R2155 dvss.n961 dvss.n896 539.294
R2156 dvss.n961 dvss.n898 539.294
R2157 dvss.n957 dvss.n898 539.294
R2158 dvss.n957 dvss.n954 539.294
R2159 dvss.n954 dvss.n903 539.294
R2160 dvss.n950 dvss.n903 539.294
R2161 dvss.n950 dvss.n905 539.294
R2162 dvss.n946 dvss.n905 539.294
R2163 dvss.n946 dvss.n930 539.294
R2164 dvss.n942 dvss.n930 539.294
R2165 dvss.n942 dvss.n623 539.294
R2166 dvss.n1270 dvss.n623 539.294
R2167 dvss.n1270 dvss.n620 539.294
R2168 dvss.n1277 dvss.n620 539.294
R2169 dvss.n1281 dvss.n619 539.294
R2170 dvss.n1289 dvss.n616 539.294
R2171 dvss.n1289 dvss.n614 539.294
R2172 dvss.n1293 dvss.n614 539.294
R2173 dvss.n1293 dvss.n608 539.294
R2174 dvss.n1304 dvss.n608 539.294
R2175 dvss.n1304 dvss.n606 539.294
R2176 dvss.n1309 dvss.n606 539.294
R2177 dvss.n1309 dvss.n598 539.294
R2178 dvss.n1319 dvss.n598 539.294
R2179 dvss.n1319 dvss.n597 539.294
R2180 dvss.n1324 dvss.n597 539.294
R2181 dvss.n1324 dvss.n590 539.294
R2182 dvss.n1334 dvss.n590 539.294
R2183 dvss.n1334 dvss.n589 539.294
R2184 dvss.n1338 dvss.n589 539.294
R2185 dvss.n1338 dvss.n584 539.294
R2186 dvss.n1457 dvss.n584 539.294
R2187 dvss.n1457 dvss.n585 539.294
R2188 dvss.n1347 dvss.n585 539.294
R2189 dvss.n1375 dvss.n1348 539.294
R2190 dvss.n1351 dvss.n1350 539.294
R2191 dvss.n1382 dvss.n1351 539.294
R2192 dvss.n1383 dvss.n1382 539.294
R2193 dvss.n1383 dvss.n1356 539.294
R2194 dvss.n1357 dvss.n1356 539.294
R2195 dvss.n1374 dvss.n1357 539.294
R2196 dvss.n1374 dvss.n1362 539.294
R2197 dvss.n1363 dvss.n1362 539.294
R2198 dvss.n1392 dvss.n1363 539.294
R2199 dvss.n1392 dvss.n1366 539.294
R2200 dvss.n1367 dvss.n1366 539.294
R2201 dvss.n1397 dvss.n1367 539.294
R2202 dvss.n1398 dvss.n1397 539.294
R2203 dvss.n1398 dvss.n1373 539.294
R2204 dvss.n1402 dvss.n1373 539.294
R2205 dvss.n1402 dvss.n503 539.294
R2206 dvss.n1753 dvss.n503 539.294
R2207 dvss.n1753 dvss.n500 539.294
R2208 dvss.n1760 dvss.n500 539.294
R2209 dvss.n1764 dvss.n499 539.294
R2210 dvss.n1772 dvss.n496 539.294
R2211 dvss.n1772 dvss.n494 539.294
R2212 dvss.n1776 dvss.n494 539.294
R2213 dvss.n1776 dvss.n488 539.294
R2214 dvss.n1787 dvss.n488 539.294
R2215 dvss.n1787 dvss.n486 539.294
R2216 dvss.n1792 dvss.n486 539.294
R2217 dvss.n1792 dvss.n478 539.294
R2218 dvss.n1802 dvss.n478 539.294
R2219 dvss.n1802 dvss.n477 539.294
R2220 dvss.n1807 dvss.n477 539.294
R2221 dvss.n1807 dvss.n470 539.294
R2222 dvss.n1817 dvss.n470 539.294
R2223 dvss.n1817 dvss.n469 539.294
R2224 dvss.n1821 dvss.n469 539.294
R2225 dvss.n1821 dvss.n464 539.294
R2226 dvss.n3406 dvss.n464 539.294
R2227 dvss.n3406 dvss.n465 539.294
R2228 dvss.n1830 dvss.n465 539.294
R2229 dvss.n1932 dvss.n1831 539.294
R2230 dvss.n1834 dvss.n1833 539.294
R2231 dvss.n1939 dvss.n1834 539.294
R2232 dvss.n1940 dvss.n1939 539.294
R2233 dvss.n1940 dvss.n1839 539.294
R2234 dvss.n1840 dvss.n1839 539.294
R2235 dvss.n1931 dvss.n1840 539.294
R2236 dvss.n1931 dvss.n1845 539.294
R2237 dvss.n1846 dvss.n1845 539.294
R2238 dvss.n1949 dvss.n1846 539.294
R2239 dvss.n1949 dvss.n1849 539.294
R2240 dvss.n1850 dvss.n1849 539.294
R2241 dvss.n1954 dvss.n1850 539.294
R2242 dvss.n1955 dvss.n1954 539.294
R2243 dvss.n1955 dvss.n1856 539.294
R2244 dvss.n1857 dvss.n1856 539.294
R2245 dvss.n1959 dvss.n1857 539.294
R2246 dvss.n1959 dvss.n1859 539.294
R2247 dvss.n1860 dvss.n1859 539.294
R2248 dvss.n1928 dvss.n1860 539.294
R2249 dvss.n1863 dvss.n1862 539.294
R2250 dvss.n1926 dvss.n1865 539.294
R2251 dvss.n1866 dvss.n1865 539.294
R2252 dvss.n1967 dvss.n1866 539.294
R2253 dvss.n1967 dvss.n1870 539.294
R2254 dvss.n1871 dvss.n1870 539.294
R2255 dvss.n1925 dvss.n1871 539.294
R2256 dvss.n1925 dvss.n1876 539.294
R2257 dvss.n1877 dvss.n1876 539.294
R2258 dvss.n1974 dvss.n1877 539.294
R2259 dvss.n1974 dvss.n1880 539.294
R2260 dvss.n1881 dvss.n1880 539.294
R2261 dvss.n1979 dvss.n1881 539.294
R2262 dvss.n1980 dvss.n1979 539.294
R2263 dvss.n1980 dvss.n1887 539.294
R2264 dvss.n1888 dvss.n1887 539.294
R2265 dvss.n1984 dvss.n1888 539.294
R2266 dvss.n1984 dvss.n1890 539.294
R2267 dvss.n1891 dvss.n1890 539.294
R2268 dvss.n1922 dvss.n1891 539.294
R2269 dvss.n1894 dvss.n1893 539.294
R2270 dvss.n1920 dvss.n1896 539.294
R2271 dvss.n1897 dvss.n1896 539.294
R2272 dvss.n1992 dvss.n1897 539.294
R2273 dvss.n1992 dvss.n1901 539.294
R2274 dvss.n1902 dvss.n1901 539.294
R2275 dvss.n1919 dvss.n1902 539.294
R2276 dvss.n1919 dvss.n1907 539.294
R2277 dvss.n1908 dvss.n1907 539.294
R2278 dvss.n3241 dvss.n1908 539.294
R2279 dvss.n3241 dvss.n1911 539.294
R2280 dvss.n1912 dvss.n1911 539.294
R2281 dvss.n3246 dvss.n1912 539.294
R2282 dvss.n3247 dvss.n3246 539.294
R2283 dvss.n3247 dvss.n1918 539.294
R2284 dvss.n3251 dvss.n1918 539.294
R2285 dvss.n3251 dvss.n257 539.294
R2286 dvss.n3884 dvss.n257 539.294
R2287 dvss.n3884 dvss.n254 539.294
R2288 dvss.n3891 dvss.n254 539.294
R2289 dvss.n3895 dvss.n253 539.294
R2290 dvss.n3903 dvss.n250 539.294
R2291 dvss.n3903 dvss.n248 539.294
R2292 dvss.n3907 dvss.n248 539.294
R2293 dvss.n3907 dvss.n242 539.294
R2294 dvss.n3918 dvss.n242 539.294
R2295 dvss.n3918 dvss.n240 539.294
R2296 dvss.n3923 dvss.n240 539.294
R2297 dvss.n3923 dvss.n232 539.294
R2298 dvss.n3933 dvss.n232 539.294
R2299 dvss.n3933 dvss.n231 539.294
R2300 dvss.n3938 dvss.n231 539.294
R2301 dvss.n3938 dvss.n224 539.294
R2302 dvss.n3948 dvss.n224 539.294
R2303 dvss.n3948 dvss.n223 539.294
R2304 dvss.n3952 dvss.n223 539.294
R2305 dvss.n3952 dvss.n218 539.294
R2306 dvss.n4063 dvss.n218 539.294
R2307 dvss.n4063 dvss.n219 539.294
R2308 dvss.n3956 dvss.n219 539.294
R2309 dvss.n3973 dvss.n3957 539.294
R2310 dvss.n3960 dvss.n3959 539.294
R2311 dvss.n3980 dvss.n3960 539.294
R2312 dvss.n3981 dvss.n3980 539.294
R2313 dvss.n3981 dvss.n3965 539.294
R2314 dvss.n3966 dvss.n3965 539.294
R2315 dvss.n3972 dvss.n3966 539.294
R2316 dvss.n3972 dvss.n3971 539.294
R2317 dvss.n3988 dvss.n3971 539.294
R2318 dvss.n4000 dvss.n3988 539.294
R2319 dvss.n4000 dvss.n3991 539.294
R2320 dvss.n3992 dvss.n3991 539.294
R2321 dvss.n4005 dvss.n3992 539.294
R2322 dvss.n4006 dvss.n4005 539.294
R2323 dvss.n4006 dvss.n3998 539.294
R2324 dvss.n3999 dvss.n3998 539.294
R2325 dvss.n4011 dvss.n3999 539.294
R2326 dvss.n4011 dvss.n60 539.294
R2327 dvss.n4308 dvss.n60 539.294
R2328 dvss.n4308 dvss.n61 539.294
R2329 dvss.n1018 dvss.n803 539.294
R2330 dvss.n1089 dvss.n803 539.294
R2331 dvss.n802 dvss.n801 539.294
R2332 dvss.n1084 dvss.n801 539.294
R2333 dvss.n1082 dvss.n1081 539.294
R2334 dvss.n1078 dvss.n1077 539.294
R2335 dvss.n1074 dvss.n1073 539.294
R2336 dvss.n1092 dvss.n794 539.294
R2337 dvss.n1093 dvss.n1092 539.294
R2338 dvss.n1095 dvss.n790 539.294
R2339 dvss.n1116 dvss.n778 539.294
R2340 dvss.n1116 dvss.n771 539.294
R2341 dvss.n1125 dvss.n771 539.294
R2342 dvss.n1125 dvss.n763 539.294
R2343 dvss.n1138 dvss.n763 539.294
R2344 dvss.n1138 dvss.n758 539.294
R2345 dvss.n1149 dvss.n758 539.294
R2346 dvss.n1149 dvss.n751 539.294
R2347 dvss.n1160 dvss.n751 539.294
R2348 dvss.n1160 dvss.n745 539.294
R2349 dvss.n1176 dvss.n745 539.294
R2350 dvss.n1177 dvss.n1176 539.294
R2351 dvss.n1177 dvss.n738 539.294
R2352 dvss.n739 dvss.n738 539.294
R2353 dvss.n1183 dvss.n739 539.294
R2354 dvss.n1183 dvss.n730 539.294
R2355 dvss.n730 dvss.n626 539.294
R2356 dvss.n1202 dvss.n626 539.294
R2357 dvss.n1203 dvss.n1202 539.294
R2358 dvss.n1205 dvss.n726 539.294
R2359 dvss.n724 dvss.n638 539.294
R2360 dvss.n1220 dvss.n638 539.294
R2361 dvss.n1220 dvss.n647 539.294
R2362 dvss.n648 dvss.n647 539.294
R2363 dvss.n649 dvss.n648 539.294
R2364 dvss.n658 dvss.n649 539.294
R2365 dvss.n1241 dvss.n658 539.294
R2366 dvss.n1241 dvss.n659 539.294
R2367 dvss.n685 dvss.n659 539.294
R2368 dvss.n685 dvss.n665 539.294
R2369 dvss.n666 dvss.n665 539.294
R2370 dvss.n693 dvss.n666 539.294
R2371 dvss.n694 dvss.n693 539.294
R2372 dvss.n694 dvss.n678 539.294
R2373 dvss.n700 dvss.n678 539.294
R2374 dvss.n700 dvss.n581 539.294
R2375 dvss.n581 dvss.n572 539.294
R2376 dvss.n572 dvss.n565 539.294
R2377 dvss.n1471 dvss.n565 539.294
R2378 dvss.n1476 dvss.n1472 539.294
R2379 dvss.n1493 dvss.n561 539.294
R2380 dvss.n1493 dvss.n555 539.294
R2381 dvss.n1507 dvss.n555 539.294
R2382 dvss.n1507 dvss.n549 539.294
R2383 dvss.n1520 dvss.n549 539.294
R2384 dvss.n1520 dvss.n543 539.294
R2385 dvss.n1536 dvss.n543 539.294
R2386 dvss.n1536 dvss.n540 539.294
R2387 dvss.n1544 dvss.n540 539.294
R2388 dvss.n1544 dvss.n534 539.294
R2389 dvss.n1563 dvss.n534 539.294
R2390 dvss.n1564 dvss.n1563 539.294
R2391 dvss.n1564 dvss.n527 539.294
R2392 dvss.n528 dvss.n527 539.294
R2393 dvss.n1570 dvss.n528 539.294
R2394 dvss.n1570 dvss.n514 539.294
R2395 dvss.n514 dvss.n506 539.294
R2396 dvss.n1586 dvss.n506 539.294
R2397 dvss.n1646 dvss.n1586 539.294
R2398 dvss.n1591 dvss.n1590 539.294
R2399 dvss.n1651 dvss.n1650 539.294
R2400 dvss.n1651 dvss.n1600 539.294
R2401 dvss.n1601 dvss.n1600 539.294
R2402 dvss.n1641 dvss.n1601 539.294
R2403 dvss.n1642 dvss.n1641 539.294
R2404 dvss.n1642 dvss.n1611 539.294
R2405 dvss.n1612 dvss.n1611 539.294
R2406 dvss.n1678 dvss.n1612 539.294
R2407 dvss.n1679 dvss.n1678 539.294
R2408 dvss.n1679 dvss.n1620 539.294
R2409 dvss.n1621 dvss.n1620 539.294
R2410 dvss.n1687 dvss.n1621 539.294
R2411 dvss.n1688 dvss.n1687 539.294
R2412 dvss.n1688 dvss.n1633 539.294
R2413 dvss.n1694 dvss.n1633 539.294
R2414 dvss.n1694 dvss.n461 539.294
R2415 dvss.n461 dvss.n452 539.294
R2416 dvss.n452 dvss.n446 539.294
R2417 dvss.n3419 dvss.n446 539.294
R2418 dvss.n3424 dvss.n3420 539.294
R2419 dvss.n3444 dvss.n442 539.294
R2420 dvss.n3444 dvss.n436 539.294
R2421 dvss.n3458 dvss.n436 539.294
R2422 dvss.n3458 dvss.n430 539.294
R2423 dvss.n3471 dvss.n430 539.294
R2424 dvss.n3471 dvss.n424 539.294
R2425 dvss.n3487 dvss.n424 539.294
R2426 dvss.n3487 dvss.n421 539.294
R2427 dvss.n3495 dvss.n421 539.294
R2428 dvss.n3495 dvss.n415 539.294
R2429 dvss.n3514 dvss.n415 539.294
R2430 dvss.n3515 dvss.n3514 539.294
R2431 dvss.n3515 dvss.n408 539.294
R2432 dvss.n409 dvss.n408 539.294
R2433 dvss.n3521 dvss.n409 539.294
R2434 dvss.n3521 dvss.n395 539.294
R2435 dvss.n395 dvss.n388 539.294
R2436 dvss.n3544 dvss.n388 539.294
R2437 dvss.n3545 dvss.n3544 539.294
R2438 dvss.n3552 dvss.n3546 539.294
R2439 dvss.n3547 dvss.n378 539.294
R2440 dvss.n378 dvss.n371 539.294
R2441 dvss.n3580 dvss.n371 539.294
R2442 dvss.n3581 dvss.n3580 539.294
R2443 dvss.n3581 dvss.n366 539.294
R2444 dvss.n366 dvss.n362 539.294
R2445 dvss.n362 dvss.n361 539.294
R2446 dvss.n361 dvss.n356 539.294
R2447 dvss.n356 dvss.n350 539.294
R2448 dvss.n3622 dvss.n350 539.294
R2449 dvss.n3623 dvss.n3622 539.294
R2450 dvss.n3623 dvss.n346 539.294
R2451 dvss.n346 dvss.n340 539.294
R2452 dvss.n341 dvss.n340 539.294
R2453 dvss.n3637 dvss.n341 539.294
R2454 dvss.n3637 dvss.n328 539.294
R2455 dvss.n3659 dvss.n328 539.294
R2456 dvss.n3659 dvss.n316 539.294
R2457 dvss.n3673 dvss.n316 539.294
R2458 dvss.n315 dvss.n313 539.294
R2459 dvss.n3677 dvss.n308 539.294
R2460 dvss.n3696 dvss.n308 539.294
R2461 dvss.n3696 dvss.n303 539.294
R2462 dvss.n3702 dvss.n303 539.294
R2463 dvss.n3702 dvss.n304 539.294
R2464 dvss.n304 dvss.n294 539.294
R2465 dvss.n299 dvss.n294 539.294
R2466 dvss.n299 dvss.n290 539.294
R2467 dvss.n3727 dvss.n290 539.294
R2468 dvss.n3727 dvss.n284 539.294
R2469 dvss.n3746 dvss.n284 539.294
R2470 dvss.n3747 dvss.n3746 539.294
R2471 dvss.n3747 dvss.n277 539.294
R2472 dvss.n278 dvss.n277 539.294
R2473 dvss.n3753 dvss.n278 539.294
R2474 dvss.n3753 dvss.n269 539.294
R2475 dvss.n269 dvss.n261 539.294
R2476 dvss.n3769 dvss.n261 539.294
R2477 dvss.n3819 dvss.n3769 539.294
R2478 dvss.n3774 dvss.n3773 539.294
R2479 dvss.n3824 dvss.n3823 539.294
R2480 dvss.n3824 dvss.n3783 539.294
R2481 dvss.n3784 dvss.n3783 539.294
R2482 dvss.n3831 dvss.n3784 539.294
R2483 dvss.n3832 dvss.n3831 539.294
R2484 dvss.n3832 dvss.n3794 539.294
R2485 dvss.n3795 dvss.n3794 539.294
R2486 dvss.n3801 dvss.n3795 539.294
R2487 dvss.n3801 dvss.n3800 539.294
R2488 dvss.n3800 dvss.n122 539.294
R2489 dvss.n128 dvss.n122 539.294
R2490 dvss.n198 dvss.n128 539.294
R2491 dvss.n200 dvss.n198 539.294
R2492 dvss.n200 dvss.n194 539.294
R2493 dvss.n209 dvss.n194 539.294
R2494 dvss.n209 dvss.n190 539.294
R2495 dvss.n190 dvss.n141 539.294
R2496 dvss.n142 dvss.n141 539.294
R2497 dvss.n181 dvss.n142 539.294
R2498 dvss.n148 dvss.n147 539.294
R2499 dvss.n186 dvss.n185 539.294
R2500 dvss.n186 dvss.n157 539.294
R2501 dvss.n158 dvss.n157 539.294
R2502 dvss.n176 dvss.n158 539.294
R2503 dvss.n177 dvss.n176 539.294
R2504 dvss.n177 dvss.n168 539.294
R2505 dvss.n169 dvss.n168 539.294
R2506 dvss.n4094 dvss.n169 539.294
R2507 dvss.n4096 dvss.n4094 539.294
R2508 dvss.n4096 dvss.n97 539.294
R2509 dvss.n4195 dvss.n97 539.294
R2510 dvss.n4196 dvss.n4195 539.294
R2511 dvss.n4196 dvss.n92 539.294
R2512 dvss.n92 dvss.n81 539.294
R2513 dvss.n4223 dvss.n81 539.294
R2514 dvss.n4224 dvss.n4223 539.294
R2515 dvss.n4224 dvss.n72 539.294
R2516 dvss.n72 dvss.n66 539.294
R2517 dvss.n4238 dvss.n66 539.294
R2518 dvss.n4239 dvss.n4238 539.294
R2519 dvss.n2572 dvss.n2113 539.294
R2520 dvss.n2115 dvss.n2113 539.294
R2521 dvss.n2116 dvss.n2115 539.294
R2522 dvss.n2210 dvss.n2116 539.294
R2523 dvss.n2210 dvss.n2120 539.294
R2524 dvss.n2121 dvss.n2120 539.294
R2525 dvss.n2214 dvss.n2121 539.294
R2526 dvss.n2214 dvss.n2126 539.294
R2527 dvss.n2127 dvss.n2126 539.294
R2528 dvss.n2218 dvss.n2127 539.294
R2529 dvss.n2218 dvss.n2130 539.294
R2530 dvss.n2131 dvss.n2130 539.294
R2531 dvss.n2229 dvss.n2131 539.294
R2532 dvss.n2229 dvss.n2228 539.294
R2533 dvss.n2228 dvss.n2137 539.294
R2534 dvss.n2138 dvss.n2137 539.294
R2535 dvss.n2223 dvss.n2138 539.294
R2536 dvss.n2223 dvss.n2140 539.294
R2537 dvss.n2141 dvss.n2140 539.294
R2538 dvss.n2143 dvss.n2141 539.294
R2539 dvss.n2522 dvss.n2143 539.294
R2540 dvss.n977 dvss.n879 533.678
R2541 dvss.n791 dvss.n790 533.678
R2542 dvss.n1103 dvss.n776 510.284
R2543 dvss.n2043 dvss.n2042 498.113
R2544 dvss.n2044 dvss.n2043 498.113
R2545 dvss.n2056 dvss.n2045 498.113
R2546 dvss.n2055 dvss.n2054 498.113
R2547 dvss.n2054 dvss.n2053 498.113
R2548 dvss.n2053 dvss.n2052 498.113
R2549 dvss.n2052 dvss.n2050 498.113
R2550 dvss.n3196 dvss.n2089 498.113
R2551 dvss.n3197 dvss.n3196 498.113
R2552 dvss.n3199 dvss.n3198 498.113
R2553 dvss.n3213 dvss.n3212 498.113
R2554 dvss.n3214 dvss.n3213 498.113
R2555 dvss.n3214 dvss.n2079 498.113
R2556 dvss.n3223 dvss.n2079 498.113
R2557 dvss.n3224 dvss.n3223 498.113
R2558 dvss.n2050 dvss.n2049 493.485
R2559 dvss.n4237 dvss.n57 491.163
R2560 dvss.n1017 dvss.n1016 486.048
R2561 dvss.n2521 dvss.n2520 479.541
R2562 dvss dvss.t592 446.038
R2563 dvss dvss.t554 446.038
R2564 dvss.n1015 dvss.n776 445.116
R2565 dvss.t570 dvss.n2044 441.038
R2566 dvss.t721 dvss.n3197 441.038
R2567 dvss.n4087 dvss.n175 432.788
R2568 dvss.n3833 dvss.n3830 432.788
R2569 dvss.n3701 dvss.n305 432.788
R2570 dvss.n3583 dvss.n3582 432.788
R2571 dvss.n3470 dvss.n431 432.788
R2572 dvss.n1671 dvss.n1640 432.788
R2573 dvss.n1519 dvss.n550 432.788
R2574 dvss.n1249 dvss.n1248 432.788
R2575 dvss.n1139 dvss.n762 432.788
R2576 dvss.n4079 dvss.t457 410.247
R2577 dvss.n3829 dvss.t35 410.247
R2578 dvss.n3698 dvss.t2 410.247
R2579 dvss.n3579 dvss.t237 410.247
R2580 dvss.n3457 dvss.t210 410.247
R2581 dvss.n1663 dvss.t331 410.247
R2582 dvss.n1506 dvss.t222 410.247
R2583 dvss.n1250 dvss.t234 410.247
R2584 dvss.n1126 dvss.t32 410.247
R2585 dvss.n2521 dvss.n2144 403.825
R2586 dvss.n2573 dvss.n2112 403.825
R2587 dvss.t463 dvss.n4088 401.229
R2588 dvss.t41 dvss.n3836 401.229
R2589 dvss.t8 dvss.n3720 401.229
R2590 dvss.t243 dvss.n3604 401.229
R2591 dvss.n432 dvss.t206 401.229
R2592 dvss.t333 dvss.n1672 401.229
R2593 dvss.n551 dvss.t216 401.229
R2594 dvss.n657 dvss.t228 401.229
R2595 dvss.n1140 dvss.t24 401.229
R2596 dvss.n4077 dvss.n179 396.721
R2597 dvss.n3825 dvss.n3817 396.721
R2598 dvss.n324 dvss.n323 396.721
R2599 dvss.n382 dvss.n381 396.721
R2600 dvss.n3443 dvss.n3442 396.721
R2601 dvss.n1661 dvss.n1644 396.721
R2602 dvss.n1492 dvss.n1491 396.721
R2603 dvss.n1257 dvss.n1256 396.721
R2604 dvss.n1117 dvss.n776 396.721
R2605 dvss.n2220 dvss.n2144 395.663
R2606 dvss.n2226 dvss.n2225 394.031
R2607 dvss.n2225 dvss.n2224 394.031
R2608 dvss.n2221 dvss.n2220 394.031
R2609 dvss.n3226 dvss.n3224 389.37
R2610 dvss.n3154 dvss.n3153 389.37
R2611 dvss.n800 dvss.n793 380.784
R2612 dvss.n2231 dvss.n2230 379.724
R2613 dvss.n2411 dvss.t75 379.31
R2614 dvss.n2042 dvss.n2040 368.271
R2615 dvss.n3187 dvss.n2089 368.271
R2616 dvss.n2208 dvss.n2112 366.872
R2617 dvss.n2209 dvss.n2208 363.512
R2618 dvss.n2213 dvss.n2212 363.512
R2619 dvss.n2217 dvss.n2216 363.512
R2620 dvss.n2232 dvss.n2231 363.512
R2621 dvss.n4237 dvss.n67 358.591
R2622 dvss.n853 dvss.t563 349.909
R2623 dvss.t117 dvss.n837 349.909
R2624 dvss.n4259 dvss.t311 348.875
R2625 dvss.n2211 dvss.t455 344.579
R2626 dvss.n3226 dvss.n3225 342.301
R2627 dvss.n2013 dvss.n2012 342.301
R2628 dvss.n2025 dvss.n2007 342.301
R2629 dvss.n2040 dvss.n2039 342.301
R2630 dvss.n3155 dvss.n3154 342.301
R2631 dvss.n3167 dvss.n3166 342.301
R2632 dvss.n3170 dvss.n3169 342.301
R2633 dvss.n3187 dvss.n3186 342.301
R2634 dvss.t451 dvss.n2215 337.005
R2635 dvss.n4199 dvss.n96 332.075
R2636 dvss.n4227 dvss.n67 332.075
R2637 dvss.n197 dvss.n196 332.075
R2638 dvss.n4068 dvss.n4067 332.075
R2639 dvss.n3748 dvss.n283 332.075
R2640 dvss.n3879 dvss.n262 332.075
R2641 dvss.n3635 dvss.n345 332.075
R2642 dvss.n3661 dvss.n3660 332.075
R2643 dvss.n3516 dvss.n414 332.075
R2644 dvss.n3543 dvss.n3542 332.075
R2645 dvss.n1686 dvss.n1685 332.075
R2646 dvss.n3441 dvss.n445 332.075
R2647 dvss.n1565 dvss.n533 332.075
R2648 dvss.n1748 dvss.n507 332.075
R2649 dvss.n692 dvss.n691 332.075
R2650 dvss.n1490 dvss.n564 332.075
R2651 dvss.n1178 dvss.n744 332.075
R2652 dvss.n1265 dvss.n627 332.075
R2653 dvss.t285 dvss.t536 331.955
R2654 dvss.t536 dvss.t574 331.955
R2655 dvss.t565 dvss.t193 327.353
R2656 dvss.t252 dvss.t123 317.724
R2657 dvss.t565 dvss.t137 317.724
R2658 dvss.n3237 dvss.t362 306.646
R2659 dvss.n2106 dvss.t604 306.646
R2660 dvss.n4088 dvss.t461 302.05
R2661 dvss.n3836 dvss.t39 302.05
R2662 dvss.n3720 dvss.t6 302.05
R2663 dvss.n3604 dvss.t241 302.05
R2664 dvss.t208 dvss.n432 302.05
R2665 dvss.n1672 dvss.t327 302.05
R2666 dvss.t218 dvss.n551 302.05
R2667 dvss.n657 dvss.t232 302.05
R2668 dvss.n1140 dvss.t30 302.05
R2669 dvss.n2056 dvss.t558 300.943
R2670 dvss.n3198 dvss.t55 300.943
R2671 dvss.n4188 dvss.t703 297.485
R2672 dvss.n4151 dvss.t374 297.485
R2673 dvss.n1997 dvss.t403 297.485
R2674 dvss.n3621 dvss.t344 297.485
R2675 dvss.n1945 dvss.t97 297.485
R2676 dvss.n1682 dvss.t425 297.485
R2677 dvss.n1388 dvss.t275 297.485
R2678 dvss.n688 dvss.t394 297.485
R2679 dvss.n1163 dvss.t133 297.485
R2680 dvss.n2224 dvss.n2222 295.522
R2681 dvss.n4079 dvss.t459 293.034
R2682 dvss.t37 dvss.n3829 293.034
R2683 dvss.n3698 dvss.t4 293.034
R2684 dvss.n3579 dvss.t239 293.034
R2685 dvss.n3457 dvss.t212 293.034
R2686 dvss.n1663 dvss.t329 293.034
R2687 dvss.n1506 dvss.t220 293.034
R2688 dvss.n1250 dvss.t230 293.034
R2689 dvss.n1126 dvss.t26 293.034
R2690 dvss.n2026 dvss.t364 292.384
R2691 dvss.t606 dvss.n3168 292.384
R2692 dvss.t294 dvss.t478 284.077
R2693 dvss.n4222 dvss.t705 283.649
R2694 dvss.n208 dvss.t384 283.649
R2695 dvss.n3754 dvss.t405 283.649
R2696 dvss.t346 dvss.n3639 283.649
R2697 dvss.n3523 dvss.t93 283.649
R2698 dvss.n1693 dvss.t429 283.649
R2699 dvss.n1571 dvss.t267 283.649
R2700 dvss.n699 dvss.t390 283.649
R2701 dvss.n1184 dvss.t129 283.649
R2702 dvss.n8 dvss.t545 283.474
R2703 dvss.n2344 dvss.t637 282.327
R2704 dvss.n2430 dvss.t154 282.327
R2705 dvss.n2511 dvss.t547 282.327
R2706 dvss.n4 dvss.t599 282.327
R2707 dvss.t516 dvss.t494 281.707
R2708 dvss.t494 dvss.t518 281.707
R2709 dvss.t518 dvss.t508 281.707
R2710 dvss.t508 dvss.t520 281.707
R2711 dvss.t520 dvss.t500 281.707
R2712 dvss.t500 dvss.t514 281.707
R2713 dvss.t514 dvss.t504 281.707
R2714 dvss.t504 dvss.t490 281.707
R2715 dvss.t490 dvss.t506 281.707
R2716 dvss.t506 dvss.t492 281.707
R2717 dvss.t492 dvss.t496 281.707
R2718 dvss.t496 dvss.t510 281.707
R2719 dvss.t498 dvss.t512 281.707
R2720 dvss.t512 dvss.t502 281.707
R2721 dvss.t592 dvss.t596 281.707
R2722 dvss.t596 dvss.t594 281.707
R2723 dvss.t594 dvss.t598 281.707
R2724 dvss.t554 dvss.t548 281.707
R2725 dvss.t548 dvss.t540 281.707
R2726 dvss.t540 dvss.t544 281.707
R2727 dvss.n2341 dvss.t633 281.13
R2728 dvss.n2423 dvss.t160 281.13
R2729 dvss.n2504 dvss.t557 281.13
R2730 dvss.n4405 dvss.t593 281.13
R2731 dvss.n5 dvss.t555 281.13
R2732 dvss.n4068 dvss.n179 276.731
R2733 dvss.n3817 dvss.n262 276.731
R2734 dvss.n3661 dvss.n324 276.731
R2735 dvss.n3543 dvss.n382 276.731
R2736 dvss.n3442 dvss.n3441 276.731
R2737 dvss.n1644 dvss.n507 276.731
R2738 dvss.n1491 dvss.n1490 276.731
R2739 dvss.n1257 dvss.n627 276.731
R2740 dvss.n2049 dvss.n2048 275.899
R2741 dvss.n2048 dvss.n2046 275.899
R2742 dvss.n121 dvss.n104 275.899
R2743 dvss.n4159 dvss.n4158 275.899
R2744 dvss.n4160 dvss.n4159 275.899
R2745 dvss.n4162 dvss.n4160 275.899
R2746 dvss.n4163 dvss.n4162 275.899
R2747 dvss.n4164 dvss.n4163 275.899
R2748 dvss.n4168 dvss.n4165 275.899
R2749 dvss.n4170 dvss.n4169 275.899
R2750 dvss.n4172 dvss.n4170 275.899
R2751 dvss.n4173 dvss.n4172 275.899
R2752 dvss.n4174 dvss.n4173 275.899
R2753 dvss.n4176 dvss.n4174 275.899
R2754 dvss.n4177 dvss.n4176 275.899
R2755 dvss.n4178 dvss.n4177 275.899
R2756 dvss.n4186 dvss.n4185 275.899
R2757 dvss.n79 dvss.n77 275.899
R2758 dvss.n77 dvss.n76 275.899
R2759 dvss.n76 dvss.n56 275.899
R2760 dvss.n4312 dvss.n56 275.899
R2761 dvss.t510 dvss.n2486 271.647
R2762 dvss.n2370 dvss.n2368 270.307
R2763 dvss.n2439 dvss.n2368 270.307
R2764 dvss.n2438 dvss.n2370 270.307
R2765 dvss.n2439 dvss.n2438 270.307
R2766 dvss.t372 dvss.n2026 263.858
R2767 dvss.n3168 dvss.t612 263.858
R2768 dvss.t502 dvss 261.586
R2769 dvss.t763 dvss.n4077 261.476
R2770 dvss.t12 dvss.n3825 261.476
R2771 dvss.n323 dvss.t247 261.476
R2772 dvss.n381 dvss.t224 261.476
R2773 dvss.n3443 dvss.t398 261.476
R2774 dvss.t709 dvss.n1661 261.476
R2775 dvss.n1492 dvss.t723 261.476
R2776 dvss.n1256 dvss.t113 261.476
R2777 dvss.n1117 dvss.t195 261.476
R2778 dvss.n2027 dvss.n259 256.726
R2779 dvss.n3185 dvss.n3184 256.726
R2780 dvss.n4222 dvss.t701 255.976
R2781 dvss.n208 dvss.t380 255.976
R2782 dvss.n3754 dvss.t413 255.976
R2783 dvss.n3639 dvss.t352 255.976
R2784 dvss.n3523 dvss.t89 255.976
R2785 dvss.n1693 dvss.t427 255.976
R2786 dvss.n1571 dvss.t269 255.976
R2787 dvss.n699 dvss.t388 255.976
R2788 dvss.n1184 dvss.t127 255.976
R2789 dvss.n1011 dvss.n839 255.845
R2790 dvss.n1005 dvss.n839 255.845
R2791 dvss.n1005 dvss.n1004 255.845
R2792 dvss.n1004 dvss.n1003 255.845
R2793 dvss.n1003 dvss.n845 255.845
R2794 dvss.n997 dvss.n845 255.845
R2795 dvss.n997 dvss.n996 255.845
R2796 dvss.n988 dvss.n864 255.845
R2797 dvss.n988 dvss.n987 255.845
R2798 dvss.n980 dvss.n877 255.845
R2799 dvss.n980 dvss.n979 255.845
R2800 dvss.n972 dvss.n878 255.845
R2801 dvss.n2215 dvss.t449 253.702
R2802 dvss.n978 dvss.n878 253.18
R2803 dvss.n972 dvss.n971 252.209
R2804 dvss.t534 dvss.t282 252.159
R2805 dvss.t282 dvss.t111 252.159
R2806 dvss.t111 dvss.t285 252.159
R2807 dvss.n3979 dvss.n3978 251.879
R2808 dvss.n3984 dvss.n3983 251.879
R2809 dvss.n3987 dvss.n3986 251.879
R2810 dvss.n4002 dvss.n4001 251.879
R2811 dvss.n4003 dvss.n4002 251.879
R2812 dvss.n4004 dvss.n4003 251.879
R2813 dvss.n4009 dvss.n4008 251.879
R2814 dvss.n4010 dvss.n4009 251.879
R2815 dvss.n4309 dvss.n59 251.879
R2816 dvss.n3905 dvss.n3904 251.879
R2817 dvss.n3919 dvss.n241 251.879
R2818 dvss.n3922 dvss.n3921 251.879
R2819 dvss.n3935 dvss.n3934 251.879
R2820 dvss.n3937 dvss.n3935 251.879
R2821 dvss.n3937 dvss.n3936 251.879
R2822 dvss.n3951 dvss.n3950 251.879
R2823 dvss.n3951 dvss.n216 251.879
R2824 dvss.n4064 dvss.n217 251.879
R2825 dvss.n1991 dvss.n1990 251.879
R2826 dvss.n1995 dvss.n1994 251.879
R2827 dvss.n3240 dvss.n3239 251.879
R2828 dvss.n3243 dvss.n3242 251.879
R2829 dvss.n3244 dvss.n3243 251.879
R2830 dvss.n3245 dvss.n3244 251.879
R2831 dvss.n3250 dvss.n3249 251.879
R2832 dvss.n3250 dvss.n258 251.879
R2833 dvss.n3883 dvss.n3882 251.879
R2834 dvss.n1966 dvss.n1965 251.879
R2835 dvss.n1970 dvss.n1969 251.879
R2836 dvss.n1973 dvss.n1972 251.879
R2837 dvss.n1976 dvss.n1975 251.879
R2838 dvss.n1977 dvss.n1976 251.879
R2839 dvss.n1978 dvss.n1977 251.879
R2840 dvss.n1983 dvss.n1982 251.879
R2841 dvss.n1985 dvss.n1983 251.879
R2842 dvss.n1988 dvss.n1987 251.879
R2843 dvss.n1938 dvss.n1937 251.879
R2844 dvss.n1943 dvss.n1942 251.879
R2845 dvss.n1948 dvss.n1947 251.879
R2846 dvss.n1951 dvss.n1950 251.879
R2847 dvss.n1952 dvss.n1951 251.879
R2848 dvss.n1953 dvss.n1952 251.879
R2849 dvss.n1958 dvss.n1957 251.879
R2850 dvss.n1960 dvss.n1958 251.879
R2851 dvss.n1963 dvss.n1962 251.879
R2852 dvss.n1774 dvss.n1773 251.879
R2853 dvss.n1788 dvss.n487 251.879
R2854 dvss.n1791 dvss.n1790 251.879
R2855 dvss.n1804 dvss.n1803 251.879
R2856 dvss.n1806 dvss.n1804 251.879
R2857 dvss.n1806 dvss.n1805 251.879
R2858 dvss.n1820 dvss.n1819 251.879
R2859 dvss.n1820 dvss.n462 251.879
R2860 dvss.n3407 dvss.n463 251.879
R2861 dvss.n1381 dvss.n1380 251.879
R2862 dvss.n1386 dvss.n1385 251.879
R2863 dvss.n1391 dvss.n1390 251.879
R2864 dvss.n1394 dvss.n1393 251.879
R2865 dvss.n1395 dvss.n1394 251.879
R2866 dvss.n1396 dvss.n1395 251.879
R2867 dvss.n1401 dvss.n1400 251.879
R2868 dvss.n1401 dvss.n504 251.879
R2869 dvss.n1752 dvss.n1751 251.879
R2870 dvss.n1291 dvss.n1290 251.879
R2871 dvss.n1305 dvss.n607 251.879
R2872 dvss.n1308 dvss.n1307 251.879
R2873 dvss.n1321 dvss.n1320 251.879
R2874 dvss.n1323 dvss.n1321 251.879
R2875 dvss.n1323 dvss.n1322 251.879
R2876 dvss.n1337 dvss.n1336 251.879
R2877 dvss.n1337 dvss.n582 251.879
R2878 dvss.n1458 dvss.n583 251.879
R2879 dvss.n971 dvss.n970 251.879
R2880 dvss.n964 dvss.n963 251.879
R2881 dvss.n956 dvss.n955 251.879
R2882 dvss.n953 dvss.n952 251.879
R2883 dvss.n952 dvss.n951 251.879
R2884 dvss.n951 dvss.n904 251.879
R2885 dvss.n944 dvss.n943 251.879
R2886 dvss.n943 dvss.n624 251.879
R2887 dvss.n1269 dvss.n1268 251.879
R2888 dvss.t598 dvss 251.524
R2889 dvss.t544 dvss 251.524
R2890 dvss.n4226 dvss.n4225 249.058
R2891 dvss.n4066 dvss.n215 249.058
R2892 dvss.n3880 dvss.n260 249.058
R2893 dvss.n3638 dvss.n327 249.058
R2894 dvss.n3522 dvss.n389 249.058
R2895 dvss.n3410 dvss.n3409 249.058
R2896 dvss.n1749 dvss.n505 249.058
R2897 dvss.n1461 dvss.n1460 249.058
R2898 dvss.n1266 dvss.n625 249.058
R2899 dvss.n986 dvss.t265 247.851
R2900 dvss.t178 dvss.n106 247.16
R2901 dvss.t621 dvss.n4184 247.16
R2902 dvss.t447 dvss.n2211 246.127
R2903 dvss.n1062 dvss.t567 245.276
R2904 dvss.n2670 dvss.t120 245.276
R2905 dvss.t53 dvss.n4164 244.286
R2906 dvss.t757 dvss.n2364 243.903
R2907 dvss.n2230 dvss.t524 242.165
R2908 dvss.n2492 dvss.t663 240.701
R2909 dvss.n864 dvss.t725 239.856
R2910 dvss.t561 dvss.n978 237.19
R2911 dvss.n4254 dvss.t281 236.975
R2912 dvss.n4256 dvss.t284 236.975
R2913 dvss.n2374 dvss.t296 236.149
R2914 dvss.n3978 dvss.n3977 230.888
R2915 dvss.n3904 dvss.n249 230.888
R2916 dvss.n1990 dvss.n1989 230.888
R2917 dvss.n1965 dvss.n1964 230.888
R2918 dvss.n1937 dvss.n1936 230.888
R2919 dvss.n1773 dvss.n495 230.888
R2920 dvss.n1380 dvss.n1379 230.888
R2921 dvss.n1290 dvss.n615 230.888
R2922 dvss.n1292 dvss.t715 226.6
R2923 dvss.n3982 dvss.t689 226.6
R2924 dvss.n3906 dvss.t141 226.6
R2925 dvss.n1993 dvss.t467 226.6
R2926 dvss.n1968 dvss.t14 226.6
R2927 dvss.n1941 dvss.t486 226.6
R2928 dvss.n1775 dvss.t441 226.6
R2929 dvss.n1384 dvss.t107 226.6
R2930 dvss.n897 dvss.t645 226.6
R2931 dvss.n4246 dvss.t293 223.559
R2932 dvss.n2233 dvss.n2232 223.409
R2933 dvss.t685 dvss.n3985 221.619
R2934 dvss.t147 dvss.n3920 221.619
R2935 dvss.t473 dvss.n1996 221.619
R2936 dvss.t20 dvss.n1971 221.619
R2937 dvss.t482 dvss.n1944 221.619
R2938 dvss.t443 dvss.n1789 221.619
R2939 dvss.t101 dvss.n1387 221.619
R2940 dvss.t719 dvss.n1306 221.619
R2941 dvss.n962 dvss.t647 221.619
R2942 dvss.n4182 dvss.n4181 220.345
R2943 dvss.t477 dvss.t294 218.643
R2944 dvss.n684 dvss.n656 217.097
R2945 dvss.n4089 dvss.n173 217.097
R2946 dvss.n3838 dvss.n3837 217.097
R2947 dvss.n3722 dvss.n3721 217.097
R2948 dvss.n3606 dvss.n3605 217.097
R2949 dvss.n3490 dvss.n3489 217.097
R2950 dvss.n1673 dvss.n1638 217.097
R2951 dvss.n1539 dvss.n1538 217.097
R2952 dvss.n1144 dvss.n759 217.097
R2953 dvss.n1052 dvss.n776 212.969
R2954 dvss.n1091 dvss.n776 212.969
R2955 dvss.n3238 dvss.n3237 210.374
R2956 dvss.n2106 dvss.n351 210.374
R2957 dvss.n4310 dvss.n4309 209.899
R2958 dvss.n3977 dvss.n217 209.899
R2959 dvss.n3882 dvss.n249 209.899
R2960 dvss.n1989 dvss.n1988 209.899
R2961 dvss.n1964 dvss.n1963 209.899
R2962 dvss.n1936 dvss.n463 209.899
R2963 dvss.n1751 dvss.n495 209.899
R2964 dvss.n1379 dvss.n583 209.899
R2965 dvss.n1268 dvss.n615 209.899
R2966 dvss.n4394 dvss.n7 207.213
R2967 dvss.n4403 dvss.n2 207.213
R2968 dvss.n2348 dvss.n2343 207.213
R2969 dvss.n2318 dvss.n2317 207.213
R2970 dvss.n2322 dvss.n2316 207.213
R2971 dvss.n2325 dvss.n2324 207.213
R2972 dvss.n2331 dvss.n2313 207.213
R2973 dvss.n2334 dvss.n2333 207.213
R2974 dvss.n2311 dvss.n2310 207.213
R2975 dvss.n2358 dvss.n2339 207.213
R2976 dvss.n2428 dvss.n2377 207.213
R2977 dvss.n2392 dvss.n2391 207.213
R2978 dvss.n2394 dvss.n2393 207.213
R2979 dvss.n2400 dvss.n2388 207.213
R2980 dvss.n2403 dvss.n2402 207.213
R2981 dvss.n2409 dvss.n2385 207.213
R2982 dvss.n2383 dvss.n2382 207.213
R2983 dvss.n2417 dvss.n2381 207.213
R2984 dvss.n2509 dvss.n2274 207.213
R2985 dvss.n2289 dvss.n2288 207.213
R2986 dvss.n2291 dvss.n2290 207.213
R2987 dvss.n2297 dvss.n2285 207.213
R2988 dvss.n2300 dvss.n2299 207.213
R2989 dvss.n2306 dvss.n2282 207.213
R2990 dvss.n2280 dvss.n2279 207.213
R2991 dvss.n2498 dvss.n2278 207.213
R2992 dvss.n2456 dvss.n2455 207.213
R2993 dvss.n2458 dvss.n2457 207.213
R2994 dvss.n2464 dvss.n2452 207.213
R2995 dvss.n2467 dvss.n2466 207.213
R2996 dvss.n2473 dvss.n2449 207.213
R2997 dvss.n2476 dvss.n2475 207.213
R2998 dvss.n2484 dvss.n2445 207.213
R2999 dvss.n4154 dvss.n4153 204.279
R3000 dvss.n4188 dvss.n4187 204.089
R3001 dvss.n4152 dvss.n4151 204.089
R3002 dvss.n3238 dvss.n1997 204.089
R3003 dvss.n3621 dvss.n351 204.089
R3004 dvss.n1946 dvss.n1945 204.089
R3005 dvss.n1682 dvss.n1681 204.089
R3006 dvss.n1389 dvss.n1388 204.089
R3007 dvss.n688 dvss.n687 204.089
R3008 dvss.n1163 dvss.n1162 204.089
R3009 dvss.t579 dvss.t312 202.685
R3010 dvss.t182 dvss.n106 201.177
R3011 dvss.n4184 dvss.t617 201.177
R3012 dvss.n2227 dvss.t552 201.119
R3013 dvss.t453 dvss.n2217 200.689
R3014 dvss.n2181 dvss.n2180 200.215
R3015 dvss.n1479 dvss.n563 200.215
R3016 dvss.n1656 dvss.n1655 200.215
R3017 dvss.n1657 dvss.n1656 200.215
R3018 dvss.n3427 dvss.n444 200.215
R3019 dvss.n3430 dvss.n444 200.215
R3020 dvss.n3562 dvss.n3561 200.215
R3021 dvss.n3563 dvss.n3562 200.215
R3022 dvss.n3665 dvss.n3664 200.215
R3023 dvss.n3666 dvss.n3665 200.215
R3024 dvss.n3816 dvss.n3815 200.215
R3025 dvss.n3816 dvss.n3811 200.215
R3026 dvss.n4072 dvss.n4071 200.215
R3027 dvss.n4073 dvss.n4072 200.215
R3028 dvss.n1259 dvss.n1258 200.215
R3029 dvss.n1258 dvss.n636 200.215
R3030 dvss.n1378 dvss.n1377 200.215
R3031 dvss.n1378 dvss.n1376 200.215
R3032 dvss.n1762 dvss.n1761 200.215
R3033 dvss.n1763 dvss.n1762 200.215
R3034 dvss.n1935 dvss.n1934 200.215
R3035 dvss.n1935 dvss.n1933 200.215
R3036 dvss.n1930 dvss.n1929 200.215
R3037 dvss.n1930 dvss.n1927 200.215
R3038 dvss.n1924 dvss.n1923 200.215
R3039 dvss.n1924 dvss.n1921 200.215
R3040 dvss.n3893 dvss.n3892 200.215
R3041 dvss.n3894 dvss.n3893 200.215
R3042 dvss.n3976 dvss.n3975 200.215
R3043 dvss.n3976 dvss.n3974 200.215
R3044 dvss.n1279 dvss.n1278 200.215
R3045 dvss.n1280 dvss.n1279 200.215
R3046 dvss.n1204 dvss.n728 200.215
R3047 dvss.n728 dvss.n727 200.215
R3048 dvss.n1475 dvss.n1474 200.215
R3049 dvss.n1474 dvss.n1473 200.215
R3050 dvss.n1648 dvss.n1647 200.215
R3051 dvss.n1649 dvss.n1648 200.215
R3052 dvss.n3423 dvss.n3422 200.215
R3053 dvss.n3422 dvss.n3421 200.215
R3054 dvss.n3550 dvss.n3549 200.215
R3055 dvss.n3551 dvss.n3550 200.215
R3056 dvss.n3675 dvss.n3674 200.215
R3057 dvss.n3676 dvss.n3675 200.215
R3058 dvss.n3821 dvss.n3820 200.215
R3059 dvss.n3822 dvss.n3821 200.215
R3060 dvss.n183 dvss.n182 200.215
R3061 dvss.n184 dvss.n183 200.215
R3062 dvss.n1094 dvss.n793 200.215
R3063 dvss.n793 dvss.n792 200.215
R3064 dvss.n1103 dvss.n1102 200.215
R3065 dvss.n1104 dvss.n1103 200.215
R3066 dvss.n1091 dvss.n1090 200.215
R3067 dvss.n1091 dvss.n796 200.215
R3068 dvss.n1091 dvss.n797 200.215
R3069 dvss.n1091 dvss.n798 200.215
R3070 dvss.n1091 dvss.n799 200.215
R3071 dvss.n1052 dvss.n1051 200.215
R3072 dvss.n1052 dvss.n828 200.215
R3073 dvss.n1052 dvss.n829 200.215
R3074 dvss.n1052 dvss.n830 200.215
R3075 dvss.n1053 dvss.n1052 200.215
R3076 dvss.n3143 dvss.n3142 200.215
R3077 dvss.n3143 dvss.n2580 200.215
R3078 dvss.n3143 dvss.n2581 200.215
R3079 dvss.n3143 dvss.n2582 200.215
R3080 dvss.n3143 dvss.n2583 200.215
R3081 dvss.n3143 dvss.n2584 200.215
R3082 dvss.n3143 dvss.n2585 200.215
R3083 dvss.n3143 dvss.n2586 200.215
R3084 dvss.n3143 dvss.n2587 200.215
R3085 dvss.n3143 dvss.n2588 200.215
R3086 dvss.n3143 dvss.n2589 200.215
R3087 dvss.n3143 dvss.n2590 200.215
R3088 dvss.n3143 dvss.n2591 200.215
R3089 dvss.n3143 dvss.n2592 200.215
R3090 dvss.n3143 dvss.n2593 200.215
R3091 dvss.n3143 dvss.n2594 200.215
R3092 dvss.n3143 dvss.n2595 200.215
R3093 dvss.n3143 dvss.n2596 200.215
R3094 dvss.n3143 dvss.n2597 200.215
R3095 dvss.n3143 dvss.n2598 200.215
R3096 dvss.n3143 dvss.n2599 200.215
R3097 dvss.n3143 dvss.n2600 200.215
R3098 dvss.n3143 dvss.n2601 200.215
R3099 dvss.n3143 dvss.n2602 200.215
R3100 dvss.n3143 dvss.n2603 200.215
R3101 dvss.n3143 dvss.n2604 200.215
R3102 dvss.n3143 dvss.n2605 200.215
R3103 dvss.n3143 dvss.n2606 200.215
R3104 dvss.n3143 dvss.n2607 200.215
R3105 dvss.n3143 dvss.n2608 200.215
R3106 dvss.n3143 dvss.n2609 200.215
R3107 dvss.n3143 dvss.n2610 200.215
R3108 dvss.n3143 dvss.n2611 200.215
R3109 dvss.n3143 dvss.n2612 200.215
R3110 dvss.n3143 dvss.n2613 200.215
R3111 dvss.n3143 dvss.n2614 200.215
R3112 dvss.n3143 dvss.n2615 200.215
R3113 dvss.n3143 dvss.n2616 200.215
R3114 dvss.n3143 dvss.n2617 200.215
R3115 dvss.n3143 dvss.n2618 200.215
R3116 dvss.n3143 dvss.n2619 200.215
R3117 dvss.n3143 dvss.n2620 200.215
R3118 dvss.n3143 dvss.n2621 200.215
R3119 dvss.n3143 dvss.n2622 200.215
R3120 dvss.n3143 dvss.n2623 200.215
R3121 dvss.n3143 dvss.n2624 200.215
R3122 dvss.n3143 dvss.n2625 200.215
R3123 dvss.n3143 dvss.n2626 200.215
R3124 dvss.n3143 dvss.n2627 200.215
R3125 dvss.n3143 dvss.n2628 200.215
R3126 dvss.n3143 dvss.n2629 200.215
R3127 dvss.n3143 dvss.n2630 200.215
R3128 dvss.n3143 dvss.n2631 200.215
R3129 dvss.n3143 dvss.n2632 200.215
R3130 dvss.n3143 dvss.n2633 200.215
R3131 dvss.n3143 dvss.n2634 200.215
R3132 dvss.n3143 dvss.n2635 200.215
R3133 dvss.n3143 dvss.n2636 200.215
R3134 dvss.n3143 dvss.n2637 200.215
R3135 dvss.n3143 dvss.n2638 200.215
R3136 dvss.n3143 dvss.n2639 200.215
R3137 dvss.n3143 dvss.n2640 200.215
R3138 dvss.n3143 dvss.n2641 200.215
R3139 dvss.n3143 dvss.n2642 200.215
R3140 dvss.n3143 dvss.n2643 200.215
R3141 dvss.n3143 dvss.n2644 200.215
R3142 dvss.n3144 dvss.n3143 200.215
R3143 dvss.t558 dvss.n2055 197.171
R3144 dvss.n3212 dvss.t55 197.171
R3145 dvss.n4266 dvss.t579 194.704
R3146 dvss.t552 dvss.n2226 192.911
R3147 dvss.n4010 dvss.n80 188.91
R3148 dvss.n4065 dvss.n216 188.91
R3149 dvss.n3881 dvss.n258 188.91
R3150 dvss.n1986 dvss.n1985 188.91
R3151 dvss.n1961 dvss.n1960 188.91
R3152 dvss.n3408 dvss.n462 188.91
R3153 dvss.n1750 dvss.n504 188.91
R3154 dvss.n1459 dvss.n582 188.91
R3155 dvss.n1267 dvss.n624 188.91
R3156 dvss.t623 dvss.n4180 188.212
R3157 dvss.n4155 dvss.t188 188.212
R3158 dvss.n396 dvss.t771 186.374
R3159 dvss.n454 dvss.t770 186.374
R3160 dvss.n574 dvss.t775 186.374
R3161 dvss.n515 dvss.t774 186.374
R3162 dvss.n3353 dvss.t773 186.374
R3163 dvss.n1824 dvss.t772 186.374
R3164 dvss.n1404 dvss.t776 186.374
R3165 dvss.n1341 dvss.t777 186.374
R3166 dvss.n1061 dvss.n1060 185
R3167 dvss.n2669 dvss.n2668 185
R3168 dvss.n2182 dvss.n2181 184.572
R3169 dvss.n3137 dvss.n2580 184.572
R3170 dvss.n3134 dvss.n2581 184.572
R3171 dvss.n3130 dvss.n2582 184.572
R3172 dvss.n3126 dvss.n2583 184.572
R3173 dvss.n3122 dvss.n2584 184.572
R3174 dvss.n3118 dvss.n2585 184.572
R3175 dvss.n3114 dvss.n2586 184.572
R3176 dvss.n3110 dvss.n2587 184.572
R3177 dvss.n3106 dvss.n2588 184.572
R3178 dvss.n3102 dvss.n2589 184.572
R3179 dvss.n3098 dvss.n2590 184.572
R3180 dvss.n3094 dvss.n2591 184.572
R3181 dvss.n3090 dvss.n2592 184.572
R3182 dvss.n3086 dvss.n2593 184.572
R3183 dvss.n3082 dvss.n2594 184.572
R3184 dvss.n3078 dvss.n2595 184.572
R3185 dvss.n3074 dvss.n2596 184.572
R3186 dvss.n3070 dvss.n2597 184.572
R3187 dvss.n3066 dvss.n2598 184.572
R3188 dvss.n3062 dvss.n2599 184.572
R3189 dvss.n3058 dvss.n2600 184.572
R3190 dvss.n3054 dvss.n2601 184.572
R3191 dvss.n3050 dvss.n2602 184.572
R3192 dvss.n3046 dvss.n2603 184.572
R3193 dvss.n3042 dvss.n2604 184.572
R3194 dvss.n3038 dvss.n2605 184.572
R3195 dvss.n3034 dvss.n2606 184.572
R3196 dvss.n3030 dvss.n2607 184.572
R3197 dvss.n3026 dvss.n2608 184.572
R3198 dvss.n3022 dvss.n2609 184.572
R3199 dvss.n3018 dvss.n2610 184.572
R3200 dvss.n3014 dvss.n2611 184.572
R3201 dvss.n3010 dvss.n2612 184.572
R3202 dvss.n3006 dvss.n2613 184.572
R3203 dvss.n3002 dvss.n2614 184.572
R3204 dvss.n2998 dvss.n2615 184.572
R3205 dvss.n2994 dvss.n2616 184.572
R3206 dvss.n2990 dvss.n2617 184.572
R3207 dvss.n2986 dvss.n2618 184.572
R3208 dvss.n2982 dvss.n2619 184.572
R3209 dvss.n2978 dvss.n2620 184.572
R3210 dvss.n2974 dvss.n2621 184.572
R3211 dvss.n2970 dvss.n2622 184.572
R3212 dvss.n2966 dvss.n2623 184.572
R3213 dvss.n2962 dvss.n2624 184.572
R3214 dvss.n2958 dvss.n2625 184.572
R3215 dvss.n2954 dvss.n2626 184.572
R3216 dvss.n2950 dvss.n2627 184.572
R3217 dvss.n2946 dvss.n2628 184.572
R3218 dvss.n2942 dvss.n2629 184.572
R3219 dvss.n2938 dvss.n2630 184.572
R3220 dvss.n2934 dvss.n2631 184.572
R3221 dvss.n2930 dvss.n2632 184.572
R3222 dvss.n2926 dvss.n2633 184.572
R3223 dvss.n2922 dvss.n2634 184.572
R3224 dvss.n2918 dvss.n2635 184.572
R3225 dvss.n2914 dvss.n2636 184.572
R3226 dvss.n2910 dvss.n2637 184.572
R3227 dvss.n2906 dvss.n2638 184.572
R3228 dvss.n2902 dvss.n2639 184.572
R3229 dvss.n2898 dvss.n2640 184.572
R3230 dvss.n2894 dvss.n2641 184.572
R3231 dvss.n2890 dvss.n2642 184.572
R3232 dvss.n2886 dvss.n2643 184.572
R3233 dvss.n2882 dvss.n2644 184.572
R3234 dvss.n3145 dvss.n3144 184.572
R3235 dvss.n1051 dvss.n1050 184.572
R3236 dvss.n1045 dvss.n828 184.572
R3237 dvss.n1042 dvss.n829 184.572
R3238 dvss.n1038 dvss.n830 184.572
R3239 dvss.n1053 dvss.n827 184.572
R3240 dvss.n1102 dvss.n1101 184.572
R3241 dvss.n1105 dvss.n1104 184.572
R3242 dvss.n1260 dvss.n1259 184.572
R3243 dvss.n639 dvss.n636 184.572
R3244 dvss.n1479 dvss.n1478 184.572
R3245 dvss.n1655 dvss.n1654 184.572
R3246 dvss.n1658 dvss.n1657 184.572
R3247 dvss.n3427 dvss.n448 184.572
R3248 dvss.n3430 dvss.n3429 184.572
R3249 dvss.n3561 dvss.n3560 184.572
R3250 dvss.n3564 dvss.n3563 184.572
R3251 dvss.n3664 dvss.n3663 184.572
R3252 dvss.n3666 dvss.n322 184.572
R3253 dvss.n3815 dvss.n3814 184.572
R3254 dvss.n3811 dvss.n3810 184.572
R3255 dvss.n4071 dvss.n4070 184.572
R3256 dvss.n4074 dvss.n4073 184.572
R3257 dvss.n1480 dvss.n1479 184.572
R3258 dvss.n1655 dvss.n1653 184.572
R3259 dvss.n1657 dvss.n1652 184.572
R3260 dvss.n3428 dvss.n3427 184.572
R3261 dvss.n3431 dvss.n3430 184.572
R3262 dvss.n3561 dvss.n383 184.572
R3263 dvss.n3563 dvss.n380 184.572
R3264 dvss.n3664 dvss.n321 184.572
R3265 dvss.n3667 dvss.n3666 184.572
R3266 dvss.n3815 dvss.n3813 184.572
R3267 dvss.n3812 dvss.n3811 184.572
R3268 dvss.n4071 dvss.n188 184.572
R3269 dvss.n4073 dvss.n187 184.572
R3270 dvss.n1259 dvss.n635 184.572
R3271 dvss.n1208 dvss.n636 184.572
R3272 dvss.n1278 dvss.n1277 184.572
R3273 dvss.n1281 dvss.n1280 184.572
R3274 dvss.n1377 dvss.n1347 184.572
R3275 dvss.n1376 dvss.n1375 184.572
R3276 dvss.n1761 dvss.n1760 184.572
R3277 dvss.n1764 dvss.n1763 184.572
R3278 dvss.n1934 dvss.n1830 184.572
R3279 dvss.n1933 dvss.n1932 184.572
R3280 dvss.n1929 dvss.n1928 184.572
R3281 dvss.n1927 dvss.n1863 184.572
R3282 dvss.n1923 dvss.n1922 184.572
R3283 dvss.n1921 dvss.n1894 184.572
R3284 dvss.n3892 dvss.n3891 184.572
R3285 dvss.n3895 dvss.n3894 184.572
R3286 dvss.n3975 dvss.n3956 184.572
R3287 dvss.n3974 dvss.n3973 184.572
R3288 dvss.n61 dvss.n58 184.572
R3289 dvss.n1377 dvss.n1348 184.572
R3290 dvss.n1376 dvss.n1350 184.572
R3291 dvss.n1761 dvss.n499 184.572
R3292 dvss.n1763 dvss.n496 184.572
R3293 dvss.n1934 dvss.n1831 184.572
R3294 dvss.n1933 dvss.n1833 184.572
R3295 dvss.n1929 dvss.n1862 184.572
R3296 dvss.n1927 dvss.n1926 184.572
R3297 dvss.n1923 dvss.n1893 184.572
R3298 dvss.n1921 dvss.n1920 184.572
R3299 dvss.n3892 dvss.n253 184.572
R3300 dvss.n3894 dvss.n250 184.572
R3301 dvss.n3975 dvss.n3957 184.572
R3302 dvss.n3974 dvss.n3959 184.572
R3303 dvss.n1278 dvss.n619 184.572
R3304 dvss.n1280 dvss.n616 184.572
R3305 dvss.n1090 dvss.n1089 184.572
R3306 dvss.n1084 dvss.n796 184.572
R3307 dvss.n1081 dvss.n797 184.572
R3308 dvss.n1077 dvss.n798 184.572
R3309 dvss.n1073 dvss.n799 184.572
R3310 dvss.n1094 dvss.n1093 184.572
R3311 dvss.n792 dvss.n791 184.572
R3312 dvss.n1204 dvss.n1203 184.572
R3313 dvss.n727 dvss.n724 184.572
R3314 dvss.n1475 dvss.n1471 184.572
R3315 dvss.n1473 dvss.n561 184.572
R3316 dvss.n1647 dvss.n1646 184.572
R3317 dvss.n1650 dvss.n1649 184.572
R3318 dvss.n3423 dvss.n3419 184.572
R3319 dvss.n3421 dvss.n442 184.572
R3320 dvss.n3549 dvss.n3545 184.572
R3321 dvss.n3551 dvss.n3547 184.572
R3322 dvss.n3674 dvss.n3673 184.572
R3323 dvss.n3677 dvss.n3676 184.572
R3324 dvss.n3820 dvss.n3819 184.572
R3325 dvss.n3823 dvss.n3822 184.572
R3326 dvss.n182 dvss.n181 184.572
R3327 dvss.n185 dvss.n184 184.572
R3328 dvss.n1205 dvss.n1204 184.572
R3329 dvss.n727 dvss.n726 184.572
R3330 dvss.n1476 dvss.n1475 184.572
R3331 dvss.n1473 dvss.n1472 184.572
R3332 dvss.n1647 dvss.n1590 184.572
R3333 dvss.n1649 dvss.n1591 184.572
R3334 dvss.n3424 dvss.n3423 184.572
R3335 dvss.n3421 dvss.n3420 184.572
R3336 dvss.n3549 dvss.n3546 184.572
R3337 dvss.n3552 dvss.n3551 184.572
R3338 dvss.n3674 dvss.n315 184.572
R3339 dvss.n3676 dvss.n313 184.572
R3340 dvss.n3820 dvss.n3773 184.572
R3341 dvss.n3822 dvss.n3774 184.572
R3342 dvss.n182 dvss.n147 184.572
R3343 dvss.n184 dvss.n148 184.572
R3344 dvss.n1095 dvss.n1094 184.572
R3345 dvss.n792 dvss.n778 184.572
R3346 dvss.n1102 dvss.n782 184.572
R3347 dvss.n1104 dvss.n775 184.572
R3348 dvss.n1090 dvss.n802 184.572
R3349 dvss.n1082 dvss.n796 184.572
R3350 dvss.n1078 dvss.n797 184.572
R3351 dvss.n1074 dvss.n798 184.572
R3352 dvss.n799 dvss.n794 184.572
R3353 dvss.n1051 dvss.n832 184.572
R3354 dvss.n1043 dvss.n828 184.572
R3355 dvss.n1039 dvss.n829 184.572
R3356 dvss.n1035 dvss.n830 184.572
R3357 dvss.n1054 dvss.n1053 184.572
R3358 dvss.n3142 dvss.n2646 184.572
R3359 dvss.n3135 dvss.n2580 184.572
R3360 dvss.n3131 dvss.n2581 184.572
R3361 dvss.n3127 dvss.n2582 184.572
R3362 dvss.n3123 dvss.n2583 184.572
R3363 dvss.n3119 dvss.n2584 184.572
R3364 dvss.n3115 dvss.n2585 184.572
R3365 dvss.n3111 dvss.n2586 184.572
R3366 dvss.n3107 dvss.n2587 184.572
R3367 dvss.n3103 dvss.n2588 184.572
R3368 dvss.n3099 dvss.n2589 184.572
R3369 dvss.n3095 dvss.n2590 184.572
R3370 dvss.n3091 dvss.n2591 184.572
R3371 dvss.n3087 dvss.n2592 184.572
R3372 dvss.n3083 dvss.n2593 184.572
R3373 dvss.n3079 dvss.n2594 184.572
R3374 dvss.n3075 dvss.n2595 184.572
R3375 dvss.n3071 dvss.n2596 184.572
R3376 dvss.n3067 dvss.n2597 184.572
R3377 dvss.n3063 dvss.n2598 184.572
R3378 dvss.n3059 dvss.n2599 184.572
R3379 dvss.n3055 dvss.n2600 184.572
R3380 dvss.n3051 dvss.n2601 184.572
R3381 dvss.n3047 dvss.n2602 184.572
R3382 dvss.n3043 dvss.n2603 184.572
R3383 dvss.n3039 dvss.n2604 184.572
R3384 dvss.n3035 dvss.n2605 184.572
R3385 dvss.n3031 dvss.n2606 184.572
R3386 dvss.n3027 dvss.n2607 184.572
R3387 dvss.n3023 dvss.n2608 184.572
R3388 dvss.n3019 dvss.n2609 184.572
R3389 dvss.n3015 dvss.n2610 184.572
R3390 dvss.n3011 dvss.n2611 184.572
R3391 dvss.n3007 dvss.n2612 184.572
R3392 dvss.n3003 dvss.n2613 184.572
R3393 dvss.n2999 dvss.n2614 184.572
R3394 dvss.n2995 dvss.n2615 184.572
R3395 dvss.n2991 dvss.n2616 184.572
R3396 dvss.n2987 dvss.n2617 184.572
R3397 dvss.n2983 dvss.n2618 184.572
R3398 dvss.n2979 dvss.n2619 184.572
R3399 dvss.n2975 dvss.n2620 184.572
R3400 dvss.n2971 dvss.n2621 184.572
R3401 dvss.n2967 dvss.n2622 184.572
R3402 dvss.n2963 dvss.n2623 184.572
R3403 dvss.n2959 dvss.n2624 184.572
R3404 dvss.n2955 dvss.n2625 184.572
R3405 dvss.n2951 dvss.n2626 184.572
R3406 dvss.n2947 dvss.n2627 184.572
R3407 dvss.n2943 dvss.n2628 184.572
R3408 dvss.n2939 dvss.n2629 184.572
R3409 dvss.n2935 dvss.n2630 184.572
R3410 dvss.n2931 dvss.n2631 184.572
R3411 dvss.n2927 dvss.n2632 184.572
R3412 dvss.n2923 dvss.n2633 184.572
R3413 dvss.n2919 dvss.n2634 184.572
R3414 dvss.n2915 dvss.n2635 184.572
R3415 dvss.n2911 dvss.n2636 184.572
R3416 dvss.n2907 dvss.n2637 184.572
R3417 dvss.n2903 dvss.n2638 184.572
R3418 dvss.n2899 dvss.n2639 184.572
R3419 dvss.n2895 dvss.n2640 184.572
R3420 dvss.n2891 dvss.n2641 184.572
R3421 dvss.n2887 dvss.n2642 184.572
R3422 dvss.n2883 dvss.n2643 184.572
R3423 dvss.n2644 dvss.n2579 184.572
R3424 dvss.n3144 dvss.n2576 184.572
R3425 dvss.n2013 dvss.t370 178.282
R3426 dvss.t610 dvss.n3167 178.282
R3427 dvss.n4199 dvss.t697 172.957
R3428 dvss.n197 dvss.t382 172.957
R3429 dvss.n3748 dvss.t411 172.957
R3430 dvss.t350 dvss.n3635 172.957
R3431 dvss.n3516 dvss.t95 172.957
R3432 dvss.n1686 dvss.t431 172.957
R3433 dvss.n1565 dvss.t273 172.957
R3434 dvss.n692 dvss.t392 172.957
R3435 dvss.n1178 dvss.t131 172.957
R3436 dvss.n4078 dvss.t763 171.311
R3437 dvss.n3826 dvss.t12 171.311
R3438 dvss.n3697 dvss.t247 171.311
R3439 dvss.n3578 dvss.t224 171.311
R3440 dvss.n3456 dvss.t398 171.311
R3441 dvss.n1662 dvss.t709 171.311
R3442 dvss.n1505 dvss.t723 171.311
R3443 dvss.n1219 dvss.t113 171.311
R3444 dvss.t195 dvss.n777 171.311
R3445 dvss.n396 dvss.t314 170.308
R3446 dvss.n454 dvss.t317 170.308
R3447 dvss.n574 dvss.t299 170.308
R3448 dvss.n515 dvss.t302 170.308
R3449 dvss.n3353 dvss.t305 170.308
R3450 dvss.n1824 dvss.t308 170.308
R3451 dvss.n1404 dvss.t290 170.308
R3452 dvss.n1341 dvss.t287 170.308
R3453 dvss.n4180 dvss.t619 169.85
R3454 dvss.n4155 dvss.t184 169.85
R3455 dvss.n4198 dvss.t322 169.498
R3456 dvss.n201 dvss.t0 169.498
R3457 dvss.t163 dvss.n3751 169.498
R3458 dvss.t337 dvss.n3636 169.498
R3459 dvss.t315 dvss.n3519 169.498
R3460 dvss.n1689 dvss.t318 169.498
R3461 dvss.t303 dvss.n1568 169.498
R3462 dvss.n695 dvss.t300 169.498
R3463 dvss.t401 dvss.n1181 169.498
R3464 dvss.t259 dvss.n986 167.899
R3465 dvss.n1306 dvss.t713 166.838
R3466 dvss.n3985 dvss.t683 166.838
R3467 dvss.n3920 dvss.t145 166.838
R3468 dvss.n1996 dvss.t471 166.838
R3469 dvss.n1971 dvss.t18 166.838
R3470 dvss.n1944 dvss.t484 166.838
R3471 dvss.n1789 dvss.t437 166.838
R3472 dvss.n1387 dvss.t103 166.838
R3473 dvss.t643 dvss.n962 166.838
R3474 dvss.t759 dvss.n4168 166.689
R3475 dvss.t370 dvss.n2007 164.019
R3476 dvss.n3170 dvss.t610 164.019
R3477 dvss.n2219 dvss.t453 162.823
R3478 dvss.t322 dvss.n4197 162.579
R3479 dvss.n207 dvss.t0 162.579
R3480 dvss.n3752 dvss.t163 162.579
R3481 dvss.n3640 dvss.t337 162.579
R3482 dvss.n3520 dvss.t315 162.579
R3483 dvss.n1692 dvss.t318 162.579
R3484 dvss.n1569 dvss.t303 162.579
R3485 dvss.n698 dvss.t300 162.579
R3486 dvss.n1182 dvss.t401 162.579
R3487 dvss.n4113 dvss 161.882
R3488 dvss.n3857 dvss 161.882
R3489 dvss.n300 dvss 161.882
R3490 dvss.n3589 dvss 161.882
R3491 dvss.n428 dvss 161.882
R3492 dvss.n1726 dvss 161.882
R3493 dvss.n547 dvss 161.882
R3494 dvss.n1228 dvss 161.882
R3495 dvss.n1133 dvss 161.882
R3496 dvss.n3968 dvss 161.882
R3497 dvss.n3913 dvss 161.882
R3498 dvss.n1904 dvss 161.882
R3499 dvss.n1873 dvss 161.882
R3500 dvss.n1842 dvss 161.882
R3501 dvss.n1782 dvss 161.882
R3502 dvss.n1359 dvss 161.882
R3503 dvss.n1299 dvss 161.882
R3504 dvss.n912 dvss 161.882
R3505 dvss.n2123 dvss 161.882
R3506 dvss.t681 dvss.n3982 161.857
R3507 dvss.n3906 dvss.t143 161.857
R3508 dvss.t469 dvss.n1993 161.857
R3509 dvss.t16 dvss.n1968 161.857
R3510 dvss.t488 dvss.n1941 161.857
R3511 dvss.n1775 dvss.t439 161.857
R3512 dvss.t105 dvss.n1384 161.857
R3513 dvss.n1292 dvss.t711 161.857
R3514 dvss.t639 dvss.n897 161.857
R3515 dvss.n2319 dvss.t736 161.522
R3516 dvss.n2287 dvss.t674 161.522
R3517 dvss.n2390 dvss.t86 161.47
R3518 dvss.n2195 dvss.n2171 161.345
R3519 dvss.n2196 dvss.n2195 161.345
R3520 dvss.n2197 dvss.n2196 161.345
R3521 dvss.n2197 dvss.n2166 161.345
R3522 dvss.n2206 dvss.n2166 161.345
R3523 dvss.n2207 dvss.n2206 161.345
R3524 dvss.n2236 dvss.n2207 161.345
R3525 dvss.n2248 dvss.n2247 161.345
R3526 dvss.n2266 dvss.n2265 161.345
R3527 dvss.n2267 dvss.n2266 161.345
R3528 dvss.n2267 dvss.n2145 161.345
R3529 dvss.n2518 dvss.n2145 161.345
R3530 dvss.n2454 dvss.t517 161.143
R3531 dvss.n816 dvss.t258 160.064
R3532 dvss.n866 dvss.t264 160.064
R3533 dvss.n996 dvss.n995 157.238
R3534 dvss.n4004 dvss.t707 154.8
R3535 dvss.n3936 dvss.t376 154.8
R3536 dvss.n3245 dvss.t407 154.8
R3537 dvss.n1978 dvss.t348 154.8
R3538 dvss.n1953 dvss.t91 154.8
R3539 dvss.n1805 dvss.t423 154.8
R3540 dvss.n1396 dvss.t271 154.8
R3541 dvss.n1322 dvss.t386 154.8
R3542 dvss.t125 dvss.n904 154.8
R3543 dvss.n397 dvss 154.56
R3544 dvss.n455 dvss 154.56
R3545 dvss.n575 dvss 154.56
R3546 dvss.n516 dvss 154.56
R3547 dvss.n3354 dvss 154.56
R3548 dvss.n1825 dvss 154.56
R3549 dvss.n1405 dvss 154.56
R3550 dvss.n1342 dvss 154.56
R3551 dvss.n1030 dvss.t251 154.305
R3552 dvss.n857 dvss.t726 154.305
R3553 dvss.n398 dvss.n397 153.462
R3554 dvss.n456 dvss.n455 153.462
R3555 dvss.n576 dvss.n575 153.462
R3556 dvss.n517 dvss.n516 153.462
R3557 dvss.n3355 dvss.n3354 153.462
R3558 dvss.n1826 dvss.n1825 153.462
R3559 dvss.n1406 dvss.n1405 153.462
R3560 dvss.n1343 dvss.n1342 153.462
R3561 dvss.t312 dvss.t477 153.21
R3562 dvss.n2340 dvss.t746 152.838
R3563 dvss.n2379 dvss.t64 152.838
R3564 dvss.n2276 dvss.t652 152.838
R3565 dvss.n2446 dvss.t503 152.838
R3566 dvss.n2227 dvss.t524 151.867
R3567 dvss.n4095 dvss.t465 148.743
R3568 dvss.n3799 dvss.t43 148.743
R3569 dvss.n3726 dvss.t10 148.743
R3570 dvss.t245 dvss.n359 148.743
R3571 dvss.n3494 dvss.t204 148.743
R3572 dvss.n1680 dvss.t325 148.743
R3573 dvss.n1543 dvss.t214 148.743
R3574 dvss.n686 dvss.t226 148.743
R3575 dvss.n1161 dvss.t28 148.743
R3576 dvss.n2440 dvss.n2439 146.25
R3577 dvss.n2441 dvss.n2440 146.25
R3578 dvss.n2370 dvss.n2369 146.25
R3579 dvss.n2369 dvss.n2365 146.25
R3580 dvss.n2235 dvss.t526 144.538
R3581 dvss.t186 dvss.n104 143.697
R3582 dvss.n4185 dvss.t615 143.697
R3583 dvss.n2251 dvss.n2250 140.614
R3584 dvss.n2233 dvss.n2219 140.103
R3585 dvss.t459 dvss.n175 139.755
R3586 dvss.n3830 dvss.t37 139.755
R3587 dvss.n3701 dvss.t4 139.755
R3588 dvss.n3583 dvss.t239 139.755
R3589 dvss.t212 dvss.n431 139.755
R3590 dvss.t329 dvss.n1640 139.755
R3591 dvss.t220 dvss.n550 139.755
R3592 dvss.t230 dvss.n1249 139.755
R3593 dvss.t26 dvss.n762 139.755
R3594 dvss.n821 dvss.t564 139.52
R3595 dvss.n2658 dvss.t118 139.52
R3596 dvss.n3987 dvss.t687 139.059
R3597 dvss.n3921 dvss.t149 139.059
R3598 dvss.t475 dvss.n3240 139.059
R3599 dvss.t22 dvss.n1973 139.059
R3600 dvss.t480 dvss.n1948 139.059
R3601 dvss.n1790 dvss.t435 139.059
R3602 dvss.t109 dvss.n1391 139.059
R3603 dvss.n1307 dvss.t717 139.059
R3604 dvss.n956 dvss.t641 139.059
R3605 dvss.n816 dvss.t256 137.442
R3606 dvss.n817 dvss.t254 137.442
R3607 dvss.n866 dvss.t262 137.442
R3608 dvss.n867 dvss.t260 137.442
R3609 dvss.n173 dvss.t465 134.488
R3610 dvss.n3838 dvss.t43 134.488
R3611 dvss.n3722 dvss.t10 134.488
R3612 dvss.n3606 dvss.t245 134.488
R3613 dvss.n3490 dvss.t204 134.488
R3614 dvss.n1638 dvss.t325 134.488
R3615 dvss.n1539 dvss.t214 134.488
R3616 dvss.t226 dvss.n684 134.488
R3617 dvss.n1144 dvss.t28 134.488
R3618 dvss.t186 dvss.n105 132.202
R3619 dvss.t461 dvss.n4087 130.738
R3620 dvss.n3833 dvss.t39 130.738
R3621 dvss.n305 dvss.t6 130.738
R3622 dvss.n3582 dvss.t241 130.738
R3623 dvss.n3470 dvss.t208 130.738
R3624 dvss.t327 dvss.n1671 130.738
R3625 dvss.n1519 dvss.t218 130.738
R3626 dvss.n1248 dvss.t232 130.738
R3627 dvss.t30 dvss.n1139 130.738
R3628 dvss.t538 dvss.n4007 128.564
R3629 dvss.t139 dvss.n3949 128.564
R3630 dvss.t761 dvss.n3248 128.564
R3631 dvss.t151 dvss.n1981 128.564
R3632 dvss.t306 dvss.n1956 128.564
R3633 dvss.t309 dvss.n1818 128.564
R3634 dvss.t291 dvss.n1399 128.564
R3635 dvss.t288 dvss.n1335 128.564
R3636 dvss.n945 dvss.t335 128.564
R3637 dvss.t625 dvss.n4198 127.987
R3638 dvss.n201 dvss.t180 127.987
R3639 dvss.n3751 dvss.t366 127.987
R3640 dvss.n3636 dvss.t608 127.987
R3641 dvss.n3519 dvss.t417 127.987
R3642 dvss.n1689 dvss.t45 127.987
R3643 dvss.n1568 dvss.t356 127.987
R3644 dvss.n695 dvss.t582 127.987
R3645 dvss.n1181 dvss.t197 127.987
R3646 dvss.t532 dvss.n2234 125.389
R3647 dvss.n4187 dvss.t617 125.389
R3648 dvss.n4152 dvss.t182 125.389
R3649 dvss.n4008 dvss.t538 123.316
R3650 dvss.n3950 dvss.t139 123.316
R3651 dvss.n3249 dvss.t761 123.316
R3652 dvss.n1982 dvss.t151 123.316
R3653 dvss.n1957 dvss.t306 123.316
R3654 dvss.n1819 dvss.t309 123.316
R3655 dvss.n1400 dvss.t291 123.316
R3656 dvss.n1336 dvss.t288 123.316
R3657 dvss.t335 dvss.n944 123.316
R3658 dvss.t530 dvss.n2249 120.108
R3659 dvss.t532 dvss.n2235 117.647
R3660 dvss.n2212 dvss.t447 117.385
R3661 dvss.n4216 dvss.t702 116.939
R3662 dvss.n4134 dvss.t381 116.939
R3663 dvss.n3765 dvss.t414 116.939
R3664 dvss.n3651 dvss.t353 116.939
R3665 dvss.n3534 dvss.t90 116.939
R3666 dvss.n3415 dvss.t428 116.939
R3667 dvss.n1582 dvss.t270 116.939
R3668 dvss.n1466 dvss.t389 116.939
R3669 dvss.n1196 dvss.t128 116.939
R3670 dvss.n4322 dvss.t620 116.939
R3671 dvss.n4369 dvss.t185 116.939
R3672 dvss.n2074 dvss.t373 116.939
R3673 dvss.n3179 dvss.t613 116.939
R3674 dvss.n2864 dvss.t416 116.939
R3675 dvss.n2825 dvss.t49 116.939
R3676 dvss.n2786 dvss.t355 116.939
R3677 dvss.n2747 dvss.t584 116.939
R3678 dvss.n2708 dvss.t199 116.939
R3679 dvss.n2260 dvss.t523 116.939
R3680 dvss.n4104 dvss.t466 116.938
R3681 dvss.n3848 dvss.t44 116.938
R3682 dvss.n3731 dvss.t11 116.938
R3683 dvss.n3615 dvss.t246 116.938
R3684 dvss.n3499 dvss.t205 116.938
R3685 dvss.n1717 dvss.t326 116.938
R3686 dvss.n1548 dvss.t215 116.938
R3687 dvss.n1236 dvss.t227 116.938
R3688 dvss.n1155 dvss.t29 116.938
R3689 dvss.n4031 dvss.t688 116.938
R3690 dvss.n3929 dvss.t150 116.938
R3691 dvss.n3269 dvss.t476 116.938
R3692 dvss.n3319 dvss.t23 116.938
R3693 dvss.n3374 dvss.t481 116.938
R3694 dvss.n1798 dvss.t436 116.938
R3695 dvss.n1425 dvss.t110 116.938
R3696 dvss.n1315 dvss.t718 116.938
R3697 dvss.n923 dvss.t642 116.938
R3698 dvss.n2547 dvss.t454 116.938
R3699 dvss.n1162 dvss.t47 116.547
R3700 dvss.n1389 dvss.t47 116.547
R3701 dvss.n1946 dvss.t47 116.547
R3702 dvss.n1681 dvss.t47 116.547
R3703 dvss.n687 dvss.t47 116.547
R3704 dvss dvss.n4204 113.316
R3705 dvss dvss.n132 113.316
R3706 dvss dvss.n3739 113.316
R3707 dvss dvss.n3628 113.316
R3708 dvss dvss.n3507 113.316
R3709 dvss dvss.n1629 113.316
R3710 dvss dvss.n1556 113.316
R3711 dvss dvss.n674 113.316
R3712 dvss dvss.n1169 113.316
R3713 dvss dvss.n3995 113.316
R3714 dvss dvss.n226 113.316
R3715 dvss dvss.n1915 113.316
R3716 dvss dvss.n1884 113.316
R3717 dvss dvss.n1853 113.316
R3718 dvss dvss.n472 113.316
R3719 dvss dvss.n1370 113.316
R3720 dvss dvss.n592 113.316
R3721 dvss dvss.n932 113.316
R3722 dvss dvss.n2134 113.316
R3723 dvss.n4001 dvss.t687 112.822
R3724 dvss.n3934 dvss.t149 112.822
R3725 dvss.n3242 dvss.t475 112.822
R3726 dvss.n1975 dvss.t22 112.822
R3727 dvss.n1950 dvss.t480 112.822
R3728 dvss.n1803 dvss.t435 112.822
R3729 dvss.n1393 dvss.t109 112.822
R3730 dvss.n1320 dvss.t717 112.822
R3731 dvss.n953 dvss.t641 112.822
R3732 dvss.t449 dvss.n2213 109.811
R3733 dvss.n4169 dvss.t759 109.21
R3734 dvss.n3153 dvss.n2575 108.963
R3735 dvss.n2249 dvss.t522 108.389
R3736 dvss.n1066 dvss.n1058 105.862
R3737 dvss.n882 dvss.n880 105.862
R3738 dvss.t615 dvss.n4182 105.582
R3739 dvss.n397 dvss.n396 101.513
R3740 dvss.n455 dvss.n454 101.513
R3741 dvss.n575 dvss.n574 101.513
R3742 dvss.n516 dvss.n515 101.513
R3743 dvss.n3354 dvss.n3353 101.513
R3744 dvss.n1825 dvss.n1824 101.513
R3745 dvss.n1405 dvss.n1404 101.513
R3746 dvss.n1342 dvss.n1341 101.513
R3747 dvss.n995 dvss.n994 98.6074
R3748 dvss.n2222 dvss.n2221 98.508
R3749 dvss.n2178 dvss.t320 97.4795
R3750 dvss.n4007 dvss.t707 97.0786
R3751 dvss.n3949 dvss.t376 97.0786
R3752 dvss.n3248 dvss.t407 97.0786
R3753 dvss.n1981 dvss.t348 97.0786
R3754 dvss.n1956 dvss.t91 97.0786
R3755 dvss.n1818 dvss.t423 97.0786
R3756 dvss.n1399 dvss.t271 97.0786
R3757 dvss.n1335 dvss.t386 97.0786
R3758 dvss.n945 dvss.t125 97.0786
R3759 dvss.n2179 dvss.n2178 95.7988
R3760 dvss.n3225 dvss.t368 92.7071
R3761 dvss.n3155 dvss.t602 92.7071
R3762 dvss.n153 dvss.n152 90.0716
R3763 dvss.n3779 dvss.n3778 90.0716
R3764 dvss.n3682 dvss.n3681 90.0716
R3765 dvss.n3569 dvss.n3568 90.0716
R3766 dvss.n3450 dvss.n3449 90.0716
R3767 dvss.n1596 dvss.n1595 90.0716
R3768 dvss.n1499 dvss.n1498 90.0716
R3769 dvss.n1212 dvss.n1211 90.0716
R3770 dvss.n1109 dvss.n1108 90.0716
R3771 dvss.n823 dvss.n822 90.0716
R3772 dvss.n31 dvss.n30 90.0716
R3773 dvss.n2036 dvss.n2035 90.0716
R3774 dvss.n3205 dvss.n3204 90.0716
R3775 dvss.n2875 dvss.n2874 90.0716
R3776 dvss.n2836 dvss.n2835 90.0716
R3777 dvss.n2797 dvss.n2796 90.0716
R3778 dvss.n2758 dvss.n2757 90.0716
R3779 dvss.n2719 dvss.n2718 90.0716
R3780 dvss.n2680 dvss.n2679 90.0716
R3781 dvss.n2660 dvss.n2659 90.0716
R3782 dvss.n2187 dvss.n2186 90.0716
R3783 dvss.n4095 dvss.t699 89.9376
R3784 dvss.n3799 dvss.t378 89.9376
R3785 dvss.n3726 dvss.t409 89.9376
R3786 dvss.n359 dvss.t342 89.9376
R3787 dvss.n3494 dvss.t99 89.9376
R3788 dvss.t433 dvss.n1680 89.9376
R3789 dvss.n1543 dvss.t277 89.9376
R3790 dvss.t396 dvss.n686 89.9376
R3791 dvss.t135 dvss.n1161 89.9376
R3792 dvss.n987 dvss.t259 87.9472
R3793 dvss.n2039 dvss.n259 85.5759
R3794 dvss.n3186 dvss.n3185 85.5759
R3795 dvss.n2435 dvss.t166 84.171
R3796 dvss.t528 dvss.n2248 84.0341
R3797 dvss.n4227 dvss.n4226 83.0194
R3798 dvss.n4067 dvss.n4066 83.0194
R3799 dvss.n3880 dvss.n3879 83.0194
R3800 dvss.n3660 dvss.n327 83.0194
R3801 dvss.n3542 dvss.n389 83.0194
R3802 dvss.n3409 dvss.n445 83.0194
R3803 dvss.n1749 dvss.n1748 83.0194
R3804 dvss.n1460 dvss.n564 83.0194
R3805 dvss.n1266 dvss.n1265 83.0194
R3806 dvss.n3983 dvss.t681 81.3362
R3807 dvss.n241 dvss.t143 81.3362
R3808 dvss.n1994 dvss.t469 81.3362
R3809 dvss.n1969 dvss.t16 81.3362
R3810 dvss.n1942 dvss.t488 81.3362
R3811 dvss.n487 dvss.t439 81.3362
R3812 dvss.n1385 dvss.t105 81.3362
R3813 dvss.n607 dvss.t711 81.3362
R3814 dvss.n964 dvss.t639 81.3362
R3815 dvss.n4269 dvss.n4268 79.7974
R3816 dvss.n2027 dvss.t372 78.4446
R3817 dvss.n3184 dvss.t612 78.4446
R3818 dvss.n4215 dvss.n86 76.7239
R3819 dvss.n4216 dvss.n4215 76.7239
R3820 dvss.n4135 dvss.n137 76.7239
R3821 dvss.n4135 dvss.n4134 76.7239
R3822 dvss.n3764 dvss.n271 76.7239
R3823 dvss.n3765 dvss.n3764 76.7239
R3824 dvss.n3650 dvss.n334 76.7239
R3825 dvss.n3651 dvss.n3650 76.7239
R3826 dvss.n3533 dvss.n402 76.7239
R3827 dvss.n3534 dvss.n3533 76.7239
R3828 dvss.n1624 dvss.n453 76.7239
R3829 dvss.n3415 dvss.n453 76.7239
R3830 dvss.n1581 dvss.n521 76.7239
R3831 dvss.n1582 dvss.n1581 76.7239
R3832 dvss.n669 dvss.n573 76.7239
R3833 dvss.n1466 dvss.n573 76.7239
R3834 dvss.n1194 dvss.n732 76.7239
R3835 dvss.n1196 dvss.n1194 76.7239
R3836 dvss.n4339 dvss.n43 76.7239
R3837 dvss.n4322 dvss.n43 76.7239
R3838 dvss.n4373 dvss.n4370 76.7239
R3839 dvss.n4370 dvss.n4369 76.7239
R3840 dvss.n3232 dvss.n2075 76.7239
R3841 dvss.n2075 dvss.n2074 76.7239
R3842 dvss.n3176 dvss.n2097 76.7239
R3843 dvss.n3179 dvss.n3176 76.7239
R3844 dvss.n2862 dvss.n2857 76.7239
R3845 dvss.n2864 dvss.n2862 76.7239
R3846 dvss.n2823 dvss.n2818 76.7239
R3847 dvss.n2825 dvss.n2823 76.7239
R3848 dvss.n2784 dvss.n2779 76.7239
R3849 dvss.n2786 dvss.n2784 76.7239
R3850 dvss.n2745 dvss.n2740 76.7239
R3851 dvss.n2747 dvss.n2745 76.7239
R3852 dvss.n2706 dvss.n2701 76.7239
R3853 dvss.n2708 dvss.n2706 76.7239
R3854 dvss.n2257 dvss.n2153 76.7239
R3855 dvss.n2260 dvss.n2257 76.7239
R3856 dvss.n4225 dvss.t701 76.1011
R3857 dvss.n215 dvss.t380 76.1011
R3858 dvss.t413 dvss.n260 76.1011
R3859 dvss.t352 dvss.n3638 76.1011
R3860 dvss.t89 dvss.n3522 76.1011
R3861 dvss.n3410 dvss.t427 76.1011
R3862 dvss.t269 dvss.n505 76.1011
R3863 dvss.n1461 dvss.t388 76.1011
R3864 dvss.t127 dvss.n625 76.1011
R3865 dvss.t683 dvss.n3984 76.0887
R3866 dvss.t145 dvss.n3919 76.0887
R3867 dvss.t471 dvss.n1995 76.0887
R3868 dvss.t18 dvss.n1970 76.0887
R3869 dvss.t484 dvss.n1943 76.0887
R3870 dvss.t437 dvss.n1788 76.0887
R3871 dvss.t103 dvss.n1386 76.0887
R3872 dvss.t713 dvss.n1305 76.0887
R3873 dvss.n963 dvss.t643 76.0887
R3874 dvss.n2046 dvss.t182 74.7229
R3875 dvss.t617 dvss.n4178 74.7229
R3876 dvss.n4291 dvss.n4290 73.1255
R3877 dvss.n4290 dvss.n4289 73.1255
R3878 dvss.n4267 dvss.n4248 73.1255
R3879 dvss.n4268 dvss.n4267 73.1255
R3880 dvss dvss.n4113 73.0358
R3881 dvss.n4103 dvss 73.0358
R3882 dvss dvss.n3857 73.0358
R3883 dvss.n3847 dvss 73.0358
R3884 dvss dvss.n300 73.0358
R3885 dvss dvss.n3710 73.0358
R3886 dvss.n3589 dvss 73.0358
R3887 dvss dvss.n3591 73.0358
R3888 dvss dvss.n428 73.0358
R3889 dvss dvss.n3478 73.0358
R3890 dvss dvss.n1726 73.0358
R3891 dvss.n1716 dvss 73.0358
R3892 dvss dvss.n547 73.0358
R3893 dvss dvss.n1527 73.0358
R3894 dvss.n1228 dvss 73.0358
R3895 dvss.n1235 dvss 73.0358
R3896 dvss.n1133 dvss 73.0358
R3897 dvss.n1154 dvss 73.0358
R3898 dvss.n3968 dvss 73.0358
R3899 dvss.n4030 dvss 73.0358
R3900 dvss.n3913 dvss 73.0358
R3901 dvss.n3928 dvss 73.0358
R3902 dvss.n1904 dvss 73.0358
R3903 dvss.n3268 dvss 73.0358
R3904 dvss.n1873 dvss 73.0358
R3905 dvss.n3318 dvss 73.0358
R3906 dvss.n1842 dvss 73.0358
R3907 dvss.n3373 dvss 73.0358
R3908 dvss.n1782 dvss 73.0358
R3909 dvss.n1797 dvss 73.0358
R3910 dvss.n1359 dvss 73.0358
R3911 dvss.n1424 dvss 73.0358
R3912 dvss.n1299 dvss 73.0358
R3913 dvss.n1314 dvss 73.0358
R3914 dvss.n912 dvss 73.0358
R3915 dvss.n920 dvss 73.0358
R3916 dvss.n2123 dvss 73.0358
R3917 dvss.n2546 dvss 73.0358
R3918 dvss.t34 dvss.t324 70.8111
R3919 dvss.t324 dvss.t190 70.8111
R3920 dvss.t190 dvss.t769 70.8111
R3921 dvss.t769 dvss.t768 70.8111
R3922 dvss.t591 dvss.t249 70.8111
R3923 dvss.t765 dvss.t400 70.8111
R3924 dvss.t614 dvss.t765 70.8111
R3925 dvss.n2251 dvss.t528 67.3778
R3926 dvss.n4246 dvss.n4245 66.9177
R3927 dvss.n4253 dvss.n4252 66.9014
R3928 dvss.n4255 dvss.n4251 66.9014
R3929 dvss.n4257 dvss.n4250 66.9014
R3930 dvss.n2372 dvss.n2371 66.771
R3931 dvss.n2436 dvss.n2373 66.771
R3932 dvss.n4259 dvss.n4258 66.6759
R3933 dvss.n180 dvss.t600 64.6673
R3934 dvss.n3818 dvss.t445 64.6673
R3935 dvss.n314 dvss.t766 64.6673
R3936 dvss.n3548 dvss.t191 64.6673
R3937 dvss.n443 dvss.t693 64.6673
R3938 dvss.n1645 dvss.t691 64.6673
R3939 dvss.n562 dvss.t589 64.6673
R3940 dvss.n637 dvss.t628 64.6673
R3941 dvss.t193 dvss.n800 63.9189
R3942 dvss.t320 dvss.n2171 63.866
R3943 dvss.n4158 dvss.t184 63.2272
R3944 dvss.t619 dvss.n79 63.2272
R3945 dvss.n80 dvss.n59 62.9701
R3946 dvss.n4065 dvss.n4064 62.9701
R3947 dvss.n3883 dvss.n3881 62.9701
R3948 dvss.n1987 dvss.n1986 62.9701
R3949 dvss.n1962 dvss.n1961 62.9701
R3950 dvss.n3408 dvss.n3407 62.9701
R3951 dvss.n1752 dvss.n1750 62.9701
R3952 dvss.n1459 dvss.n1458 62.9701
R3953 dvss.n1269 dvss.n1267 62.9701
R3954 dvss.t574 dvss.n4266 57.4543
R3955 dvss.n86 dvss.n85 57.0829
R3956 dvss.n4214 dvss.n88 57.0829
R3957 dvss.n137 dvss.n136 57.0829
R3958 dvss.n4138 dvss.n4136 57.0829
R3959 dvss.n271 dvss.n270 57.0829
R3960 dvss.n3763 dvss.n273 57.0829
R3961 dvss.n334 dvss.n333 57.0829
R3962 dvss.n3649 dvss.n336 57.0829
R3963 dvss.n402 dvss.n401 57.0829
R3964 dvss.n3532 dvss.n404 57.0829
R3965 dvss.n1624 dvss.n1623 57.0829
R3966 dvss.n1702 dvss.n1700 57.0829
R3967 dvss.n521 dvss.n520 57.0829
R3968 dvss.n1580 dvss.n523 57.0829
R3969 dvss.n669 dvss.n668 57.0829
R3970 dvss.n708 dvss.n706 57.0829
R3971 dvss.n732 dvss.n731 57.0829
R3972 dvss.n1193 dvss.n734 57.0829
R3973 dvss.n4339 dvss.n4338 57.0829
R3974 dvss.n4331 dvss.n4330 57.0829
R3975 dvss.n4373 dvss.n4371 57.0829
R3976 dvss.n21 dvss.n20 57.0829
R3977 dvss.n3232 dvss.n2076 57.0829
R3978 dvss.n2003 dvss.n2002 57.0829
R3979 dvss.n2097 dvss.n2096 57.0829
R3980 dvss.n3175 dvss.n2099 57.0829
R3981 dvss.n2857 dvss.n2855 57.0829
R3982 dvss.n2861 dvss.n2859 57.0829
R3983 dvss.n2818 dvss.n2816 57.0829
R3984 dvss.n2822 dvss.n2820 57.0829
R3985 dvss.n2779 dvss.n2777 57.0829
R3986 dvss.n2783 dvss.n2781 57.0829
R3987 dvss.n2740 dvss.n2738 57.0829
R3988 dvss.n2744 dvss.n2742 57.0829
R3989 dvss.n2701 dvss.n2699 57.0829
R3990 dvss.n2705 dvss.n2703 57.0829
R3991 dvss.n2153 dvss.n2152 57.0829
R3992 dvss.n2256 dvss.n2155 57.0829
R3993 dvss.n2045 dvss.t570 57.076
R3994 dvss.n3199 dvss.t721 57.076
R3995 dvss.n3143 dvss.t175 56.4983
R3996 dvss.t400 dvss.n4269 51.5162
R3997 dvss.t364 dvss.n2025 49.9195
R3998 dvss.n3169 dvss.t606 49.9195
R3999 dvss.n4270 dvss.t614 49.3028
R4000 dvss.n4197 dvss.t705 48.4282
R4001 dvss.t384 dvss.n207 48.4282
R4002 dvss.t405 dvss.n3752 48.4282
R4003 dvss.n3640 dvss.t346 48.4282
R4004 dvss.t93 dvss.n3520 48.4282
R4005 dvss.t429 dvss.n1692 48.4282
R4006 dvss.t267 dvss.n1569 48.4282
R4007 dvss.t390 dvss.n698 48.4282
R4008 dvss.t129 dvss.n1182 48.4282
R4009 dvss.n163 dvss.n162 46.2505
R4010 dvss.n165 dvss.n164 46.2505
R4011 dvss.n3789 dvss.n3788 46.2505
R4012 dvss.n3791 dvss.n3790 46.2505
R4013 dvss.n3692 dvss.n3688 46.2505
R4014 dvss.n3709 dvss.n3708 46.2505
R4015 dvss.n368 dvss.n367 46.2505
R4016 dvss.n3595 dvss.n3590 46.2505
R4017 dvss.n3463 dvss.n3462 46.2505
R4018 dvss.n3477 dvss.n3476 46.2505
R4019 dvss.n1606 dvss.n1605 46.2505
R4020 dvss.n1608 dvss.n1607 46.2505
R4021 dvss.n1512 dvss.n1511 46.2505
R4022 dvss.n1526 dvss.n1525 46.2505
R4023 dvss.n722 dvss.n721 46.2505
R4024 dvss.n1232 dvss.n1231 46.2505
R4025 dvss.n768 dvss.n767 46.2505
R4026 dvss.n755 dvss.n754 46.2505
R4027 dvss.n4048 dvss.n3962 46.2505
R4028 dvss.n4039 dvss.n3969 46.2505
R4029 dvss.n246 dvss.n245 46.2505
R4030 dvss.n237 dvss.n236 46.2505
R4031 dvss.n3286 dvss.n1899 46.2505
R4032 dvss.n3277 dvss.n1905 46.2505
R4033 dvss.n3336 dvss.n1868 46.2505
R4034 dvss.n3327 dvss.n1874 46.2505
R4035 dvss.n3391 dvss.n1836 46.2505
R4036 dvss.n3382 dvss.n1843 46.2505
R4037 dvss.n492 dvss.n491 46.2505
R4038 dvss.n483 dvss.n482 46.2505
R4039 dvss.n1442 dvss.n1353 46.2505
R4040 dvss.n1433 dvss.n1360 46.2505
R4041 dvss.n612 dvss.n611 46.2505
R4042 dvss.n603 dvss.n602 46.2505
R4043 dvss.n909 dvss.n908 46.2505
R4044 dvss.n917 dvss.n916 46.2505
R4045 dvss.n2564 dvss.n2118 46.2505
R4046 dvss.n2555 dvss.n2124 46.2505
R4047 dvss.n2412 dvss.n2411 45.0005
R4048 dvss.n2438 dvss.n2367 45.0005
R4049 dvss.n2367 dvss.t157 45.0005
R4050 dvss.n2368 dvss.n2366 45.0005
R4051 dvss.t157 dvss.n2366 45.0005
R4052 dvss.n2364 dvss.n2363 45.0005
R4053 dvss.n2493 dvss.n2492 45.0005
R4054 dvss.n4288 dvss.t34 44.9596
R4055 dvss.n4103 dvss 44.424
R4056 dvss.n3847 dvss 44.424
R4057 dvss.n3710 dvss 44.424
R4058 dvss.n3591 dvss 44.424
R4059 dvss.n3478 dvss 44.424
R4060 dvss.n1716 dvss 44.424
R4061 dvss.n1527 dvss 44.424
R4062 dvss.n1235 dvss 44.424
R4063 dvss.n1154 dvss 44.424
R4064 dvss.n4030 dvss 44.424
R4065 dvss.n3928 dvss 44.424
R4066 dvss.n3268 dvss 44.424
R4067 dvss.n3318 dvss 44.424
R4068 dvss.n3373 dvss 44.424
R4069 dvss.n1797 dvss 44.424
R4070 dvss.n1424 dvss 44.424
R4071 dvss.n1314 dvss 44.424
R4072 dvss.n920 dvss 44.424
R4073 dvss.n2546 dvss 44.424
R4074 dvss.n2236 dvss.t532 43.698
R4075 dvss.t567 dvss.n1061 43.2419
R4076 dvss.t120 dvss.n2669 43.2419
R4077 dvss.n3238 dvss.t368 39.2225
R4078 dvss.t602 dvss.n351 39.2225
R4079 dvss.n4187 dvss.t699 38.0508
R4080 dvss.n4152 dvss.t378 38.0508
R4081 dvss.n3238 dvss.t409 38.0508
R4082 dvss.t342 dvss.n351 38.0508
R4083 dvss.n1946 dvss.t99 38.0508
R4084 dvss.n1681 dvss.t433 38.0508
R4085 dvss.n1389 dvss.t277 38.0508
R4086 dvss.n687 dvss.t396 38.0508
R4087 dvss.n1162 dvss.t135 38.0508
R4088 dvss.n1058 dvss.t124 37.7206
R4089 dvss.n880 dvss.t562 37.7206
R4090 dvss.n2265 dvss.t522 36.9753
R4091 dvss.n2486 dvss.n2485 36.563
R4092 dvss.t250 dvss.t252 36.1649
R4093 dvss.n2183 dvss.n2175 36.1417
R4094 dvss.n2183 dvss.n2176 36.1417
R4095 dvss.n2176 dvss.n2173 36.1417
R4096 dvss.n2193 dvss.n2173 36.1417
R4097 dvss.n2193 dvss.n2169 36.1417
R4098 dvss.n2199 dvss.n2169 36.1417
R4099 dvss.n2199 dvss.n2168 36.1417
R4100 dvss.n2204 dvss.n2168 36.1417
R4101 dvss.n2204 dvss.n2164 36.1417
R4102 dvss.n2238 dvss.n2164 36.1417
R4103 dvss.n2238 dvss.n2163 36.1417
R4104 dvss.n2245 dvss.n2163 36.1417
R4105 dvss.n2245 dvss.n2156 36.1417
R4106 dvss.n2253 dvss.n2156 36.1417
R4107 dvss.n2253 dvss.n2159 36.1417
R4108 dvss.n2159 dvss.n2151 36.1417
R4109 dvss.n2263 dvss.n2151 36.1417
R4110 dvss.n2263 dvss.n2148 36.1417
R4111 dvss.n2269 dvss.n2148 36.1417
R4112 dvss.n2269 dvss.n2147 36.1417
R4113 dvss.n2516 dvss.n2147 36.1417
R4114 dvss.n3141 dvss.n3140 36.1417
R4115 dvss.n3140 dvss.n3139 36.1417
R4116 dvss.n3139 dvss.n3138 36.1417
R4117 dvss.n3138 dvss.n3136 36.1417
R4118 dvss.n3136 dvss.n3133 36.1417
R4119 dvss.n3133 dvss.n3132 36.1417
R4120 dvss.n3132 dvss.n3129 36.1417
R4121 dvss.n3129 dvss.n3128 36.1417
R4122 dvss.n3128 dvss.n3125 36.1417
R4123 dvss.n3125 dvss.n3124 36.1417
R4124 dvss.n3124 dvss.n3121 36.1417
R4125 dvss.n3121 dvss.n3120 36.1417
R4126 dvss.n3120 dvss.n3117 36.1417
R4127 dvss.n3117 dvss.n3116 36.1417
R4128 dvss.n3116 dvss.n3113 36.1417
R4129 dvss.n3113 dvss.n3112 36.1417
R4130 dvss.n3109 dvss.n3108 36.1417
R4131 dvss.n3108 dvss.n3105 36.1417
R4132 dvss.n3105 dvss.n3104 36.1417
R4133 dvss.n3104 dvss.n3101 36.1417
R4134 dvss.n3101 dvss.n3100 36.1417
R4135 dvss.n3100 dvss.n3097 36.1417
R4136 dvss.n3097 dvss.n3096 36.1417
R4137 dvss.n3096 dvss.n3093 36.1417
R4138 dvss.n3093 dvss.n3092 36.1417
R4139 dvss.n3092 dvss.n3089 36.1417
R4140 dvss.n3089 dvss.n3088 36.1417
R4141 dvss.n3088 dvss.n3085 36.1417
R4142 dvss.n3085 dvss.n3084 36.1417
R4143 dvss.n3084 dvss.n3081 36.1417
R4144 dvss.n3081 dvss.n3080 36.1417
R4145 dvss.n3080 dvss.n3077 36.1417
R4146 dvss.n3077 dvss.n3076 36.1417
R4147 dvss.n3076 dvss.n3073 36.1417
R4148 dvss.n3073 dvss.n3072 36.1417
R4149 dvss.n3072 dvss.n3069 36.1417
R4150 dvss.n3069 dvss.n3068 36.1417
R4151 dvss.n3065 dvss.n3064 36.1417
R4152 dvss.n3064 dvss.n3061 36.1417
R4153 dvss.n3061 dvss.n3060 36.1417
R4154 dvss.n3060 dvss.n3057 36.1417
R4155 dvss.n3057 dvss.n3056 36.1417
R4156 dvss.n3056 dvss.n3053 36.1417
R4157 dvss.n3053 dvss.n3052 36.1417
R4158 dvss.n3052 dvss.n3049 36.1417
R4159 dvss.n3049 dvss.n3048 36.1417
R4160 dvss.n3048 dvss.n3045 36.1417
R4161 dvss.n3045 dvss.n3044 36.1417
R4162 dvss.n3044 dvss.n3041 36.1417
R4163 dvss.n3041 dvss.n3040 36.1417
R4164 dvss.n3040 dvss.n3037 36.1417
R4165 dvss.n3037 dvss.n3036 36.1417
R4166 dvss.n3036 dvss.n3033 36.1417
R4167 dvss.n3033 dvss.n3032 36.1417
R4168 dvss.n3032 dvss.n3029 36.1417
R4169 dvss.n3029 dvss.n3028 36.1417
R4170 dvss.n3028 dvss.n3025 36.1417
R4171 dvss.n3025 dvss.n3024 36.1417
R4172 dvss.n3021 dvss.n3020 36.1417
R4173 dvss.n3020 dvss.n3017 36.1417
R4174 dvss.n3017 dvss.n3016 36.1417
R4175 dvss.n3016 dvss.n3013 36.1417
R4176 dvss.n3013 dvss.n3012 36.1417
R4177 dvss.n3012 dvss.n3009 36.1417
R4178 dvss.n3009 dvss.n3008 36.1417
R4179 dvss.n3008 dvss.n3005 36.1417
R4180 dvss.n3005 dvss.n3004 36.1417
R4181 dvss.n3004 dvss.n3001 36.1417
R4182 dvss.n3001 dvss.n3000 36.1417
R4183 dvss.n3000 dvss.n2997 36.1417
R4184 dvss.n2997 dvss.n2996 36.1417
R4185 dvss.n2996 dvss.n2993 36.1417
R4186 dvss.n2993 dvss.n2992 36.1417
R4187 dvss.n2992 dvss.n2989 36.1417
R4188 dvss.n2989 dvss.n2988 36.1417
R4189 dvss.n2988 dvss.n2985 36.1417
R4190 dvss.n2985 dvss.n2984 36.1417
R4191 dvss.n2984 dvss.n2981 36.1417
R4192 dvss.n2981 dvss.n2980 36.1417
R4193 dvss.n2977 dvss.n2976 36.1417
R4194 dvss.n2976 dvss.n2973 36.1417
R4195 dvss.n2973 dvss.n2972 36.1417
R4196 dvss.n2972 dvss.n2969 36.1417
R4197 dvss.n2969 dvss.n2968 36.1417
R4198 dvss.n2968 dvss.n2965 36.1417
R4199 dvss.n2965 dvss.n2964 36.1417
R4200 dvss.n2964 dvss.n2961 36.1417
R4201 dvss.n2961 dvss.n2960 36.1417
R4202 dvss.n2960 dvss.n2957 36.1417
R4203 dvss.n2957 dvss.n2956 36.1417
R4204 dvss.n2956 dvss.n2953 36.1417
R4205 dvss.n2953 dvss.n2952 36.1417
R4206 dvss.n2952 dvss.n2949 36.1417
R4207 dvss.n2949 dvss.n2948 36.1417
R4208 dvss.n2948 dvss.n2945 36.1417
R4209 dvss.n2945 dvss.n2944 36.1417
R4210 dvss.n2944 dvss.n2941 36.1417
R4211 dvss.n2941 dvss.n2940 36.1417
R4212 dvss.n2940 dvss.n2937 36.1417
R4213 dvss.n2937 dvss.n2936 36.1417
R4214 dvss.n2933 dvss.n2932 36.1417
R4215 dvss.n2932 dvss.n2929 36.1417
R4216 dvss.n2929 dvss.n2928 36.1417
R4217 dvss.n2928 dvss.n2925 36.1417
R4218 dvss.n2925 dvss.n2924 36.1417
R4219 dvss.n2924 dvss.n2921 36.1417
R4220 dvss.n2921 dvss.n2920 36.1417
R4221 dvss.n2920 dvss.n2917 36.1417
R4222 dvss.n2917 dvss.n2916 36.1417
R4223 dvss.n2916 dvss.n2913 36.1417
R4224 dvss.n2913 dvss.n2912 36.1417
R4225 dvss.n2912 dvss.n2909 36.1417
R4226 dvss.n2909 dvss.n2908 36.1417
R4227 dvss.n2908 dvss.n2905 36.1417
R4228 dvss.n2905 dvss.n2904 36.1417
R4229 dvss.n2904 dvss.n2901 36.1417
R4230 dvss.n2901 dvss.n2900 36.1417
R4231 dvss.n2900 dvss.n2897 36.1417
R4232 dvss.n2897 dvss.n2896 36.1417
R4233 dvss.n2896 dvss.n2893 36.1417
R4234 dvss.n2893 dvss.n2892 36.1417
R4235 dvss.n2889 dvss.n2888 36.1417
R4236 dvss.n2888 dvss.n2885 36.1417
R4237 dvss.n2885 dvss.n2884 36.1417
R4238 dvss.n2884 dvss.n2881 36.1417
R4239 dvss.n2881 dvss.n2578 36.1417
R4240 dvss.n3146 dvss.n2578 36.1417
R4241 dvss.n3146 dvss.n2577 36.1417
R4242 dvss.n3151 dvss.n2577 36.1417
R4243 dvss.n3151 dvss.n2109 36.1417
R4244 dvss.n3157 dvss.n2109 36.1417
R4245 dvss.n3157 dvss.n2108 36.1417
R4246 dvss.n3164 dvss.n2108 36.1417
R4247 dvss.n3164 dvss.n2100 36.1417
R4248 dvss.n3172 dvss.n2100 36.1417
R4249 dvss.n3172 dvss.n2103 36.1417
R4250 dvss.n2103 dvss.n2095 36.1417
R4251 dvss.n3182 dvss.n2095 36.1417
R4252 dvss.n3182 dvss.n2092 36.1417
R4253 dvss.n3189 dvss.n2092 36.1417
R4254 dvss.n3189 dvss.n2091 36.1417
R4255 dvss.n3194 dvss.n2091 36.1417
R4256 dvss.n3201 dvss.n2087 36.1417
R4257 dvss.n3201 dvss.n2085 36.1417
R4258 dvss.n3210 dvss.n2085 36.1417
R4259 dvss.n3210 dvss.n2082 36.1417
R4260 dvss.n3216 dvss.n2082 36.1417
R4261 dvss.n3216 dvss.n2081 36.1417
R4262 dvss.n3221 dvss.n2081 36.1417
R4263 dvss.n3221 dvss.n2077 36.1417
R4264 dvss.n3228 dvss.n2077 36.1417
R4265 dvss.n3228 dvss.n2000 36.1417
R4266 dvss.n3235 dvss.n2000 36.1417
R4267 dvss.n3235 dvss.n2001 36.1417
R4268 dvss.n2015 dvss.n2001 36.1417
R4269 dvss.n2015 dvss.n2009 36.1417
R4270 dvss.n2023 dvss.n2009 36.1417
R4271 dvss.n2023 dvss.n2010 36.1417
R4272 dvss.n2010 dvss.n2005 36.1417
R4273 dvss.n2071 dvss.n2005 36.1417
R4274 dvss.n2071 dvss.n2070 36.1417
R4275 dvss.n2070 dvss.n2031 36.1417
R4276 dvss.n2066 dvss.n2031 36.1417
R4277 dvss.n2065 dvss.n2034 36.1417
R4278 dvss.n2058 dvss.n2034 36.1417
R4279 dvss.n2058 dvss.n10 36.1417
R4280 dvss.n4387 dvss.n10 36.1417
R4281 dvss.n4387 dvss.n4386 36.1417
R4282 dvss.n4386 dvss.n13 36.1417
R4283 dvss.n4382 dvss.n13 36.1417
R4284 dvss.n4382 dvss.n4381 36.1417
R4285 dvss.n4381 dvss.n16 36.1417
R4286 dvss.n4377 dvss.n16 36.1417
R4287 dvss.n4377 dvss.n4376 36.1417
R4288 dvss.n4376 dvss.n19 36.1417
R4289 dvss.n118 dvss.n19 36.1417
R4290 dvss.n118 dvss.n108 36.1417
R4291 dvss.n112 dvss.n108 36.1417
R4292 dvss.n112 dvss.n102 36.1417
R4293 dvss.n102 dvss.n23 36.1417
R4294 dvss.n4366 dvss.n23 36.1417
R4295 dvss.n4366 dvss.n4365 36.1417
R4296 dvss.n4365 dvss.n26 36.1417
R4297 dvss.n4361 dvss.n26 36.1417
R4298 dvss.n4360 dvss.n29 36.1417
R4299 dvss.n33 dvss.n29 36.1417
R4300 dvss.n4353 dvss.n33 36.1417
R4301 dvss.n4353 dvss.n4352 36.1417
R4302 dvss.n4352 dvss.n36 36.1417
R4303 dvss.n4348 dvss.n36 36.1417
R4304 dvss.n4348 dvss.n4347 36.1417
R4305 dvss.n4347 dvss.n39 36.1417
R4306 dvss.n4343 dvss.n39 36.1417
R4307 dvss.n4343 dvss.n4342 36.1417
R4308 dvss.n4342 dvss.n42 36.1417
R4309 dvss.n4335 dvss.n42 36.1417
R4310 dvss.n4335 dvss.n4334 36.1417
R4311 dvss.n4334 dvss.n47 36.1417
R4312 dvss.n4327 dvss.n47 36.1417
R4313 dvss.n4327 dvss.n4326 36.1417
R4314 dvss.n4326 dvss.n51 36.1417
R4315 dvss.n4319 dvss.n51 36.1417
R4316 dvss.n4319 dvss.n4318 36.1417
R4317 dvss.n4318 dvss.n54 36.1417
R4318 dvss.n4314 dvss.n54 36.1417
R4319 dvss.n835 dvss.n834 36.1417
R4320 dvss.n1049 dvss.n834 36.1417
R4321 dvss.n1049 dvss.n1048 36.1417
R4322 dvss.n1048 dvss.n1047 36.1417
R4323 dvss.n1047 dvss.n1046 36.1417
R4324 dvss.n1046 dvss.n1044 36.1417
R4325 dvss.n1044 dvss.n1041 36.1417
R4326 dvss.n1041 dvss.n1040 36.1417
R4327 dvss.n1040 dvss.n1037 36.1417
R4328 dvss.n1037 dvss.n1036 36.1417
R4329 dvss.n1036 dvss.n826 36.1417
R4330 dvss.n1055 dvss.n826 36.1417
R4331 dvss.n1055 dvss.n784 36.1417
R4332 dvss.n1100 dvss.n784 36.1417
R4333 dvss.n1100 dvss.n1099 36.1417
R4334 dvss.n1099 dvss.n780 36.1417
R4335 dvss.n1106 dvss.n780 36.1417
R4336 dvss.n1106 dvss.n773 36.1417
R4337 dvss.n1119 dvss.n773 36.1417
R4338 dvss.n1120 dvss.n1119 36.1417
R4339 dvss.n1120 dvss.n769 36.1417
R4340 dvss.n1129 dvss.n769 36.1417
R4341 dvss.n1129 dvss.n765 36.1417
R4342 dvss.n765 dvss.n761 36.1417
R4343 dvss.n761 dvss.n756 36.1417
R4344 dvss.n1143 dvss.n756 36.1417
R4345 dvss.n1143 dvss.n747 36.1417
R4346 dvss.n1165 dvss.n747 36.1417
R4347 dvss.n1166 dvss.n1165 36.1417
R4348 dvss.n1166 dvss.n743 36.1417
R4349 dvss.n743 dvss.n735 36.1417
R4350 dvss.n740 dvss.n735 36.1417
R4351 dvss.n1186 dvss.n740 36.1417
R4352 dvss.n1186 dvss.n630 36.1417
R4353 dvss.n1263 dvss.n630 36.1417
R4354 dvss.n1263 dvss.n1262 36.1417
R4355 dvss.n1262 dvss.n1261 36.1417
R4356 dvss.n1261 dvss.n634 36.1417
R4357 dvss.n1209 dvss.n634 36.1417
R4358 dvss.n1209 dvss.n641 36.1417
R4359 dvss.n1254 dvss.n641 36.1417
R4360 dvss.n1254 dvss.n1253 36.1417
R4361 dvss.n1253 dvss.n1252 36.1417
R4362 dvss.n1252 dvss.n645 36.1417
R4363 dvss.n1246 dvss.n645 36.1417
R4364 dvss.n1246 dvss.n1245 36.1417
R4365 dvss.n1245 dvss.n1244 36.1417
R4366 dvss.n1244 dvss.n654 36.1417
R4367 dvss.n681 dvss.n654 36.1417
R4368 dvss.n681 dvss.n664 36.1417
R4369 dvss.n671 dvss.n664 36.1417
R4370 dvss.n672 dvss.n671 36.1417
R4371 dvss.n680 dvss.n672 36.1417
R4372 dvss.n680 dvss.n676 36.1417
R4373 dvss.n676 dvss.n579 36.1417
R4374 dvss.n1463 dvss.n579 36.1417
R4375 dvss.n1463 dvss.n568 36.1417
R4376 dvss.n1488 dvss.n568 36.1417
R4377 dvss.n1488 dvss.n1487 36.1417
R4378 dvss.n1487 dvss.n570 36.1417
R4379 dvss.n1481 dvss.n570 36.1417
R4380 dvss.n1481 dvss.n559 36.1417
R4381 dvss.n559 dvss.n557 36.1417
R4382 dvss.n1503 dvss.n557 36.1417
R4383 dvss.n1503 dvss.n553 36.1417
R4384 dvss.n1516 dvss.n553 36.1417
R4385 dvss.n1516 dvss.n545 36.1417
R4386 dvss.n1531 dvss.n545 36.1417
R4387 dvss.n1532 dvss.n1531 36.1417
R4388 dvss.n1532 dvss.n542 36.1417
R4389 dvss.n542 dvss.n536 36.1417
R4390 dvss.n1552 dvss.n536 36.1417
R4391 dvss.n1553 dvss.n1552 36.1417
R4392 dvss.n1553 dvss.n532 36.1417
R4393 dvss.n532 dvss.n524 36.1417
R4394 dvss.n529 dvss.n524 36.1417
R4395 dvss.n1573 dvss.n529 36.1417
R4396 dvss.n1573 dvss.n510 36.1417
R4397 dvss.n1746 dvss.n510 36.1417
R4398 dvss.n1746 dvss.n511 36.1417
R4399 dvss.n1588 dvss.n511 36.1417
R4400 dvss.n1589 dvss.n1588 36.1417
R4401 dvss.n1593 dvss.n1589 36.1417
R4402 dvss.n1594 dvss.n1593 36.1417
R4403 dvss.n1659 dvss.n1594 36.1417
R4404 dvss.n1659 dvss.n1598 36.1417
R4405 dvss.n1603 dvss.n1598 36.1417
R4406 dvss.n1666 dvss.n1603 36.1417
R4407 dvss.n1669 dvss.n1666 36.1417
R4408 dvss.n1669 dvss.n1609 36.1417
R4409 dvss.n1614 dvss.n1609 36.1417
R4410 dvss.n1615 dvss.n1614 36.1417
R4411 dvss.n1636 dvss.n1615 36.1417
R4412 dvss.n1636 dvss.n1618 36.1417
R4413 dvss.n1626 dvss.n1618 36.1417
R4414 dvss.n1627 dvss.n1626 36.1417
R4415 dvss.n1635 dvss.n1627 36.1417
R4416 dvss.n1635 dvss.n1631 36.1417
R4417 dvss.n1631 dvss.n459 36.1417
R4418 dvss.n3412 dvss.n459 36.1417
R4419 dvss.n3412 dvss.n449 36.1417
R4420 dvss.n3439 dvss.n449 36.1417
R4421 dvss.n3439 dvss.n450 36.1417
R4422 dvss.n3426 dvss.n450 36.1417
R4423 dvss.n3432 dvss.n3426 36.1417
R4424 dvss.n3432 dvss.n440 36.1417
R4425 dvss.n440 dvss.n438 36.1417
R4426 dvss.n3454 dvss.n438 36.1417
R4427 dvss.n3454 dvss.n434 36.1417
R4428 dvss.n3467 dvss.n434 36.1417
R4429 dvss.n3467 dvss.n426 36.1417
R4430 dvss.n3482 dvss.n426 36.1417
R4431 dvss.n3483 dvss.n3482 36.1417
R4432 dvss.n3483 dvss.n423 36.1417
R4433 dvss.n423 dvss.n417 36.1417
R4434 dvss.n3503 dvss.n417 36.1417
R4435 dvss.n3504 dvss.n3503 36.1417
R4436 dvss.n3504 dvss.n413 36.1417
R4437 dvss.n413 dvss.n405 36.1417
R4438 dvss.n410 dvss.n405 36.1417
R4439 dvss.n3525 dvss.n410 36.1417
R4440 dvss.n3525 dvss.n391 36.1417
R4441 dvss.n3540 dvss.n391 36.1417
R4442 dvss.n3540 dvss.n385 36.1417
R4443 dvss.n3559 dvss.n385 36.1417
R4444 dvss.n3559 dvss.n386 36.1417
R4445 dvss.n386 dvss.n379 36.1417
R4446 dvss.n3565 dvss.n379 36.1417
R4447 dvss.n3565 dvss.n374 36.1417
R4448 dvss.n3576 dvss.n374 36.1417
R4449 dvss.n3576 dvss.n369 36.1417
R4450 dvss.n3585 dvss.n369 36.1417
R4451 dvss.n3585 dvss.n364 36.1417
R4452 dvss.n3602 dvss.n364 36.1417
R4453 dvss.n3602 dvss.n357 36.1417
R4454 dvss.n3609 dvss.n357 36.1417
R4455 dvss.n3609 dvss.n353 36.1417
R4456 dvss.n3619 dvss.n353 36.1417
R4457 dvss.n3619 dvss.n348 36.1417
R4458 dvss.n3633 dvss.n348 36.1417
R4459 dvss.n3633 dvss.n337 36.1417
R4460 dvss.n3642 dvss.n337 36.1417
R4461 dvss.n3642 dvss.n331 36.1417
R4462 dvss.n3654 dvss.n331 36.1417
R4463 dvss.n3655 dvss.n3654 36.1417
R4464 dvss.n3655 dvss.n326 36.1417
R4465 dvss.n326 dvss.n319 36.1417
R4466 dvss.n320 dvss.n319 36.1417
R4467 dvss.n3668 dvss.n320 36.1417
R4468 dvss.n3668 dvss.n310 36.1417
R4469 dvss.n3686 dvss.n310 36.1417
R4470 dvss.n3687 dvss.n3686 36.1417
R4471 dvss.n3687 dvss.n307 36.1417
R4472 dvss.n307 dvss.n301 36.1417
R4473 dvss.n301 dvss.n296 36.1417
R4474 dvss.n3718 dvss.n296 36.1417
R4475 dvss.n3718 dvss.n297 36.1417
R4476 dvss.n297 dvss.n292 36.1417
R4477 dvss.n292 dvss.n286 36.1417
R4478 dvss.n3735 dvss.n286 36.1417
R4479 dvss.n3736 dvss.n3735 36.1417
R4480 dvss.n3736 dvss.n282 36.1417
R4481 dvss.n282 dvss.n274 36.1417
R4482 dvss.n279 dvss.n274 36.1417
R4483 dvss.n3756 dvss.n279 36.1417
R4484 dvss.n3756 dvss.n265 36.1417
R4485 dvss.n3877 dvss.n265 36.1417
R4486 dvss.n3877 dvss.n266 36.1417
R4487 dvss.n3771 dvss.n266 36.1417
R4488 dvss.n3772 dvss.n3771 36.1417
R4489 dvss.n3776 dvss.n3772 36.1417
R4490 dvss.n3777 dvss.n3776 36.1417
R4491 dvss.n3808 dvss.n3777 36.1417
R4492 dvss.n3808 dvss.n3781 36.1417
R4493 dvss.n3786 dvss.n3781 36.1417
R4494 dvss.n3804 dvss.n3786 36.1417
R4495 dvss.n3807 dvss.n3804 36.1417
R4496 dvss.n3807 dvss.n3792 36.1417
R4497 dvss.n3797 dvss.n3792 36.1417
R4498 dvss.n3841 dvss.n3797 36.1417
R4499 dvss.n3841 dvss.n125 36.1417
R4500 dvss.n4149 dvss.n125 36.1417
R4501 dvss.n4149 dvss.n126 36.1417
R4502 dvss.n130 dvss.n126 36.1417
R4503 dvss.n203 dvss.n130 36.1417
R4504 dvss.n205 dvss.n203 36.1417
R4505 dvss.n205 dvss.n192 36.1417
R4506 dvss.n213 dvss.n192 36.1417
R4507 dvss.n213 dvss.n139 36.1417
R4508 dvss.n144 dvss.n139 36.1417
R4509 dvss.n145 dvss.n144 36.1417
R4510 dvss.n146 dvss.n145 36.1417
R4511 dvss.n150 dvss.n146 36.1417
R4512 dvss.n151 dvss.n150 36.1417
R4513 dvss.n4075 dvss.n151 36.1417
R4514 dvss.n4075 dvss.n155 36.1417
R4515 dvss.n160 dvss.n155 36.1417
R4516 dvss.n4082 dvss.n160 36.1417
R4517 dvss.n4085 dvss.n4082 36.1417
R4518 dvss.n4085 dvss.n166 36.1417
R4519 dvss.n171 dvss.n166 36.1417
R4520 dvss.n172 dvss.n171 36.1417
R4521 dvss.n172 dvss.n99 36.1417
R4522 dvss.n4190 dvss.n99 36.1417
R4523 dvss.n4190 dvss.n93 36.1417
R4524 dvss.n4201 dvss.n93 36.1417
R4525 dvss.n4201 dvss.n89 36.1417
R4526 dvss.n89 dvss.n84 36.1417
R4527 dvss.n4220 dvss.n84 36.1417
R4528 dvss.n4220 dvss.n74 36.1417
R4529 dvss.n4229 dvss.n74 36.1417
R4530 dvss.n4229 dvss.n70 36.1417
R4531 dvss.n4235 dvss.n70 36.1417
R4532 dvss.n4235 dvss.n64 36.1417
R4533 dvss.n1009 dvss.n1008 36.1417
R4534 dvss.n1008 dvss.n1007 36.1417
R4535 dvss.n1007 dvss.n843 36.1417
R4536 dvss.n1001 dvss.n843 36.1417
R4537 dvss.n1001 dvss.n1000 36.1417
R4538 dvss.n1000 dvss.n999 36.1417
R4539 dvss.n999 dvss.n851 36.1417
R4540 dvss.n992 dvss.n851 36.1417
R4541 dvss.n992 dvss.n991 36.1417
R4542 dvss.n991 dvss.n990 36.1417
R4543 dvss.n990 dvss.n862 36.1417
R4544 dvss.n984 dvss.n862 36.1417
R4545 dvss.n984 dvss.n983 36.1417
R4546 dvss.n983 dvss.n982 36.1417
R4547 dvss.n982 dvss.n875 36.1417
R4548 dvss.n976 dvss.n875 36.1417
R4549 dvss.n975 dvss.n974 36.1417
R4550 dvss.n974 dvss.n888 36.1417
R4551 dvss.n968 dvss.n888 36.1417
R4552 dvss.n968 dvss.n967 36.1417
R4553 dvss.n967 dvss.n966 36.1417
R4554 dvss.n966 dvss.n895 36.1417
R4555 dvss.n960 dvss.n895 36.1417
R4556 dvss.n960 dvss.n959 36.1417
R4557 dvss.n959 dvss.n958 36.1417
R4558 dvss.n958 dvss.n902 36.1417
R4559 dvss.n906 dvss.n902 36.1417
R4560 dvss.n949 dvss.n906 36.1417
R4561 dvss.n949 dvss.n948 36.1417
R4562 dvss.n948 dvss.n947 36.1417
R4563 dvss.n947 dvss.n929 36.1417
R4564 dvss.n941 dvss.n929 36.1417
R4565 dvss.n941 dvss.n622 36.1417
R4566 dvss.n1271 dvss.n622 36.1417
R4567 dvss.n1271 dvss.n621 36.1417
R4568 dvss.n1276 dvss.n621 36.1417
R4569 dvss.n1276 dvss.n618 36.1417
R4570 dvss.n1282 dvss.n618 36.1417
R4571 dvss.n1282 dvss.n617 36.1417
R4572 dvss.n1288 dvss.n617 36.1417
R4573 dvss.n1288 dvss.n613 36.1417
R4574 dvss.n1294 dvss.n613 36.1417
R4575 dvss.n1294 dvss.n609 36.1417
R4576 dvss.n1303 dvss.n609 36.1417
R4577 dvss.n1303 dvss.n605 36.1417
R4578 dvss.n1310 dvss.n605 36.1417
R4579 dvss.n1310 dvss.n599 36.1417
R4580 dvss.n1318 dvss.n599 36.1417
R4581 dvss.n1318 dvss.n596 36.1417
R4582 dvss.n1325 dvss.n596 36.1417
R4583 dvss.n1325 dvss.n591 36.1417
R4584 dvss.n1333 dvss.n591 36.1417
R4585 dvss.n1333 dvss.n588 36.1417
R4586 dvss.n1339 dvss.n588 36.1417
R4587 dvss.n1339 dvss.n586 36.1417
R4588 dvss.n1456 dvss.n586 36.1417
R4589 dvss.n1456 dvss.n587 36.1417
R4590 dvss.n1452 dvss.n587 36.1417
R4591 dvss.n1452 dvss.n1451 36.1417
R4592 dvss.n1451 dvss.n1349 36.1417
R4593 dvss.n1447 dvss.n1349 36.1417
R4594 dvss.n1447 dvss.n1446 36.1417
R4595 dvss.n1446 dvss.n1352 36.1417
R4596 dvss.n1355 dvss.n1352 36.1417
R4597 dvss.n1438 dvss.n1355 36.1417
R4598 dvss.n1438 dvss.n1437 36.1417
R4599 dvss.n1437 dvss.n1358 36.1417
R4600 dvss.n1429 dvss.n1358 36.1417
R4601 dvss.n1429 dvss.n1428 36.1417
R4602 dvss.n1428 dvss.n1364 36.1417
R4603 dvss.n1421 dvss.n1364 36.1417
R4604 dvss.n1421 dvss.n1420 36.1417
R4605 dvss.n1420 dvss.n1368 36.1417
R4606 dvss.n1372 dvss.n1368 36.1417
R4607 dvss.n1411 dvss.n1372 36.1417
R4608 dvss.n1411 dvss.n1410 36.1417
R4609 dvss.n1410 dvss.n502 36.1417
R4610 dvss.n1754 dvss.n502 36.1417
R4611 dvss.n1754 dvss.n501 36.1417
R4612 dvss.n1759 dvss.n501 36.1417
R4613 dvss.n1759 dvss.n498 36.1417
R4614 dvss.n1765 dvss.n498 36.1417
R4615 dvss.n1765 dvss.n497 36.1417
R4616 dvss.n1771 dvss.n497 36.1417
R4617 dvss.n1771 dvss.n493 36.1417
R4618 dvss.n1777 dvss.n493 36.1417
R4619 dvss.n1777 dvss.n489 36.1417
R4620 dvss.n1786 dvss.n489 36.1417
R4621 dvss.n1786 dvss.n485 36.1417
R4622 dvss.n1793 dvss.n485 36.1417
R4623 dvss.n1793 dvss.n479 36.1417
R4624 dvss.n1801 dvss.n479 36.1417
R4625 dvss.n1801 dvss.n476 36.1417
R4626 dvss.n1808 dvss.n476 36.1417
R4627 dvss.n1808 dvss.n471 36.1417
R4628 dvss.n1816 dvss.n471 36.1417
R4629 dvss.n1816 dvss.n468 36.1417
R4630 dvss.n1822 dvss.n468 36.1417
R4631 dvss.n1822 dvss.n466 36.1417
R4632 dvss.n3405 dvss.n466 36.1417
R4633 dvss.n3405 dvss.n467 36.1417
R4634 dvss.n3401 dvss.n467 36.1417
R4635 dvss.n3401 dvss.n3400 36.1417
R4636 dvss.n3400 dvss.n1832 36.1417
R4637 dvss.n3396 dvss.n1832 36.1417
R4638 dvss.n3396 dvss.n3395 36.1417
R4639 dvss.n3395 dvss.n1835 36.1417
R4640 dvss.n1838 dvss.n1835 36.1417
R4641 dvss.n3387 dvss.n1838 36.1417
R4642 dvss.n3387 dvss.n3386 36.1417
R4643 dvss.n3386 dvss.n1841 36.1417
R4644 dvss.n3378 dvss.n1841 36.1417
R4645 dvss.n3378 dvss.n3377 36.1417
R4646 dvss.n3377 dvss.n1847 36.1417
R4647 dvss.n3370 dvss.n1847 36.1417
R4648 dvss.n3370 dvss.n3369 36.1417
R4649 dvss.n3369 dvss.n1851 36.1417
R4650 dvss.n1855 dvss.n1851 36.1417
R4651 dvss.n3360 dvss.n1855 36.1417
R4652 dvss.n3360 dvss.n3359 36.1417
R4653 dvss.n3359 dvss.n1858 36.1417
R4654 dvss.n3350 dvss.n1858 36.1417
R4655 dvss.n3350 dvss.n3349 36.1417
R4656 dvss.n3349 dvss.n1861 36.1417
R4657 dvss.n3345 dvss.n1861 36.1417
R4658 dvss.n3345 dvss.n3344 36.1417
R4659 dvss.n3344 dvss.n1864 36.1417
R4660 dvss.n3340 dvss.n1864 36.1417
R4661 dvss.n3340 dvss.n3339 36.1417
R4662 dvss.n3339 dvss.n1867 36.1417
R4663 dvss.n3332 dvss.n1867 36.1417
R4664 dvss.n3332 dvss.n3331 36.1417
R4665 dvss.n3331 dvss.n1872 36.1417
R4666 dvss.n3323 dvss.n1872 36.1417
R4667 dvss.n3323 dvss.n3322 36.1417
R4668 dvss.n3322 dvss.n1878 36.1417
R4669 dvss.n3315 dvss.n1878 36.1417
R4670 dvss.n3315 dvss.n3314 36.1417
R4671 dvss.n3314 dvss.n1882 36.1417
R4672 dvss.n1886 dvss.n1882 36.1417
R4673 dvss.n3305 dvss.n1886 36.1417
R4674 dvss.n3305 dvss.n3304 36.1417
R4675 dvss.n3304 dvss.n1889 36.1417
R4676 dvss.n3300 dvss.n1889 36.1417
R4677 dvss.n3300 dvss.n3299 36.1417
R4678 dvss.n3299 dvss.n1892 36.1417
R4679 dvss.n3295 dvss.n1892 36.1417
R4680 dvss.n3295 dvss.n3294 36.1417
R4681 dvss.n3294 dvss.n1895 36.1417
R4682 dvss.n3290 dvss.n1895 36.1417
R4683 dvss.n3290 dvss.n3289 36.1417
R4684 dvss.n3289 dvss.n1898 36.1417
R4685 dvss.n3282 dvss.n1898 36.1417
R4686 dvss.n3282 dvss.n3281 36.1417
R4687 dvss.n3281 dvss.n1903 36.1417
R4688 dvss.n3273 dvss.n1903 36.1417
R4689 dvss.n3273 dvss.n3272 36.1417
R4690 dvss.n3272 dvss.n1909 36.1417
R4691 dvss.n3265 dvss.n1909 36.1417
R4692 dvss.n3265 dvss.n3264 36.1417
R4693 dvss.n3264 dvss.n1913 36.1417
R4694 dvss.n1917 dvss.n1913 36.1417
R4695 dvss.n3255 dvss.n1917 36.1417
R4696 dvss.n3255 dvss.n3254 36.1417
R4697 dvss.n3254 dvss.n256 36.1417
R4698 dvss.n3885 dvss.n256 36.1417
R4699 dvss.n3885 dvss.n255 36.1417
R4700 dvss.n3890 dvss.n255 36.1417
R4701 dvss.n3890 dvss.n252 36.1417
R4702 dvss.n3896 dvss.n252 36.1417
R4703 dvss.n3896 dvss.n251 36.1417
R4704 dvss.n3902 dvss.n251 36.1417
R4705 dvss.n3902 dvss.n247 36.1417
R4706 dvss.n3908 dvss.n247 36.1417
R4707 dvss.n3908 dvss.n243 36.1417
R4708 dvss.n3917 dvss.n243 36.1417
R4709 dvss.n3917 dvss.n239 36.1417
R4710 dvss.n3924 dvss.n239 36.1417
R4711 dvss.n3924 dvss.n233 36.1417
R4712 dvss.n3932 dvss.n233 36.1417
R4713 dvss.n3932 dvss.n230 36.1417
R4714 dvss.n3939 dvss.n230 36.1417
R4715 dvss.n3939 dvss.n225 36.1417
R4716 dvss.n3947 dvss.n225 36.1417
R4717 dvss.n3947 dvss.n222 36.1417
R4718 dvss.n3953 dvss.n222 36.1417
R4719 dvss.n3953 dvss.n220 36.1417
R4720 dvss.n4062 dvss.n220 36.1417
R4721 dvss.n4062 dvss.n221 36.1417
R4722 dvss.n4058 dvss.n221 36.1417
R4723 dvss.n4058 dvss.n4057 36.1417
R4724 dvss.n4057 dvss.n3958 36.1417
R4725 dvss.n4053 dvss.n3958 36.1417
R4726 dvss.n4053 dvss.n4052 36.1417
R4727 dvss.n4052 dvss.n3961 36.1417
R4728 dvss.n3964 dvss.n3961 36.1417
R4729 dvss.n4044 dvss.n3964 36.1417
R4730 dvss.n4044 dvss.n4043 36.1417
R4731 dvss.n4043 dvss.n3967 36.1417
R4732 dvss.n4035 dvss.n3967 36.1417
R4733 dvss.n4035 dvss.n4034 36.1417
R4734 dvss.n4034 dvss.n3989 36.1417
R4735 dvss.n4027 dvss.n3989 36.1417
R4736 dvss.n4027 dvss.n4026 36.1417
R4737 dvss.n4026 dvss.n3993 36.1417
R4738 dvss.n3997 dvss.n3993 36.1417
R4739 dvss.n4017 dvss.n3997 36.1417
R4740 dvss.n4017 dvss.n4016 36.1417
R4741 dvss.n4016 dvss.n4012 36.1417
R4742 dvss.n4012 dvss.n62 36.1417
R4743 dvss.n4307 dvss.n62 36.1417
R4744 dvss.n4307 dvss.n63 36.1417
R4745 dvss.n4303 dvss.n63 36.1417
R4746 dvss.n1019 dvss.n804 36.1417
R4747 dvss.n1088 dvss.n804 36.1417
R4748 dvss.n1088 dvss.n1087 36.1417
R4749 dvss.n1087 dvss.n1086 36.1417
R4750 dvss.n1086 dvss.n1085 36.1417
R4751 dvss.n1085 dvss.n1083 36.1417
R4752 dvss.n1083 dvss.n1080 36.1417
R4753 dvss.n1080 dvss.n1079 36.1417
R4754 dvss.n1079 dvss.n1076 36.1417
R4755 dvss.n1076 dvss.n1075 36.1417
R4756 dvss.n1075 dvss.n1072 36.1417
R4757 dvss.n1072 dvss.n1071 36.1417
R4758 dvss.n1071 dvss.n795 36.1417
R4759 dvss.n795 dvss.n786 36.1417
R4760 dvss.n1096 dvss.n786 36.1417
R4761 dvss.n1096 dvss.n789 36.1417
R4762 dvss.n1114 dvss.n779 36.1417
R4763 dvss.n1115 dvss.n1114 36.1417
R4764 dvss.n1115 dvss.n772 36.1417
R4765 dvss.n1124 dvss.n772 36.1417
R4766 dvss.n1124 dvss.n764 36.1417
R4767 dvss.n1137 dvss.n764 36.1417
R4768 dvss.n1137 dvss.n757 36.1417
R4769 dvss.n1150 dvss.n757 36.1417
R4770 dvss.n1150 dvss.n752 36.1417
R4771 dvss.n1159 dvss.n752 36.1417
R4772 dvss.n1159 dvss.n746 36.1417
R4773 dvss.n1175 dvss.n746 36.1417
R4774 dvss.n1175 dvss.n737 36.1417
R4775 dvss.n1190 dvss.n737 36.1417
R4776 dvss.n1190 dvss.n1189 36.1417
R4777 dvss.n1189 dvss.n729 36.1417
R4778 dvss.n1199 dvss.n729 36.1417
R4779 dvss.n1200 dvss.n1199 36.1417
R4780 dvss.n1201 dvss.n1200 36.1417
R4781 dvss.n1201 dvss.n725 36.1417
R4782 dvss.n1206 dvss.n725 36.1417
R4783 dvss.n1217 dvss.n723 36.1417
R4784 dvss.n1218 dvss.n1217 36.1417
R4785 dvss.n1221 dvss.n1218 36.1417
R4786 dvss.n1222 dvss.n1221 36.1417
R4787 dvss.n1224 dvss.n1222 36.1417
R4788 dvss.n1224 dvss.n1223 36.1417
R4789 dvss.n1223 dvss.n660 36.1417
R4790 dvss.n1240 dvss.n660 36.1417
R4791 dvss.n1240 dvss.n1239 36.1417
R4792 dvss.n1239 dvss.n661 36.1417
R4793 dvss.n717 dvss.n661 36.1417
R4794 dvss.n717 dvss.n716 36.1417
R4795 dvss.n716 dvss.n667 36.1417
R4796 dvss.n677 dvss.n667 36.1417
R4797 dvss.n703 dvss.n677 36.1417
R4798 dvss.n703 dvss.n702 36.1417
R4799 dvss.n702 dvss.n571 36.1417
R4800 dvss.n1469 dvss.n571 36.1417
R4801 dvss.n1470 dvss.n1469 36.1417
R4802 dvss.n1485 dvss.n1470 36.1417
R4803 dvss.n1485 dvss.n1484 36.1417
R4804 dvss.n1495 dvss.n560 36.1417
R4805 dvss.n1495 dvss.n1494 36.1417
R4806 dvss.n1494 dvss.n554 36.1417
R4807 dvss.n1508 dvss.n554 36.1417
R4808 dvss.n1508 dvss.n548 36.1417
R4809 dvss.n1521 dvss.n548 36.1417
R4810 dvss.n1521 dvss.n544 36.1417
R4811 dvss.n1535 dvss.n544 36.1417
R4812 dvss.n1535 dvss.n539 36.1417
R4813 dvss.n1545 dvss.n539 36.1417
R4814 dvss.n1545 dvss.n535 36.1417
R4815 dvss.n1562 dvss.n535 36.1417
R4816 dvss.n1562 dvss.n526 36.1417
R4817 dvss.n1577 dvss.n526 36.1417
R4818 dvss.n1577 dvss.n1576 36.1417
R4819 dvss.n1576 dvss.n513 36.1417
R4820 dvss.n1585 dvss.n513 36.1417
R4821 dvss.n1744 dvss.n1585 36.1417
R4822 dvss.n1744 dvss.n1743 36.1417
R4823 dvss.n1743 dvss.n1587 36.1417
R4824 dvss.n1739 dvss.n1587 36.1417
R4825 dvss.n1738 dvss.n1592 36.1417
R4826 dvss.n1599 dvss.n1592 36.1417
R4827 dvss.n1731 dvss.n1599 36.1417
R4828 dvss.n1731 dvss.n1730 36.1417
R4829 dvss.n1730 dvss.n1602 36.1417
R4830 dvss.n1610 dvss.n1602 36.1417
R4831 dvss.n1722 dvss.n1610 36.1417
R4832 dvss.n1722 dvss.n1721 36.1417
R4833 dvss.n1721 dvss.n1613 36.1417
R4834 dvss.n1619 dvss.n1613 36.1417
R4835 dvss.n1711 dvss.n1619 36.1417
R4836 dvss.n1711 dvss.n1710 36.1417
R4837 dvss.n1710 dvss.n1622 36.1417
R4838 dvss.n1632 dvss.n1622 36.1417
R4839 dvss.n1697 dvss.n1632 36.1417
R4840 dvss.n1697 dvss.n1696 36.1417
R4841 dvss.n1696 dvss.n451 36.1417
R4842 dvss.n3418 dvss.n451 36.1417
R4843 dvss.n3437 dvss.n3418 36.1417
R4844 dvss.n3437 dvss.n3436 36.1417
R4845 dvss.n3436 dvss.n3425 36.1417
R4846 dvss.n3446 dvss.n441 36.1417
R4847 dvss.n3446 dvss.n3445 36.1417
R4848 dvss.n3445 dvss.n435 36.1417
R4849 dvss.n3459 dvss.n435 36.1417
R4850 dvss.n3459 dvss.n429 36.1417
R4851 dvss.n3472 dvss.n429 36.1417
R4852 dvss.n3472 dvss.n425 36.1417
R4853 dvss.n3486 dvss.n425 36.1417
R4854 dvss.n3486 dvss.n420 36.1417
R4855 dvss.n3496 dvss.n420 36.1417
R4856 dvss.n3496 dvss.n416 36.1417
R4857 dvss.n3513 dvss.n416 36.1417
R4858 dvss.n3513 dvss.n407 36.1417
R4859 dvss.n3529 dvss.n407 36.1417
R4860 dvss.n3529 dvss.n3528 36.1417
R4861 dvss.n3528 dvss.n394 36.1417
R4862 dvss.n3537 dvss.n394 36.1417
R4863 dvss.n3538 dvss.n3537 36.1417
R4864 dvss.n3538 dvss.n387 36.1417
R4865 dvss.n3557 dvss.n387 36.1417
R4866 dvss.n3557 dvss.n3556 36.1417
R4867 dvss.n3553 dvss.n377 36.1417
R4868 dvss.n3573 dvss.n377 36.1417
R4869 dvss.n3574 dvss.n3573 36.1417
R4870 dvss.n3574 dvss.n372 36.1417
R4871 dvss.n372 dvss.n365 36.1417
R4872 dvss.n3599 dvss.n365 36.1417
R4873 dvss.n3600 dvss.n3599 36.1417
R4874 dvss.n3600 dvss.n355 36.1417
R4875 dvss.n3611 dvss.n355 36.1417
R4876 dvss.n3612 dvss.n3611 36.1417
R4877 dvss.n3612 dvss.n349 36.1417
R4878 dvss.n3624 dvss.n349 36.1417
R4879 dvss.n3624 dvss.n339 36.1417
R4880 dvss.n3646 dvss.n339 36.1417
R4881 dvss.n3646 dvss.n3645 36.1417
R4882 dvss.n3645 dvss.n342 36.1417
R4883 dvss.n342 dvss.n329 36.1417
R4884 dvss.n3658 dvss.n329 36.1417
R4885 dvss.n3658 dvss.n317 36.1417
R4886 dvss.n3672 dvss.n317 36.1417
R4887 dvss.n3672 dvss.n318 36.1417
R4888 dvss.n3678 dvss.n312 36.1417
R4889 dvss.n3678 dvss.n309 36.1417
R4890 dvss.n3695 dvss.n309 36.1417
R4891 dvss.n3695 dvss.n302 36.1417
R4892 dvss.n3703 dvss.n302 36.1417
R4893 dvss.n3703 dvss.n298 36.1417
R4894 dvss.n3716 dvss.n298 36.1417
R4895 dvss.n3716 dvss.n3715 36.1417
R4896 dvss.n3715 dvss.n289 36.1417
R4897 dvss.n3728 dvss.n289 36.1417
R4898 dvss.n3728 dvss.n285 36.1417
R4899 dvss.n3745 dvss.n285 36.1417
R4900 dvss.n3745 dvss.n276 36.1417
R4901 dvss.n3760 dvss.n276 36.1417
R4902 dvss.n3760 dvss.n3759 36.1417
R4903 dvss.n3759 dvss.n268 36.1417
R4904 dvss.n3768 dvss.n268 36.1417
R4905 dvss.n3875 dvss.n3768 36.1417
R4906 dvss.n3875 dvss.n3874 36.1417
R4907 dvss.n3874 dvss.n3770 36.1417
R4908 dvss.n3870 dvss.n3770 36.1417
R4909 dvss.n3869 dvss.n3775 36.1417
R4910 dvss.n3782 dvss.n3775 36.1417
R4911 dvss.n3862 dvss.n3782 36.1417
R4912 dvss.n3862 dvss.n3861 36.1417
R4913 dvss.n3861 dvss.n3785 36.1417
R4914 dvss.n3793 dvss.n3785 36.1417
R4915 dvss.n3853 dvss.n3793 36.1417
R4916 dvss.n3853 dvss.n3852 36.1417
R4917 dvss.n3852 dvss.n3796 36.1417
R4918 dvss.n3796 dvss.n127 36.1417
R4919 dvss.n4147 dvss.n127 36.1417
R4920 dvss.n4147 dvss.n4146 36.1417
R4921 dvss.n4146 dvss.n129 36.1417
R4922 dvss.n199 dvss.n129 36.1417
R4923 dvss.n199 dvss.n193 36.1417
R4924 dvss.n210 dvss.n193 36.1417
R4925 dvss.n210 dvss.n140 36.1417
R4926 dvss.n4131 dvss.n140 36.1417
R4927 dvss.n4131 dvss.n4130 36.1417
R4928 dvss.n4130 dvss.n143 36.1417
R4929 dvss.n4126 dvss.n143 36.1417
R4930 dvss.n4125 dvss.n149 36.1417
R4931 dvss.n156 dvss.n149 36.1417
R4932 dvss.n4118 dvss.n156 36.1417
R4933 dvss.n4118 dvss.n4117 36.1417
R4934 dvss.n4117 dvss.n159 36.1417
R4935 dvss.n167 dvss.n159 36.1417
R4936 dvss.n4109 dvss.n167 36.1417
R4937 dvss.n4109 dvss.n4108 36.1417
R4938 dvss.n4108 dvss.n170 36.1417
R4939 dvss.n4097 dvss.n170 36.1417
R4940 dvss.n4097 dvss.n98 36.1417
R4941 dvss.n4194 dvss.n98 36.1417
R4942 dvss.n4194 dvss.n91 36.1417
R4943 dvss.n4211 dvss.n91 36.1417
R4944 dvss.n4211 dvss.n4210 36.1417
R4945 dvss.n4210 dvss.n82 36.1417
R4946 dvss.n82 dvss.n71 36.1417
R4947 dvss.n4231 dvss.n71 36.1417
R4948 dvss.n4232 dvss.n4231 36.1417
R4949 dvss.n4232 dvss.n65 36.1417
R4950 dvss.n4240 dvss.n65 36.1417
R4951 dvss.n2571 dvss.n2114 36.1417
R4952 dvss.n2568 dvss.n2114 36.1417
R4953 dvss.n2568 dvss.n2567 36.1417
R4954 dvss.n2567 dvss.n2117 36.1417
R4955 dvss.n2560 dvss.n2117 36.1417
R4956 dvss.n2560 dvss.n2559 36.1417
R4957 dvss.n2559 dvss.n2122 36.1417
R4958 dvss.n2551 dvss.n2122 36.1417
R4959 dvss.n2551 dvss.n2550 36.1417
R4960 dvss.n2550 dvss.n2128 36.1417
R4961 dvss.n2543 dvss.n2128 36.1417
R4962 dvss.n2543 dvss.n2542 36.1417
R4963 dvss.n2542 dvss.n2132 36.1417
R4964 dvss.n2136 dvss.n2132 36.1417
R4965 dvss.n2533 dvss.n2136 36.1417
R4966 dvss.n2533 dvss.n2532 36.1417
R4967 dvss.n2532 dvss.n2139 36.1417
R4968 dvss.n2528 dvss.n2139 36.1417
R4969 dvss.n2528 dvss.n2527 36.1417
R4970 dvss.n2527 dvss.n2142 36.1417
R4971 dvss.n2523 dvss.n2142 36.1417
R4972 dvss.n976 dvss.n975 35.7652
R4973 dvss.n2012 dvss.t362 35.6569
R4974 dvss.n3166 dvss.t604 35.6569
R4975 dvss.t768 dvss.n4287 35.4058
R4976 dvss.n4287 dvss.t249 35.4058
R4977 dvss.t703 dvss.n96 34.5917
R4978 dvss.n196 dvss.t374 34.5917
R4979 dvss.t403 dvss.n283 34.5917
R4980 dvss.t344 dvss.n345 34.5917
R4981 dvss.t97 dvss.n414 34.5917
R4982 dvss.n1685 dvss.t425 34.5917
R4983 dvss.t275 dvss.n533 34.5917
R4984 dvss.n691 dvss.t394 34.5917
R4985 dvss.t133 dvss.n744 34.5917
R4986 dvss.n4206 dvss 33.9483
R4987 dvss.n4142 dvss 33.9483
R4988 dvss.n3741 dvss 33.9483
R4989 dvss.n3630 dvss 33.9483
R4990 dvss.n3509 dvss 33.9483
R4991 dvss.n1706 dvss 33.9483
R4992 dvss.n1558 dvss 33.9483
R4993 dvss.n712 dvss 33.9483
R4994 dvss.n1171 dvss 33.9483
R4995 dvss.n4022 dvss 33.9483
R4996 dvss.n3943 dvss 33.9483
R4997 dvss.n3260 dvss 33.9483
R4998 dvss.n3310 dvss 33.9483
R4999 dvss.n3365 dvss 33.9483
R5000 dvss.n1812 dvss 33.9483
R5001 dvss.n1416 dvss 33.9483
R5002 dvss.n1329 dvss 33.9483
R5003 dvss.n935 dvss 33.9483
R5004 dvss.n2538 dvss 33.9483
R5005 dvss.n4181 dvss.t623 32.1345
R5006 dvss.t188 dvss.n4154 32.1345
R5007 dvss.n4165 dvss.t53 31.6138
R5008 dvss.t697 dvss.t625 31.1326
R5009 dvss.t382 dvss.t180 31.1326
R5010 dvss.t411 dvss.t366 31.1326
R5011 dvss.t608 dvss.t350 31.1326
R5012 dvss.t95 dvss.t417 31.1326
R5013 dvss.t431 dvss.t45 31.1326
R5014 dvss.t273 dvss.t356 31.1326
R5015 dvss.t392 dvss.t582 31.1326
R5016 dvss.t131 dvss.t197 31.1326
R5017 dvss.n817 dvss.n816 30.6481
R5018 dvss.n867 dvss.n866 30.6481
R5019 dvss.t178 dvss.n121 28.7399
R5020 dvss.t621 dvss.n4186 28.7399
R5021 dvss.n152 dvss.t764 28.1205
R5022 dvss.n3778 dvss.t13 28.1205
R5023 dvss.n3681 dvss.t248 28.1205
R5024 dvss.n3568 dvss.t225 28.1205
R5025 dvss.n3449 dvss.t399 28.1205
R5026 dvss.n1595 dvss.t710 28.1205
R5027 dvss.n1498 dvss.t724 28.1205
R5028 dvss.n1211 dvss.t114 28.1205
R5029 dvss.n1108 dvss.t196 28.1205
R5030 dvss.n30 dvss.t760 28.1205
R5031 dvss.n2035 dvss.t559 28.1205
R5032 dvss.n3204 dvss.t56 28.1205
R5033 dvss.n2874 dvss.t638 28.1205
R5034 dvss.n2835 dvss.t560 28.1205
R5035 dvss.n2796 dvss.t361 28.1205
R5036 dvss.n2757 dvss.t415 28.1205
R5037 dvss.n2718 dvss.t627 28.1205
R5038 dvss.n2679 dvss.t341 28.1205
R5039 dvss.n2186 dvss.t321 28.1205
R5040 dvss.n4093 dvss.n173 27.2737
R5041 dvss.n3839 dvss.n3838 27.2737
R5042 dvss.n3723 dvss.n3722 27.2737
R5043 dvss.n3607 dvss.n3606 27.2737
R5044 dvss.n3491 dvss.n3490 27.2737
R5045 dvss.n1677 dvss.n1638 27.2737
R5046 dvss.n1540 dvss.n1539 27.2737
R5047 dvss.n684 dvss.n683 27.2737
R5048 dvss.n1145 dvss.n1144 27.2737
R5049 dvss.n2216 dvss.t451 26.5065
R5050 dvss.n838 dvss.t47 25.3944
R5051 dvss.n7 dvss.t549 24.9236
R5052 dvss.n7 dvss.t541 24.9236
R5053 dvss.n2 dvss.t597 24.9236
R5054 dvss.n2 dvss.t595 24.9236
R5055 dvss.n2343 dvss.t635 24.9236
R5056 dvss.n2343 dvss.t631 24.9236
R5057 dvss.n2317 dvss.t748 24.9236
R5058 dvss.n2317 dvss.t738 24.9236
R5059 dvss.n2316 dvss.t750 24.9236
R5060 dvss.n2316 dvss.t730 24.9236
R5061 dvss.n2324 dvss.t754 24.9236
R5062 dvss.n2324 dvss.t756 24.9236
R5063 dvss.n2313 dvss.t744 24.9236
R5064 dvss.n2313 dvss.t734 24.9236
R5065 dvss.n2333 dvss.t740 24.9236
R5066 dvss.n2333 dvss.t758 24.9236
R5067 dvss.n2310 dvss.t742 24.9236
R5068 dvss.n2310 dvss.t728 24.9236
R5069 dvss.n2339 dvss.t752 24.9236
R5070 dvss.n2339 dvss.t732 24.9236
R5071 dvss.n2377 dvss.t156 24.9236
R5072 dvss.n2377 dvss.t162 24.9236
R5073 dvss.n2391 dvss.t66 24.9236
R5074 dvss.n2391 dvss.t88 24.9236
R5075 dvss.n2393 dvss.t68 24.9236
R5076 dvss.n2393 dvss.t80 24.9236
R5077 dvss.n2388 dvss.t72 24.9236
R5078 dvss.n2388 dvss.t74 24.9236
R5079 dvss.n2402 dvss.t62 24.9236
R5080 dvss.n2402 dvss.t84 24.9236
R5081 dvss.n2385 dvss.t58 24.9236
R5082 dvss.n2385 dvss.t76 24.9236
R5083 dvss.n2382 dvss.t60 24.9236
R5084 dvss.n2382 dvss.t78 24.9236
R5085 dvss.n2381 dvss.t70 24.9236
R5086 dvss.n2381 dvss.t82 24.9236
R5087 dvss.n2274 dvss.t551 24.9236
R5088 dvss.n2274 dvss.t543 24.9236
R5089 dvss.n2288 dvss.t654 24.9236
R5090 dvss.n2288 dvss.t676 24.9236
R5091 dvss.n2290 dvss.t656 24.9236
R5092 dvss.n2290 dvss.t668 24.9236
R5093 dvss.n2285 dvss.t660 24.9236
R5094 dvss.n2285 dvss.t662 24.9236
R5095 dvss.n2299 dvss.t650 24.9236
R5096 dvss.n2299 dvss.t672 24.9236
R5097 dvss.n2282 dvss.t678 24.9236
R5098 dvss.n2282 dvss.t664 24.9236
R5099 dvss.n2279 dvss.t680 24.9236
R5100 dvss.n2279 dvss.t666 24.9236
R5101 dvss.n2278 dvss.t658 24.9236
R5102 dvss.n2278 dvss.t670 24.9236
R5103 dvss.n2455 dvss.t495 24.9236
R5104 dvss.n2455 dvss.t519 24.9236
R5105 dvss.n2457 dvss.t509 24.9236
R5106 dvss.n2457 dvss.t521 24.9236
R5107 dvss.n2452 dvss.t501 24.9236
R5108 dvss.n2452 dvss.t515 24.9236
R5109 dvss.n2466 dvss.t505 24.9236
R5110 dvss.n2466 dvss.t491 24.9236
R5111 dvss.n2449 dvss.t507 24.9236
R5112 dvss.n2449 dvss.t493 24.9236
R5113 dvss.n2475 dvss.t497 24.9236
R5114 dvss.n2475 dvss.t511 24.9236
R5115 dvss.n2445 dvss.t499 24.9236
R5116 dvss.n2445 dvss.t513 24.9236
R5117 dvss.n823 dvss.n821 22.5639
R5118 dvss.n2660 dvss.n2658 22.5639
R5119 dvss.t457 dvss.n4078 22.5415
R5120 dvss.n3826 dvss.t35 22.5415
R5121 dvss.t2 dvss.n3697 22.5415
R5122 dvss.t237 dvss.n3578 22.5415
R5123 dvss.t210 dvss.n3456 22.5415
R5124 dvss.t331 dvss.n1662 22.5415
R5125 dvss.t222 dvss.n1505 22.5415
R5126 dvss.n1219 dvss.t234 22.5415
R5127 dvss.n777 dvss.t32 22.5415
R5128 dvss.n4301 dvss.n4295 22.2727
R5129 dvss.n1058 dvss.t253 22.0013
R5130 dvss.n880 dvss.t266 22.0013
R5131 dvss.n4206 dvss.n4203 21.8222
R5132 dvss.n4143 dvss.n4142 21.8222
R5133 dvss.n3742 dvss.n3741 21.8222
R5134 dvss.n3631 dvss.n3630 21.8222
R5135 dvss.n3510 dvss.n3509 21.8222
R5136 dvss.n1707 dvss.n1706 21.8222
R5137 dvss.n1559 dvss.n1558 21.8222
R5138 dvss.n713 dvss.n712 21.8222
R5139 dvss.n1172 dvss.n1171 21.8222
R5140 dvss.n4023 dvss.n4022 21.8222
R5141 dvss.n3943 dvss.n3942 21.8222
R5142 dvss.n3261 dvss.n3260 21.8222
R5143 dvss.n3311 dvss.n3310 21.8222
R5144 dvss.n3366 dvss.n3365 21.8222
R5145 dvss.n1812 dvss.n1811 21.8222
R5146 dvss.n1417 dvss.n1416 21.8222
R5147 dvss.n1329 dvss.n1328 21.8222
R5148 dvss.n935 dvss.n931 21.8222
R5149 dvss.n2539 dvss.n2538 21.8222
R5150 dvss.n152 dvss.t601 21.2805
R5151 dvss.n3778 dvss.t446 21.2805
R5152 dvss.n3681 dvss.t767 21.2805
R5153 dvss.n3568 dvss.t192 21.2805
R5154 dvss.n3449 dvss.t694 21.2805
R5155 dvss.n1595 dvss.t692 21.2805
R5156 dvss.n1498 dvss.t590 21.2805
R5157 dvss.n1211 dvss.t629 21.2805
R5158 dvss.n1108 dvss.t194 21.2805
R5159 dvss.n822 dvss.t568 21.2805
R5160 dvss.n822 dvss.t566 21.2805
R5161 dvss.n30 dvss.t54 21.2805
R5162 dvss.n2035 dvss.t571 21.2805
R5163 dvss.n3204 dvss.t722 21.2805
R5164 dvss.n2874 dvss.t236 21.2805
R5165 dvss.n2835 dvss.t569 21.2805
R5166 dvss.n2796 dvss.t177 21.2805
R5167 dvss.n2757 dvss.t339 21.2805
R5168 dvss.n2718 dvss.t176 21.2805
R5169 dvss.n2679 dvss.t340 21.2805
R5170 dvss.n2659 dvss.t122 21.2805
R5171 dvss.n2659 dvss.t121 21.2805
R5172 dvss.n2186 dvss.t696 21.2805
R5173 dvss.n2250 dvss.t530 20.507
R5174 dvss.n1061 dvss.t138 20.3576
R5175 dvss.n2669 dvss.t116 20.3576
R5176 dvss.n4204 dvss.t626 20.0005
R5177 dvss.n4204 dvss.t323 20.0005
R5178 dvss.n132 dvss.t181 20.0005
R5179 dvss.n132 dvss.t1 20.0005
R5180 dvss.n3739 dvss.t367 20.0005
R5181 dvss.n3739 dvss.t164 20.0005
R5182 dvss.n3628 dvss.t609 20.0005
R5183 dvss.n3628 dvss.t338 20.0005
R5184 dvss.n3507 dvss.t418 20.0005
R5185 dvss.n3507 dvss.t316 20.0005
R5186 dvss.n1629 dvss.t46 20.0005
R5187 dvss.n1629 dvss.t319 20.0005
R5188 dvss.n1556 dvss.t357 20.0005
R5189 dvss.n1556 dvss.t304 20.0005
R5190 dvss.n674 dvss.t583 20.0005
R5191 dvss.n674 dvss.t301 20.0005
R5192 dvss.n1169 dvss.t198 20.0005
R5193 dvss.n1169 dvss.t402 20.0005
R5194 dvss.n3995 dvss.t708 20.0005
R5195 dvss.n3995 dvss.t539 20.0005
R5196 dvss.n226 dvss.t377 20.0005
R5197 dvss.n226 dvss.t140 20.0005
R5198 dvss.n1915 dvss.t408 20.0005
R5199 dvss.n1915 dvss.t762 20.0005
R5200 dvss.n1884 dvss.t349 20.0005
R5201 dvss.n1884 dvss.t152 20.0005
R5202 dvss.n1853 dvss.t92 20.0005
R5203 dvss.n1853 dvss.t307 20.0005
R5204 dvss.n472 dvss.t424 20.0005
R5205 dvss.n472 dvss.t310 20.0005
R5206 dvss.n1370 dvss.t272 20.0005
R5207 dvss.n1370 dvss.t292 20.0005
R5208 dvss.n592 dvss.t387 20.0005
R5209 dvss.n592 dvss.t289 20.0005
R5210 dvss.n932 dvss.t126 20.0005
R5211 dvss.n932 dvss.t336 20.0005
R5212 dvss.n2134 dvss.t525 20.0005
R5213 dvss.n2134 dvss.t553 20.0005
R5214 dvss.n4269 dvss.t591 19.2955
R5215 dvss.t455 dvss.n2209 18.9334
R5216 dvss.n180 dvss.n179 18.8324
R5217 dvss.n3818 dvss.n3817 18.8324
R5218 dvss.n324 dvss.n314 18.8324
R5219 dvss.n3548 dvss.n382 18.8324
R5220 dvss.n3442 dvss.n443 18.8324
R5221 dvss.n1645 dvss.n1644 18.8324
R5222 dvss.n1491 dvss.n562 18.8324
R5223 dvss.n1257 dvss.n637 18.8324
R5224 dvss.n979 dvss.t561 18.6559
R5225 dvss.n800 dvss.n776 18.6144
R5226 dvss.n3986 dvss.t685 18.3666
R5227 dvss.n3922 dvss.t147 18.3666
R5228 dvss.n3239 dvss.t473 18.3666
R5229 dvss.n1972 dvss.t20 18.3666
R5230 dvss.n1947 dvss.t482 18.3666
R5231 dvss.n1791 dvss.t443 18.3666
R5232 dvss.n1390 dvss.t101 18.3666
R5233 dvss.n1308 dvss.t719 18.3666
R5234 dvss.n955 dvss.t647 18.3666
R5235 dvss.n2516 dvss 18.0711
R5236 dvss.n3112 dvss 18.0711
R5237 dvss.n3109 dvss 18.0711
R5238 dvss.n3068 dvss 18.0711
R5239 dvss.n3065 dvss 18.0711
R5240 dvss.n3024 dvss 18.0711
R5241 dvss.n3021 dvss 18.0711
R5242 dvss.n2980 dvss 18.0711
R5243 dvss.n2977 dvss 18.0711
R5244 dvss.n2936 dvss 18.0711
R5245 dvss.n2933 dvss 18.0711
R5246 dvss.n2892 dvss 18.0711
R5247 dvss.n2889 dvss 18.0711
R5248 dvss.n3194 dvss 18.0711
R5249 dvss dvss.n2087 18.0711
R5250 dvss.n2066 dvss 18.0711
R5251 dvss dvss.n2065 18.0711
R5252 dvss.n4361 dvss 18.0711
R5253 dvss dvss.n4360 18.0711
R5254 dvss.n4314 dvss 18.0711
R5255 dvss.n789 dvss 18.0711
R5256 dvss.n1206 dvss 18.0711
R5257 dvss dvss.n723 18.0711
R5258 dvss.n1484 dvss 18.0711
R5259 dvss dvss.n560 18.0711
R5260 dvss.n1739 dvss 18.0711
R5261 dvss dvss.n1738 18.0711
R5262 dvss.n3425 dvss 18.0711
R5263 dvss dvss.n441 18.0711
R5264 dvss.n3556 dvss 18.0711
R5265 dvss.n3553 dvss 18.0711
R5266 dvss.n318 dvss 18.0711
R5267 dvss dvss.n312 18.0711
R5268 dvss.n3870 dvss 18.0711
R5269 dvss dvss.n3869 18.0711
R5270 dvss.n4126 dvss 18.0711
R5271 dvss dvss.n4125 18.0711
R5272 dvss.n4240 dvss 18.0711
R5273 dvss.n4258 dvss.t313 18.0005
R5274 dvss dvss.n779 17.6946
R5275 dvss.n4252 dvss.t535 17.4005
R5276 dvss.n4252 dvss.t283 17.4005
R5277 dvss.n4251 dvss.t112 17.4005
R5278 dvss.n4251 dvss.t286 17.4005
R5279 dvss.n4250 dvss.t537 17.4005
R5280 dvss.n4250 dvss.t575 17.4005
R5281 dvss.n4258 dvss.t580 17.4005
R5282 dvss.n4245 dvss.t295 17.4005
R5283 dvss.n4245 dvss.t479 17.4005
R5284 dvss.n2371 dvss.t280 17.4005
R5285 dvss.n2371 dvss.t298 17.4005
R5286 dvss.n2373 dvss.t158 17.4005
R5287 dvss.n2373 dvss.t168 17.4005
R5288 dvss.n4153 dvss.n103 17.2441
R5289 dvss.n4280 dvss.n4279 17.1002
R5290 dvss.n4281 dvss.n4280 16.9365
R5291 dvss.n2247 dvss.t526 16.8072
R5292 dvss.n1345 dvss.n1344 16.666
R5293 dvss.n1828 dvss.n1827 16.6189
R5294 dvss.n1408 dvss.n1407 16.6189
R5295 dvss.n458 dvss.n457 16.615
R5296 dvss.n578 dvss.n577 16.615
R5297 dvss.n400 dvss.n399 16.611
R5298 dvss.n519 dvss.n518 16.6032
R5299 dvss.n3357 dvss.n3356 16.5915
R5300 dvss.n4272 dvss.n4243 16.3843
R5301 dvss.n2326 dvss.n2323 16.3561
R5302 dvss.n2330 dvss.n2314 16.3561
R5303 dvss.n2335 dvss.n2332 16.3561
R5304 dvss.n2357 dvss.n2356 16.3561
R5305 dvss.n2353 dvss.n2352 16.3561
R5306 dvss.n2349 dvss.n2348 16.3561
R5307 dvss.n2348 dvss.n2347 16.3561
R5308 dvss.n2296 dvss.n2286 16.3561
R5309 dvss.n2301 dvss.n2298 16.3561
R5310 dvss.n2305 dvss.n2283 16.3561
R5311 dvss.n2500 dvss.n2499 16.3561
R5312 dvss.n2505 dvss.n2503 16.3561
R5313 dvss.n2509 dvss.n2275 16.3561
R5314 dvss.n2510 dvss.n2509 16.3561
R5315 dvss.n1242 dvss.n656 16.2675
R5316 dvss.n4090 dvss.n4089 16.2668
R5317 dvss.n3837 dvss.n3802 16.2668
R5318 dvss.n3721 dvss.n293 16.2668
R5319 dvss.n3605 dvss.n360 16.2668
R5320 dvss.n3489 dvss.n3488 16.2668
R5321 dvss.n1674 dvss.n1673 16.2668
R5322 dvss.n1538 dvss.n1537 16.2668
R5323 dvss.n1148 dvss.n759 16.2668
R5324 dvss.n2321 dvss.n2318 16.1783
R5325 dvss.n2292 dvss.n2289 16.1783
R5326 dvss.n2399 dvss.n2389 16.132
R5327 dvss.n2404 dvss.n2401 16.132
R5328 dvss.n2408 dvss.n2386 16.132
R5329 dvss.n2419 dvss.n2418 16.132
R5330 dvss.n2424 dvss.n2422 16.132
R5331 dvss.n2428 dvss.n2378 16.132
R5332 dvss.n2429 dvss.n2428 16.132
R5333 dvss.n994 dvss.t725 15.9908
R5334 dvss.n2395 dvss.n2392 15.9567
R5335 dvss.n2359 dvss.n2358 15.8227
R5336 dvss.n2498 dvss.n2497 15.8227
R5337 dvss.n2363 dvss.n2362 15.6449
R5338 dvss.n2494 dvss.n2493 15.6449
R5339 dvss.n2417 dvss.n2416 15.606
R5340 dvss.n2347 dvss.n2344 15.2894
R5341 dvss.n2511 dvss.n2510 15.2894
R5342 dvss.n2430 dvss.n2429 15.08
R5343 dvss.n2349 dvss.n2341 14.9338
R5344 dvss.n2504 dvss.n2275 14.9338
R5345 dvss.n2423 dvss.n2378 14.7293
R5346 dvss.n2463 dvss.n2453 14.7205
R5347 dvss.n2468 dvss.n2465 14.7205
R5348 dvss.n2472 dvss.n2450 14.7205
R5349 dvss.n2477 dvss.n2474 14.7205
R5350 dvss.n2483 dvss.n2447 14.7205
R5351 dvss.n4406 dvss.n1 14.7205
R5352 dvss.n4404 dvss.n4403 14.7205
R5353 dvss.n4403 dvss.n3 14.7205
R5354 dvss.n4399 dvss.n4398 14.7205
R5355 dvss.n4395 dvss.n4394 14.7205
R5356 dvss.n4394 dvss.n4393 14.7205
R5357 dvss.n3143 dvss.n2575 14.5906
R5358 dvss.n2459 dvss.n2456 14.5605
R5359 dvss.n2413 dvss.n2412 14.5539
R5360 dvss.n838 dvss.t117 14.1215
R5361 dvss.n2359 dvss.n2311 14.0449
R5362 dvss.n2356 dvss.n2340 14.0449
R5363 dvss.n2497 dvss.n2280 14.0449
R5364 dvss.n2500 dvss.n2276 14.0449
R5365 dvss.n2416 dvss.n2383 13.8526
R5366 dvss.n2419 dvss.n2379 13.8526
R5367 dvss.n4 dvss.n3 13.7605
R5368 dvss.n2322 dvss.n2321 13.6894
R5369 dvss.n2292 dvss.n2291 13.6894
R5370 dvss.n2395 dvss.n2394 13.5019
R5371 dvss.n4405 dvss.n4404 13.4405
R5372 dvss.n4395 dvss.n5 13.4405
R5373 dvss.n4278 dvss.n4272 13.3982
R5374 dvss.n4393 dvss.n8 13.2077
R5375 dvss.n3979 dvss.t689 13.1192
R5376 dvss.t141 dvss.n3905 13.1192
R5377 dvss.t467 dvss.n1991 13.1192
R5378 dvss.t14 dvss.n1966 13.1192
R5379 dvss.n1938 dvss.t486 13.1192
R5380 dvss.t441 dvss.n1774 13.1192
R5381 dvss.n1381 dvss.t107 13.1192
R5382 dvss.t715 dvss.n1291 13.1192
R5383 dvss.n970 dvss.t645 13.1192
R5384 dvss.n4278 dvss.n4277 13.0828
R5385 dvss.n2476 dvss.n2444 12.6405
R5386 dvss.n2447 dvss.n2446 12.6405
R5387 dvss.n4207 dvss.n4206 12.5222
R5388 dvss.n4142 dvss.n131 12.5222
R5389 dvss.n3741 dvss.n3738 12.5222
R5390 dvss.n3630 dvss.n3627 12.5222
R5391 dvss.n3509 dvss.n3506 12.5222
R5392 dvss.n1706 dvss.n1628 12.5222
R5393 dvss.n1558 dvss.n1555 12.5222
R5394 dvss.n712 dvss.n673 12.5222
R5395 dvss.n1171 dvss.n1168 12.5222
R5396 dvss.n4022 dvss.n3994 12.5222
R5397 dvss.n3943 dvss.n229 12.5222
R5398 dvss.n3260 dvss.n1914 12.5222
R5399 dvss.n3310 dvss.n1883 12.5222
R5400 dvss.n3365 dvss.n1852 12.5222
R5401 dvss.n1812 dvss.n475 12.5222
R5402 dvss.n1416 dvss.n1369 12.5222
R5403 dvss.n1329 dvss.n595 12.5222
R5404 dvss.n936 dvss.n935 12.5222
R5405 dvss.n2538 dvss.n2133 12.5222
R5406 dvss.n2459 dvss.n2458 12.3205
R5407 dvss.n824 dvss.n823 12.2361
R5408 dvss.n2661 dvss.n2660 12.2361
R5409 dvss.n818 dvss.n817 12.1422
R5410 dvss.n869 dvss.n867 12.1422
R5411 dvss.t228 dvss.n656 11.3665
R5412 dvss.n4089 dvss.t463 11.3663
R5413 dvss.n3837 dvss.t41 11.3663
R5414 dvss.n3721 dvss.t8 11.3663
R5415 dvss.n3605 dvss.t243 11.3663
R5416 dvss.n3489 dvss.t206 11.3663
R5417 dvss.n1673 dvss.t333 11.3663
R5418 dvss.n1538 dvss.t216 11.3663
R5419 dvss.t24 dvss.n759 11.3663
R5420 dvss.n2334 dvss.n2309 11.2005
R5421 dvss.n2307 dvss.n2306 11.2005
R5422 dvss.n2410 dvss.n2409 11.0471
R5423 dvss.n2326 dvss.n2325 10.8449
R5424 dvss.n2297 dvss.n2296 10.8449
R5425 dvss.n4391 dvss.n8 10.7826
R5426 dvss.n2400 dvss.n2399 10.6964
R5427 dvss.n164 dvss.t462 10.6405
R5428 dvss.n164 dvss.t464 10.6405
R5429 dvss.n162 dvss.t458 10.6405
R5430 dvss.n162 dvss.t460 10.6405
R5431 dvss.n3790 dvss.t40 10.6405
R5432 dvss.n3790 dvss.t42 10.6405
R5433 dvss.n3788 dvss.t36 10.6405
R5434 dvss.n3788 dvss.t38 10.6405
R5435 dvss.n3708 dvss.t7 10.6405
R5436 dvss.n3708 dvss.t9 10.6405
R5437 dvss.n3688 dvss.t3 10.6405
R5438 dvss.n3688 dvss.t5 10.6405
R5439 dvss.n3590 dvss.t242 10.6405
R5440 dvss.n3590 dvss.t244 10.6405
R5441 dvss.n367 dvss.t238 10.6405
R5442 dvss.n367 dvss.t240 10.6405
R5443 dvss.n3476 dvss.t209 10.6405
R5444 dvss.n3476 dvss.t207 10.6405
R5445 dvss.n3462 dvss.t211 10.6405
R5446 dvss.n3462 dvss.t213 10.6405
R5447 dvss.n1607 dvss.t328 10.6405
R5448 dvss.n1607 dvss.t334 10.6405
R5449 dvss.n1605 dvss.t332 10.6405
R5450 dvss.n1605 dvss.t330 10.6405
R5451 dvss.n1525 dvss.t219 10.6405
R5452 dvss.n1525 dvss.t217 10.6405
R5453 dvss.n1511 dvss.t223 10.6405
R5454 dvss.n1511 dvss.t221 10.6405
R5455 dvss.n1231 dvss.t233 10.6405
R5456 dvss.n1231 dvss.t229 10.6405
R5457 dvss.n721 dvss.t235 10.6405
R5458 dvss.n721 dvss.t231 10.6405
R5459 dvss.n754 dvss.t31 10.6405
R5460 dvss.n754 dvss.t25 10.6405
R5461 dvss.n767 dvss.t33 10.6405
R5462 dvss.n767 dvss.t27 10.6405
R5463 dvss.n85 dvss.t700 10.6405
R5464 dvss.n85 dvss.t704 10.6405
R5465 dvss.n88 dvss.t698 10.6405
R5466 dvss.n88 dvss.t706 10.6405
R5467 dvss.n136 dvss.t379 10.6405
R5468 dvss.n136 dvss.t375 10.6405
R5469 dvss.n4136 dvss.t383 10.6405
R5470 dvss.n4136 dvss.t385 10.6405
R5471 dvss.n270 dvss.t410 10.6405
R5472 dvss.n270 dvss.t404 10.6405
R5473 dvss.n273 dvss.t412 10.6405
R5474 dvss.n273 dvss.t406 10.6405
R5475 dvss.n333 dvss.t343 10.6405
R5476 dvss.n333 dvss.t345 10.6405
R5477 dvss.n336 dvss.t351 10.6405
R5478 dvss.n336 dvss.t347 10.6405
R5479 dvss.n401 dvss.t100 10.6405
R5480 dvss.n401 dvss.t98 10.6405
R5481 dvss.n404 dvss.t96 10.6405
R5482 dvss.n404 dvss.t94 10.6405
R5483 dvss.n1623 dvss.t434 10.6405
R5484 dvss.n1623 dvss.t426 10.6405
R5485 dvss.n1700 dvss.t432 10.6405
R5486 dvss.n1700 dvss.t430 10.6405
R5487 dvss.n520 dvss.t278 10.6405
R5488 dvss.n520 dvss.t276 10.6405
R5489 dvss.n523 dvss.t274 10.6405
R5490 dvss.n523 dvss.t268 10.6405
R5491 dvss.n668 dvss.t397 10.6405
R5492 dvss.n668 dvss.t395 10.6405
R5493 dvss.n706 dvss.t393 10.6405
R5494 dvss.n706 dvss.t391 10.6405
R5495 dvss.n731 dvss.t136 10.6405
R5496 dvss.n731 dvss.t134 10.6405
R5497 dvss.n734 dvss.t132 10.6405
R5498 dvss.n734 dvss.t130 10.6405
R5499 dvss.n3969 dvss.t684 10.6405
R5500 dvss.n3969 dvss.t686 10.6405
R5501 dvss.n3962 dvss.t690 10.6405
R5502 dvss.n3962 dvss.t682 10.6405
R5503 dvss.n236 dvss.t146 10.6405
R5504 dvss.n236 dvss.t148 10.6405
R5505 dvss.n245 dvss.t142 10.6405
R5506 dvss.n245 dvss.t144 10.6405
R5507 dvss.n1905 dvss.t472 10.6405
R5508 dvss.n1905 dvss.t474 10.6405
R5509 dvss.n1899 dvss.t468 10.6405
R5510 dvss.n1899 dvss.t470 10.6405
R5511 dvss.n1874 dvss.t19 10.6405
R5512 dvss.n1874 dvss.t21 10.6405
R5513 dvss.n1868 dvss.t15 10.6405
R5514 dvss.n1868 dvss.t17 10.6405
R5515 dvss.n1843 dvss.t485 10.6405
R5516 dvss.n1843 dvss.t483 10.6405
R5517 dvss.n1836 dvss.t487 10.6405
R5518 dvss.n1836 dvss.t489 10.6405
R5519 dvss.n482 dvss.t438 10.6405
R5520 dvss.n482 dvss.t444 10.6405
R5521 dvss.n491 dvss.t442 10.6405
R5522 dvss.n491 dvss.t440 10.6405
R5523 dvss.n1360 dvss.t104 10.6405
R5524 dvss.n1360 dvss.t102 10.6405
R5525 dvss.n1353 dvss.t108 10.6405
R5526 dvss.n1353 dvss.t106 10.6405
R5527 dvss.n602 dvss.t714 10.6405
R5528 dvss.n602 dvss.t720 10.6405
R5529 dvss.n611 dvss.t716 10.6405
R5530 dvss.n611 dvss.t712 10.6405
R5531 dvss.n916 dvss.t644 10.6405
R5532 dvss.n916 dvss.t648 10.6405
R5533 dvss.n908 dvss.t646 10.6405
R5534 dvss.n908 dvss.t640 10.6405
R5535 dvss.n4338 dvss.t618 10.6405
R5536 dvss.n4338 dvss.t622 10.6405
R5537 dvss.n4330 dvss.t616 10.6405
R5538 dvss.n4330 dvss.t624 10.6405
R5539 dvss.n4371 dvss.t183 10.6405
R5540 dvss.n4371 dvss.t179 10.6405
R5541 dvss.n20 dvss.t187 10.6405
R5542 dvss.n20 dvss.t189 10.6405
R5543 dvss.n2076 dvss.t369 10.6405
R5544 dvss.n2076 dvss.t363 10.6405
R5545 dvss.n2002 dvss.t371 10.6405
R5546 dvss.n2002 dvss.t365 10.6405
R5547 dvss.n2096 dvss.t603 10.6405
R5548 dvss.n2096 dvss.t605 10.6405
R5549 dvss.n2099 dvss.t611 10.6405
R5550 dvss.n2099 dvss.t607 10.6405
R5551 dvss.n2855 dvss.t422 10.6405
R5552 dvss.n2855 dvss.t421 10.6405
R5553 dvss.n2859 dvss.t420 10.6405
R5554 dvss.n2859 dvss.t419 10.6405
R5555 dvss.n2816 dvss.t52 10.6405
R5556 dvss.n2816 dvss.t48 10.6405
R5557 dvss.n2820 dvss.t51 10.6405
R5558 dvss.n2820 dvss.t50 10.6405
R5559 dvss.n2777 dvss.t360 10.6405
R5560 dvss.n2777 dvss.t359 10.6405
R5561 dvss.n2781 dvss.t358 10.6405
R5562 dvss.n2781 dvss.t354 10.6405
R5563 dvss.n2738 dvss.t588 10.6405
R5564 dvss.n2738 dvss.t587 10.6405
R5565 dvss.n2742 dvss.t586 10.6405
R5566 dvss.n2742 dvss.t585 10.6405
R5567 dvss.n2699 dvss.t203 10.6405
R5568 dvss.n2699 dvss.t202 10.6405
R5569 dvss.n2703 dvss.t201 10.6405
R5570 dvss.n2703 dvss.t200 10.6405
R5571 dvss.n2152 dvss.t533 10.6405
R5572 dvss.n2152 dvss.t527 10.6405
R5573 dvss.n2155 dvss.t529 10.6405
R5574 dvss.n2155 dvss.t531 10.6405
R5575 dvss.n2124 dvss.t450 10.6405
R5576 dvss.n2124 dvss.t452 10.6405
R5577 dvss.n2118 dvss.t456 10.6405
R5578 dvss.n2118 dvss.t448 10.6405
R5579 dvss.n163 dvss.n161 10.64
R5580 dvss.n3789 dvss.n3787 10.64
R5581 dvss.n3693 dvss.n3692 10.64
R5582 dvss.n376 dvss.n368 10.64
R5583 dvss.n3463 dvss.n3461 10.64
R5584 dvss.n1606 dvss.n1604 10.64
R5585 dvss.n1512 dvss.n1510 10.64
R5586 dvss.n722 dvss.n720 10.64
R5587 dvss.n1122 dvss.n768 10.64
R5588 dvss.n4049 dvss.n4048 10.64
R5589 dvss.n3899 dvss.n246 10.64
R5590 dvss.n3287 dvss.n3286 10.64
R5591 dvss.n3337 dvss.n3336 10.64
R5592 dvss.n3392 dvss.n3391 10.64
R5593 dvss.n1768 dvss.n492 10.64
R5594 dvss.n1443 dvss.n1442 10.64
R5595 dvss.n1285 dvss.n612 10.64
R5596 dvss.n909 dvss.n907 10.64
R5597 dvss.n2565 dvss.n2564 10.64
R5598 dvss.n4283 dvss.n4265 10.6369
R5599 dvss.n4287 dvss.n4265 10.6369
R5600 dvss.n4286 dvss.n4285 10.6369
R5601 dvss.n4287 dvss.n4286 10.6369
R5602 dvss.n4263 dvss.n4262 10.6369
R5603 dvss.n4266 dvss.n4263 10.6369
R5604 dvss.n4292 dvss.n4249 10.6369
R5605 dvss.n4266 dvss.n4249 10.6369
R5606 dvss.t175 dvss.t119 10.555
R5607 dvss.n2345 dvss.n2344 10.3672
R5608 dvss.n2512 dvss.n2511 10.3672
R5609 dvss.n2431 dvss.n2430 10.3526
R5610 dvss.t119 dvss.t115 10.2446
R5611 dvss.n2474 dvss.n2473 10.0805
R5612 dvss.n2486 dvss.t498 10.0615
R5613 dvss.n2464 dvss.n2463 9.7605
R5614 dvss.n3141 dvss 9.31486
R5615 dvss.n2175 dvss 9.31486
R5616 dvss.n2571 dvss 9.31486
R5617 dvss.n1009 dvss 9.30735
R5618 dvss.n1020 dvss.n835 9.30085
R5619 dvss.n825 dvss.n824 9.3005
R5620 dvss.n824 dvss.n820 9.3005
R5621 dvss.n1064 dvss.n1063 9.3005
R5622 dvss.n1063 dvss.n1057 9.3005
R5623 dvss.n1111 dvss.n1110 9.3005
R5624 dvss.n1112 dvss.n1111 9.3005
R5625 dvss.n1196 dvss.n1195 9.3005
R5626 dvss.n1197 dvss.n1196 9.3005
R5627 dvss.n1193 dvss.n733 9.3005
R5628 dvss.n1193 dvss.n1192 9.3005
R5629 dvss.n748 dvss.n732 9.3005
R5630 dvss.n1157 dvss.n732 9.3005
R5631 dvss.n1214 dvss.n1213 9.3005
R5632 dvss.n1215 dvss.n1214 9.3005
R5633 dvss.n1467 dvss.n1466 9.3005
R5634 dvss.n1466 dvss.n1465 9.3005
R5635 dvss.n709 dvss.n708 9.3005
R5636 dvss.n708 dvss.n707 9.3005
R5637 dvss.n670 dvss.n669 9.3005
R5638 dvss.n669 dvss.n663 9.3005
R5639 dvss.n1501 dvss.n1500 9.3005
R5640 dvss.n1500 dvss.n1497 9.3005
R5641 dvss.n1582 dvss.n512 9.3005
R5642 dvss.n1583 dvss.n1582 9.3005
R5643 dvss.n1580 dvss.n522 9.3005
R5644 dvss.n1580 dvss.n1579 9.3005
R5645 dvss.n1550 dvss.n521 9.3005
R5646 dvss.n538 dvss.n521 9.3005
R5647 dvss.n1734 dvss.n1733 9.3005
R5648 dvss.n1735 dvss.n1734 9.3005
R5649 dvss.n3416 dvss.n3415 9.3005
R5650 dvss.n3415 dvss.n3414 9.3005
R5651 dvss.n1703 dvss.n1702 9.3005
R5652 dvss.n1702 dvss.n1701 9.3005
R5653 dvss.n1625 dvss.n1624 9.3005
R5654 dvss.n1624 dvss.n1617 9.3005
R5655 dvss.n3452 dvss.n3451 9.3005
R5656 dvss.n3451 dvss.n3448 9.3005
R5657 dvss.n3534 dvss.n392 9.3005
R5658 dvss.n3535 dvss.n3534 9.3005
R5659 dvss.n3532 dvss.n403 9.3005
R5660 dvss.n3532 dvss.n3531 9.3005
R5661 dvss.n3501 dvss.n402 9.3005
R5662 dvss.n419 dvss.n402 9.3005
R5663 dvss.n3571 dvss.n3570 9.3005
R5664 dvss.n3570 dvss.n3567 9.3005
R5665 dvss.n3651 dvss.n330 9.3005
R5666 dvss.n3652 dvss.n3651 9.3005
R5667 dvss.n3649 dvss.n335 9.3005
R5668 dvss.n3649 dvss.n3648 9.3005
R5669 dvss.n3617 dvss.n334 9.3005
R5670 dvss.n354 dvss.n334 9.3005
R5671 dvss.n3684 dvss.n3683 9.3005
R5672 dvss.n3683 dvss.n3680 9.3005
R5673 dvss.n3765 dvss.n267 9.3005
R5674 dvss.n3766 dvss.n3765 9.3005
R5675 dvss.n3763 dvss.n272 9.3005
R5676 dvss.n3763 dvss.n3762 9.3005
R5677 dvss.n3733 dvss.n271 9.3005
R5678 dvss.n288 dvss.n271 9.3005
R5679 dvss.n3865 dvss.n3864 9.3005
R5680 dvss.n3866 dvss.n3865 9.3005
R5681 dvss.n4134 dvss.n4133 9.3005
R5682 dvss.n4134 dvss.n138 9.3005
R5683 dvss.n4139 dvss.n4138 9.3005
R5684 dvss.n4138 dvss.n4137 9.3005
R5685 dvss.n137 dvss.n135 9.3005
R5686 dvss.n3843 dvss.n137 9.3005
R5687 dvss.n4121 dvss.n4120 9.3005
R5688 dvss.n4122 dvss.n4121 9.3005
R5689 dvss.n4216 dvss.n73 9.3005
R5690 dvss.n4217 dvss.n4216 9.3005
R5691 dvss.n4214 dvss.n87 9.3005
R5692 dvss.n4214 dvss.n4213 9.3005
R5693 dvss.n4192 dvss.n86 9.3005
R5694 dvss.n4099 dvss.n86 9.3005
R5695 dvss.n1031 dvss.n1030 9.3005
R5696 dvss.n1030 dvss.n1029 9.3005
R5697 dvss.n1066 dvss.n1065 9.3005
R5698 dvss.n1067 dvss.n1066 9.3005
R5699 dvss.n1170 dvss.n736 9.3005
R5700 dvss.n1168 dvss.n1167 9.3005
R5701 dvss.n1155 dvss.n753 9.3005
R5702 dvss.n1132 dvss.n1131 9.3005
R5703 dvss.n1135 dvss.n1134 9.3005
R5704 dvss.n1153 dvss.n1152 9.3005
R5705 dvss.n1156 dvss.n1155 9.3005
R5706 dvss.n711 dvss.n710 9.3005
R5707 dvss.n705 dvss.n673 9.3005
R5708 dvss.n1237 dvss.n1236 9.3005
R5709 dvss.n1227 dvss.n1226 9.3005
R5710 dvss.n1230 dvss.n1229 9.3005
R5711 dvss.n1234 dvss.n1233 9.3005
R5712 dvss.n1236 dvss.n719 9.3005
R5713 dvss.n1557 dvss.n525 9.3005
R5714 dvss.n1555 dvss.n1554 9.3005
R5715 dvss.n1548 dvss.n1547 9.3005
R5716 dvss.n1514 dvss.n1513 9.3005
R5717 dvss.n1524 dvss.n1523 9.3005
R5718 dvss.n1529 dvss.n1528 9.3005
R5719 dvss.n1549 dvss.n1548 9.3005
R5720 dvss.n1705 dvss.n1704 9.3005
R5721 dvss.n1699 dvss.n1628 9.3005
R5722 dvss.n1718 dvss.n1717 9.3005
R5723 dvss.n1728 dvss.n1727 9.3005
R5724 dvss.n1725 dvss.n1724 9.3005
R5725 dvss.n1715 dvss.n1714 9.3005
R5726 dvss.n1717 dvss.n1713 9.3005
R5727 dvss.n3508 dvss.n406 9.3005
R5728 dvss.n3506 dvss.n3505 9.3005
R5729 dvss.n3499 dvss.n3498 9.3005
R5730 dvss.n3465 dvss.n3464 9.3005
R5731 dvss.n3475 dvss.n3474 9.3005
R5732 dvss.n3480 dvss.n3479 9.3005
R5733 dvss.n3500 dvss.n3499 9.3005
R5734 dvss.n3629 dvss.n338 9.3005
R5735 dvss.n3627 dvss.n3626 9.3005
R5736 dvss.n3615 dvss.n3614 9.3005
R5737 dvss.n3588 dvss.n3587 9.3005
R5738 dvss.n3597 dvss.n3596 9.3005
R5739 dvss.n3594 dvss.n3593 9.3005
R5740 dvss.n3616 dvss.n3615 9.3005
R5741 dvss.n3740 dvss.n275 9.3005
R5742 dvss.n3738 dvss.n3737 9.3005
R5743 dvss.n3731 dvss.n3730 9.3005
R5744 dvss.n3691 dvss.n3690 9.3005
R5745 dvss.n3707 dvss.n3706 9.3005
R5746 dvss.n3712 dvss.n3711 9.3005
R5747 dvss.n3732 dvss.n3731 9.3005
R5748 dvss.n4141 dvss.n4140 9.3005
R5749 dvss.n134 dvss.n131 9.3005
R5750 dvss.n3849 dvss.n3848 9.3005
R5751 dvss.n3859 dvss.n3858 9.3005
R5752 dvss.n3856 dvss.n3855 9.3005
R5753 dvss.n3846 dvss.n3845 9.3005
R5754 dvss.n3848 dvss.n3844 9.3005
R5755 dvss.n4205 dvss.n90 9.3005
R5756 dvss.n4208 dvss.n4207 9.3005
R5757 dvss.n4105 dvss.n4104 9.3005
R5758 dvss.n4115 dvss.n4114 9.3005
R5759 dvss.n4112 dvss.n4111 9.3005
R5760 dvss.n4102 dvss.n4101 9.3005
R5761 dvss.n4104 dvss.n4100 9.3005
R5762 dvss.n818 dvss.n815 9.3005
R5763 dvss.n819 dvss.n818 9.3005
R5764 dvss.n858 dvss.n857 9.3005
R5765 dvss.n857 dvss.n856 9.3005
R5766 dvss.n883 dvss.n882 9.3005
R5767 dvss.n882 dvss.n881 9.3005
R5768 dvss.n934 dvss.n933 9.3005
R5769 dvss.n937 dvss.n936 9.3005
R5770 dvss.n923 dvss.n922 9.3005
R5771 dvss.n911 dvss.n910 9.3005
R5772 dvss.n915 dvss.n914 9.3005
R5773 dvss.n919 dvss.n918 9.3005
R5774 dvss.n924 dvss.n923 9.3005
R5775 dvss.n1331 dvss.n1330 9.3005
R5776 dvss.n595 dvss.n594 9.3005
R5777 dvss.n1315 dvss.n600 9.3005
R5778 dvss.n1298 dvss.n1297 9.3005
R5779 dvss.n1301 dvss.n1300 9.3005
R5780 dvss.n1313 dvss.n1312 9.3005
R5781 dvss.n1316 dvss.n1315 9.3005
R5782 dvss.n1415 dvss.n1414 9.3005
R5783 dvss.n1413 dvss.n1369 9.3005
R5784 dvss.n1426 dvss.n1425 9.3005
R5785 dvss.n1441 dvss.n1440 9.3005
R5786 dvss.n1435 dvss.n1434 9.3005
R5787 dvss.n1432 dvss.n1431 9.3005
R5788 dvss.n1425 dvss.n1423 9.3005
R5789 dvss.n1814 dvss.n1813 9.3005
R5790 dvss.n475 dvss.n474 9.3005
R5791 dvss.n1798 dvss.n480 9.3005
R5792 dvss.n1781 dvss.n1780 9.3005
R5793 dvss.n1784 dvss.n1783 9.3005
R5794 dvss.n1796 dvss.n1795 9.3005
R5795 dvss.n1799 dvss.n1798 9.3005
R5796 dvss.n3364 dvss.n3363 9.3005
R5797 dvss.n3362 dvss.n1852 9.3005
R5798 dvss.n3375 dvss.n3374 9.3005
R5799 dvss.n3390 dvss.n3389 9.3005
R5800 dvss.n3384 dvss.n3383 9.3005
R5801 dvss.n3381 dvss.n3380 9.3005
R5802 dvss.n3374 dvss.n3372 9.3005
R5803 dvss.n3309 dvss.n3308 9.3005
R5804 dvss.n3307 dvss.n1883 9.3005
R5805 dvss.n3320 dvss.n3319 9.3005
R5806 dvss.n3335 dvss.n3334 9.3005
R5807 dvss.n3329 dvss.n3328 9.3005
R5808 dvss.n3326 dvss.n3325 9.3005
R5809 dvss.n3319 dvss.n3317 9.3005
R5810 dvss.n3259 dvss.n3258 9.3005
R5811 dvss.n3257 dvss.n1914 9.3005
R5812 dvss.n3270 dvss.n3269 9.3005
R5813 dvss.n3285 dvss.n3284 9.3005
R5814 dvss.n3279 dvss.n3278 9.3005
R5815 dvss.n3276 dvss.n3275 9.3005
R5816 dvss.n3269 dvss.n3267 9.3005
R5817 dvss.n3945 dvss.n3944 9.3005
R5818 dvss.n229 dvss.n228 9.3005
R5819 dvss.n3929 dvss.n234 9.3005
R5820 dvss.n3912 dvss.n3911 9.3005
R5821 dvss.n3915 dvss.n3914 9.3005
R5822 dvss.n3927 dvss.n3926 9.3005
R5823 dvss.n3930 dvss.n3929 9.3005
R5824 dvss.n4021 dvss.n4020 9.3005
R5825 dvss.n4019 dvss.n3994 9.3005
R5826 dvss.n4032 dvss.n4031 9.3005
R5827 dvss.n4047 dvss.n4046 9.3005
R5828 dvss.n4041 dvss.n4040 9.3005
R5829 dvss.n4038 dvss.n4037 9.3005
R5830 dvss.n4031 dvss.n4029 9.3005
R5831 dvss.n870 dvss.n869 9.3005
R5832 dvss.n869 dvss.n868 9.3005
R5833 dvss.n2662 dvss.n2661 9.3005
R5834 dvss.n2661 dvss.n2657 9.3005
R5835 dvss.n2672 dvss.n2671 9.3005
R5836 dvss.n2671 dvss.n2667 9.3005
R5837 dvss.n2682 dvss.n2681 9.3005
R5838 dvss.n2681 dvss.n2678 9.3005
R5839 dvss.n2709 dvss.n2708 9.3005
R5840 dvss.n2708 dvss.n2707 9.3005
R5841 dvss.n2705 dvss.n2702 9.3005
R5842 dvss.n2705 dvss.n2704 9.3005
R5843 dvss.n2701 dvss.n2698 9.3005
R5844 dvss.n2701 dvss.n2700 9.3005
R5845 dvss.n2721 dvss.n2720 9.3005
R5846 dvss.n2720 dvss.n2717 9.3005
R5847 dvss.n2748 dvss.n2747 9.3005
R5848 dvss.n2747 dvss.n2746 9.3005
R5849 dvss.n2744 dvss.n2741 9.3005
R5850 dvss.n2744 dvss.n2743 9.3005
R5851 dvss.n2740 dvss.n2737 9.3005
R5852 dvss.n2740 dvss.n2739 9.3005
R5853 dvss.n2760 dvss.n2759 9.3005
R5854 dvss.n2759 dvss.n2756 9.3005
R5855 dvss.n2787 dvss.n2786 9.3005
R5856 dvss.n2786 dvss.n2785 9.3005
R5857 dvss.n2783 dvss.n2780 9.3005
R5858 dvss.n2783 dvss.n2782 9.3005
R5859 dvss.n2779 dvss.n2776 9.3005
R5860 dvss.n2779 dvss.n2778 9.3005
R5861 dvss.n2799 dvss.n2798 9.3005
R5862 dvss.n2798 dvss.n2795 9.3005
R5863 dvss.n2826 dvss.n2825 9.3005
R5864 dvss.n2825 dvss.n2824 9.3005
R5865 dvss.n2822 dvss.n2819 9.3005
R5866 dvss.n2822 dvss.n2821 9.3005
R5867 dvss.n2818 dvss.n2815 9.3005
R5868 dvss.n2818 dvss.n2817 9.3005
R5869 dvss.n2838 dvss.n2837 9.3005
R5870 dvss.n2837 dvss.n2834 9.3005
R5871 dvss.n2865 dvss.n2864 9.3005
R5872 dvss.n2864 dvss.n2863 9.3005
R5873 dvss.n2861 dvss.n2858 9.3005
R5874 dvss.n2861 dvss.n2860 9.3005
R5875 dvss.n2857 dvss.n2854 9.3005
R5876 dvss.n2857 dvss.n2856 9.3005
R5877 dvss.n2877 dvss.n2876 9.3005
R5878 dvss.n2876 dvss.n2873 9.3005
R5879 dvss.n3179 dvss.n3178 9.3005
R5880 dvss.n3180 dvss.n3179 9.3005
R5881 dvss.n3175 dvss.n2098 9.3005
R5882 dvss.n3175 dvss.n3174 9.3005
R5883 dvss.n3161 dvss.n2097 9.3005
R5884 dvss.n3159 dvss.n2097 9.3005
R5885 dvss.n3207 dvss.n3206 9.3005
R5886 dvss.n3206 dvss.n3203 9.3005
R5887 dvss.n2074 dvss.n2073 9.3005
R5888 dvss.n2074 dvss.n2004 9.3005
R5889 dvss.n2019 dvss.n2003 9.3005
R5890 dvss.n2017 dvss.n2003 9.3005
R5891 dvss.n3233 dvss.n3232 9.3005
R5892 dvss.n3232 dvss.n3231 9.3005
R5893 dvss.n2061 dvss.n2060 9.3005
R5894 dvss.n2062 dvss.n2061 9.3005
R5895 dvss.n4369 dvss.n4368 9.3005
R5896 dvss.n4369 dvss.n22 9.3005
R5897 dvss.n114 dvss.n21 9.3005
R5898 dvss.n116 dvss.n21 9.3005
R5899 dvss.n4374 dvss.n4373 9.3005
R5900 dvss.n4373 dvss.n4372 9.3005
R5901 dvss.n4356 dvss.n4355 9.3005
R5902 dvss.n4357 dvss.n4356 9.3005
R5903 dvss.n4322 dvss.n4321 9.3005
R5904 dvss.n4323 dvss.n4322 9.3005
R5905 dvss.n4331 dvss.n4329 9.3005
R5906 dvss.n4332 dvss.n4331 9.3005
R5907 dvss.n4339 dvss.n4337 9.3005
R5908 dvss.n4340 dvss.n4339 9.3005
R5909 dvss.n2189 dvss.n2188 9.3005
R5910 dvss.n2188 dvss.n2185 9.3005
R5911 dvss.n2260 dvss.n2259 9.3005
R5912 dvss.n2261 dvss.n2260 9.3005
R5913 dvss.n2256 dvss.n2154 9.3005
R5914 dvss.n2256 dvss.n2255 9.3005
R5915 dvss.n2242 dvss.n2153 9.3005
R5916 dvss.n2240 dvss.n2153 9.3005
R5917 dvss.n2184 dvss.n2183 9.3005
R5918 dvss.n2176 dvss.n2174 9.3005
R5919 dvss.n2190 dvss.n2173 9.3005
R5920 dvss.n2193 dvss.n2192 9.3005
R5921 dvss.n2191 dvss.n2169 9.3005
R5922 dvss.n2200 dvss.n2199 9.3005
R5923 dvss.n2201 dvss.n2168 9.3005
R5924 dvss.n2204 dvss.n2203 9.3005
R5925 dvss.n2202 dvss.n2164 9.3005
R5926 dvss.n2239 dvss.n2238 9.3005
R5927 dvss.n2241 dvss.n2163 9.3005
R5928 dvss.n2245 dvss.n2244 9.3005
R5929 dvss.n2243 dvss.n2156 9.3005
R5930 dvss.n2254 dvss.n2253 9.3005
R5931 dvss.n2159 dvss.n2158 9.3005
R5932 dvss.n2157 dvss.n2151 9.3005
R5933 dvss.n2263 dvss.n2262 9.3005
R5934 dvss.n2258 dvss.n2148 9.3005
R5935 dvss.n2270 dvss.n2269 9.3005
R5936 dvss.n2271 dvss.n2147 9.3005
R5937 dvss.n2516 dvss.n2515 9.3005
R5938 dvss.n3140 dvss.n2647 9.3005
R5939 dvss.n3139 dvss.n2648 9.3005
R5940 dvss.n3138 dvss.n2649 9.3005
R5941 dvss.n3136 dvss.n2650 9.3005
R5942 dvss.n3133 dvss.n2651 9.3005
R5943 dvss.n3132 dvss.n2652 9.3005
R5944 dvss.n3129 dvss.n2653 9.3005
R5945 dvss.n3128 dvss.n2654 9.3005
R5946 dvss.n3125 dvss.n2655 9.3005
R5947 dvss.n3124 dvss.n2656 9.3005
R5948 dvss.n3121 dvss.n2663 9.3005
R5949 dvss.n3120 dvss.n2664 9.3005
R5950 dvss.n3117 dvss.n2665 9.3005
R5951 dvss.n3116 dvss.n2666 9.3005
R5952 dvss.n3113 dvss.n2673 9.3005
R5953 dvss.n3112 dvss.n2674 9.3005
R5954 dvss.n3109 dvss.n2675 9.3005
R5955 dvss.n3108 dvss.n2676 9.3005
R5956 dvss.n3105 dvss.n2677 9.3005
R5957 dvss.n3104 dvss.n2683 9.3005
R5958 dvss.n3101 dvss.n2684 9.3005
R5959 dvss.n3100 dvss.n2685 9.3005
R5960 dvss.n3097 dvss.n2686 9.3005
R5961 dvss.n3096 dvss.n2687 9.3005
R5962 dvss.n3093 dvss.n2688 9.3005
R5963 dvss.n3092 dvss.n2689 9.3005
R5964 dvss.n3089 dvss.n2690 9.3005
R5965 dvss.n3088 dvss.n2691 9.3005
R5966 dvss.n3085 dvss.n2692 9.3005
R5967 dvss.n3084 dvss.n2693 9.3005
R5968 dvss.n3081 dvss.n2694 9.3005
R5969 dvss.n3080 dvss.n2695 9.3005
R5970 dvss.n3077 dvss.n2696 9.3005
R5971 dvss.n3076 dvss.n2697 9.3005
R5972 dvss.n3073 dvss.n2710 9.3005
R5973 dvss.n3072 dvss.n2711 9.3005
R5974 dvss.n3069 dvss.n2712 9.3005
R5975 dvss.n3068 dvss.n2713 9.3005
R5976 dvss.n3065 dvss.n2714 9.3005
R5977 dvss.n3064 dvss.n2715 9.3005
R5978 dvss.n3061 dvss.n2716 9.3005
R5979 dvss.n3060 dvss.n2722 9.3005
R5980 dvss.n3057 dvss.n2723 9.3005
R5981 dvss.n3056 dvss.n2724 9.3005
R5982 dvss.n3053 dvss.n2725 9.3005
R5983 dvss.n3052 dvss.n2726 9.3005
R5984 dvss.n3049 dvss.n2727 9.3005
R5985 dvss.n3048 dvss.n2728 9.3005
R5986 dvss.n3045 dvss.n2729 9.3005
R5987 dvss.n3044 dvss.n2730 9.3005
R5988 dvss.n3041 dvss.n2731 9.3005
R5989 dvss.n3040 dvss.n2732 9.3005
R5990 dvss.n3037 dvss.n2733 9.3005
R5991 dvss.n3036 dvss.n2734 9.3005
R5992 dvss.n3033 dvss.n2735 9.3005
R5993 dvss.n3032 dvss.n2736 9.3005
R5994 dvss.n3029 dvss.n2749 9.3005
R5995 dvss.n3028 dvss.n2750 9.3005
R5996 dvss.n3025 dvss.n2751 9.3005
R5997 dvss.n3024 dvss.n2752 9.3005
R5998 dvss.n3021 dvss.n2753 9.3005
R5999 dvss.n3020 dvss.n2754 9.3005
R6000 dvss.n3017 dvss.n2755 9.3005
R6001 dvss.n3016 dvss.n2761 9.3005
R6002 dvss.n3013 dvss.n2762 9.3005
R6003 dvss.n3012 dvss.n2763 9.3005
R6004 dvss.n3009 dvss.n2764 9.3005
R6005 dvss.n3008 dvss.n2765 9.3005
R6006 dvss.n3005 dvss.n2766 9.3005
R6007 dvss.n3004 dvss.n2767 9.3005
R6008 dvss.n3001 dvss.n2768 9.3005
R6009 dvss.n3000 dvss.n2769 9.3005
R6010 dvss.n2997 dvss.n2770 9.3005
R6011 dvss.n2996 dvss.n2771 9.3005
R6012 dvss.n2993 dvss.n2772 9.3005
R6013 dvss.n2992 dvss.n2773 9.3005
R6014 dvss.n2989 dvss.n2774 9.3005
R6015 dvss.n2988 dvss.n2775 9.3005
R6016 dvss.n2985 dvss.n2788 9.3005
R6017 dvss.n2984 dvss.n2789 9.3005
R6018 dvss.n2981 dvss.n2790 9.3005
R6019 dvss.n2980 dvss.n2791 9.3005
R6020 dvss.n2977 dvss.n2792 9.3005
R6021 dvss.n2976 dvss.n2793 9.3005
R6022 dvss.n2973 dvss.n2794 9.3005
R6023 dvss.n2972 dvss.n2800 9.3005
R6024 dvss.n2969 dvss.n2801 9.3005
R6025 dvss.n2968 dvss.n2802 9.3005
R6026 dvss.n2965 dvss.n2803 9.3005
R6027 dvss.n2964 dvss.n2804 9.3005
R6028 dvss.n2961 dvss.n2805 9.3005
R6029 dvss.n2960 dvss.n2806 9.3005
R6030 dvss.n2957 dvss.n2807 9.3005
R6031 dvss.n2956 dvss.n2808 9.3005
R6032 dvss.n2953 dvss.n2809 9.3005
R6033 dvss.n2952 dvss.n2810 9.3005
R6034 dvss.n2949 dvss.n2811 9.3005
R6035 dvss.n2948 dvss.n2812 9.3005
R6036 dvss.n2945 dvss.n2813 9.3005
R6037 dvss.n2944 dvss.n2814 9.3005
R6038 dvss.n2941 dvss.n2827 9.3005
R6039 dvss.n2940 dvss.n2828 9.3005
R6040 dvss.n2937 dvss.n2829 9.3005
R6041 dvss.n2936 dvss.n2830 9.3005
R6042 dvss.n2933 dvss.n2831 9.3005
R6043 dvss.n2932 dvss.n2832 9.3005
R6044 dvss.n2929 dvss.n2833 9.3005
R6045 dvss.n2928 dvss.n2839 9.3005
R6046 dvss.n2925 dvss.n2840 9.3005
R6047 dvss.n2924 dvss.n2841 9.3005
R6048 dvss.n2921 dvss.n2842 9.3005
R6049 dvss.n2920 dvss.n2843 9.3005
R6050 dvss.n2917 dvss.n2844 9.3005
R6051 dvss.n2916 dvss.n2845 9.3005
R6052 dvss.n2913 dvss.n2846 9.3005
R6053 dvss.n2912 dvss.n2847 9.3005
R6054 dvss.n2909 dvss.n2848 9.3005
R6055 dvss.n2908 dvss.n2849 9.3005
R6056 dvss.n2905 dvss.n2850 9.3005
R6057 dvss.n2904 dvss.n2851 9.3005
R6058 dvss.n2901 dvss.n2852 9.3005
R6059 dvss.n2900 dvss.n2853 9.3005
R6060 dvss.n2897 dvss.n2866 9.3005
R6061 dvss.n2896 dvss.n2867 9.3005
R6062 dvss.n2893 dvss.n2868 9.3005
R6063 dvss.n2892 dvss.n2869 9.3005
R6064 dvss.n2889 dvss.n2870 9.3005
R6065 dvss.n2888 dvss.n2871 9.3005
R6066 dvss.n2885 dvss.n2872 9.3005
R6067 dvss.n2884 dvss.n2878 9.3005
R6068 dvss.n2881 dvss.n2880 9.3005
R6069 dvss.n2879 dvss.n2578 9.3005
R6070 dvss.n3147 dvss.n3146 9.3005
R6071 dvss.n3148 dvss.n2577 9.3005
R6072 dvss.n3151 dvss.n3150 9.3005
R6073 dvss.n3149 dvss.n2109 9.3005
R6074 dvss.n3158 dvss.n3157 9.3005
R6075 dvss.n3160 dvss.n2108 9.3005
R6076 dvss.n3164 dvss.n3163 9.3005
R6077 dvss.n3162 dvss.n2100 9.3005
R6078 dvss.n3173 dvss.n3172 9.3005
R6079 dvss.n2103 dvss.n2102 9.3005
R6080 dvss.n2101 dvss.n2095 9.3005
R6081 dvss.n3182 dvss.n3181 9.3005
R6082 dvss.n3177 dvss.n2092 9.3005
R6083 dvss.n3190 dvss.n3189 9.3005
R6084 dvss.n3191 dvss.n2091 9.3005
R6085 dvss.n3194 dvss.n3193 9.3005
R6086 dvss.n3192 dvss.n2087 9.3005
R6087 dvss.n3202 dvss.n3201 9.3005
R6088 dvss.n2086 dvss.n2085 9.3005
R6089 dvss.n3210 dvss.n3209 9.3005
R6090 dvss.n3208 dvss.n2082 9.3005
R6091 dvss.n3217 dvss.n3216 9.3005
R6092 dvss.n3218 dvss.n2081 9.3005
R6093 dvss.n3221 dvss.n3220 9.3005
R6094 dvss.n3219 dvss.n2077 9.3005
R6095 dvss.n3229 dvss.n3228 9.3005
R6096 dvss.n3230 dvss.n2000 9.3005
R6097 dvss.n3235 dvss.n3234 9.3005
R6098 dvss.n2011 dvss.n2001 9.3005
R6099 dvss.n2016 dvss.n2015 9.3005
R6100 dvss.n2018 dvss.n2009 9.3005
R6101 dvss.n2023 dvss.n2022 9.3005
R6102 dvss.n2021 dvss.n2010 9.3005
R6103 dvss.n2020 dvss.n2005 9.3005
R6104 dvss.n2072 dvss.n2071 9.3005
R6105 dvss.n2070 dvss.n2069 9.3005
R6106 dvss.n2068 dvss.n2031 9.3005
R6107 dvss.n2067 dvss.n2066 9.3005
R6108 dvss.n2065 dvss.n2064 9.3005
R6109 dvss.n2063 dvss.n2034 9.3005
R6110 dvss.n2059 dvss.n2058 9.3005
R6111 dvss.n10 dvss.n9 9.3005
R6112 dvss.n4388 dvss.n4387 9.3005
R6113 dvss.n4386 dvss.n4385 9.3005
R6114 dvss.n4384 dvss.n13 9.3005
R6115 dvss.n4383 dvss.n4382 9.3005
R6116 dvss.n4381 dvss.n4380 9.3005
R6117 dvss.n4379 dvss.n16 9.3005
R6118 dvss.n4378 dvss.n4377 9.3005
R6119 dvss.n4376 dvss.n4375 9.3005
R6120 dvss.n109 dvss.n19 9.3005
R6121 dvss.n118 dvss.n117 9.3005
R6122 dvss.n115 dvss.n108 9.3005
R6123 dvss.n113 dvss.n112 9.3005
R6124 dvss.n111 dvss.n102 9.3005
R6125 dvss.n110 dvss.n23 9.3005
R6126 dvss.n4367 dvss.n4366 9.3005
R6127 dvss.n4365 dvss.n4364 9.3005
R6128 dvss.n4363 dvss.n26 9.3005
R6129 dvss.n4362 dvss.n4361 9.3005
R6130 dvss.n4360 dvss.n4359 9.3005
R6131 dvss.n4358 dvss.n29 9.3005
R6132 dvss.n33 dvss.n32 9.3005
R6133 dvss.n4354 dvss.n4353 9.3005
R6134 dvss.n4352 dvss.n4351 9.3005
R6135 dvss.n4350 dvss.n36 9.3005
R6136 dvss.n4349 dvss.n4348 9.3005
R6137 dvss.n4347 dvss.n4346 9.3005
R6138 dvss.n4345 dvss.n39 9.3005
R6139 dvss.n4344 dvss.n4343 9.3005
R6140 dvss.n4342 dvss.n4341 9.3005
R6141 dvss.n44 dvss.n42 9.3005
R6142 dvss.n4336 dvss.n4335 9.3005
R6143 dvss.n4334 dvss.n4333 9.3005
R6144 dvss.n48 dvss.n47 9.3005
R6145 dvss.n4328 dvss.n4327 9.3005
R6146 dvss.n4326 dvss.n4325 9.3005
R6147 dvss.n4324 dvss.n51 9.3005
R6148 dvss.n4320 dvss.n4319 9.3005
R6149 dvss.n4318 dvss.n4317 9.3005
R6150 dvss.n4316 dvss.n54 9.3005
R6151 dvss.n4315 dvss.n4314 9.3005
R6152 dvss.n1021 dvss.n834 9.3005
R6153 dvss.n1049 dvss.n1023 9.3005
R6154 dvss.n1048 dvss.n1024 9.3005
R6155 dvss.n1047 dvss.n1025 9.3005
R6156 dvss.n1046 dvss.n1026 9.3005
R6157 dvss.n1044 dvss.n1027 9.3005
R6158 dvss.n1041 dvss.n1028 9.3005
R6159 dvss.n1040 dvss.n1032 9.3005
R6160 dvss.n1037 dvss.n1033 9.3005
R6161 dvss.n1036 dvss.n1034 9.3005
R6162 dvss.n826 dvss.n825 9.3005
R6163 dvss.n1056 dvss.n1055 9.3005
R6164 dvss.n1069 dvss.n784 9.3005
R6165 dvss.n1100 dvss.n785 9.3005
R6166 dvss.n1099 dvss.n1098 9.3005
R6167 dvss.n787 dvss.n780 9.3005
R6168 dvss.n1107 dvss.n1106 9.3005
R6169 dvss.n1113 dvss.n773 9.3005
R6170 dvss.n1119 dvss.n774 9.3005
R6171 dvss.n1121 dvss.n1120 9.3005
R6172 dvss.n1123 dvss.n769 9.3005
R6173 dvss.n1130 dvss.n1129 9.3005
R6174 dvss.n1136 dvss.n765 9.3005
R6175 dvss.n766 dvss.n761 9.3005
R6176 dvss.n1151 dvss.n756 9.3005
R6177 dvss.n1143 dvss.n1142 9.3005
R6178 dvss.n1158 dvss.n747 9.3005
R6179 dvss.n1165 dvss.n749 9.3005
R6180 dvss.n1174 dvss.n1166 9.3005
R6181 dvss.n1173 dvss.n743 9.3005
R6182 dvss.n1191 dvss.n735 9.3005
R6183 dvss.n1188 dvss.n740 9.3005
R6184 dvss.n1187 dvss.n1186 9.3005
R6185 dvss.n1198 dvss.n630 9.3005
R6186 dvss.n1263 dvss.n631 9.3005
R6187 dvss.n1262 dvss.n632 9.3005
R6188 dvss.n1261 dvss.n633 9.3005
R6189 dvss.n1207 dvss.n634 9.3005
R6190 dvss.n1210 dvss.n1209 9.3005
R6191 dvss.n1216 dvss.n641 9.3005
R6192 dvss.n1254 dvss.n642 9.3005
R6193 dvss.n1253 dvss.n643 9.3005
R6194 dvss.n1252 dvss.n644 9.3005
R6195 dvss.n1225 dvss.n645 9.3005
R6196 dvss.n1246 dvss.n651 9.3005
R6197 dvss.n1245 dvss.n652 9.3005
R6198 dvss.n1244 dvss.n653 9.3005
R6199 dvss.n1238 dvss.n654 9.3005
R6200 dvss.n681 dvss.n662 9.3005
R6201 dvss.n718 dvss.n664 9.3005
R6202 dvss.n715 dvss.n671 9.3005
R6203 dvss.n714 dvss.n672 9.3005
R6204 dvss.n680 dvss.n675 9.3005
R6205 dvss.n704 dvss.n676 9.3005
R6206 dvss.n701 dvss.n579 9.3005
R6207 dvss.n1464 dvss.n1463 9.3005
R6208 dvss.n1468 dvss.n568 9.3005
R6209 dvss.n1488 dvss.n569 9.3005
R6210 dvss.n1487 dvss.n1486 9.3005
R6211 dvss.n1483 dvss.n570 9.3005
R6212 dvss.n1482 dvss.n1481 9.3005
R6213 dvss.n1496 dvss.n559 9.3005
R6214 dvss.n558 dvss.n557 9.3005
R6215 dvss.n1503 dvss.n1502 9.3005
R6216 dvss.n1509 dvss.n553 9.3005
R6217 dvss.n1516 dvss.n1515 9.3005
R6218 dvss.n1522 dvss.n545 9.3005
R6219 dvss.n1531 dvss.n1530 9.3005
R6220 dvss.n1534 dvss.n1532 9.3005
R6221 dvss.n1533 dvss.n542 9.3005
R6222 dvss.n1546 dvss.n536 9.3005
R6223 dvss.n1552 dvss.n1551 9.3005
R6224 dvss.n1561 dvss.n1553 9.3005
R6225 dvss.n1560 dvss.n532 9.3005
R6226 dvss.n1578 dvss.n524 9.3005
R6227 dvss.n1575 dvss.n529 9.3005
R6228 dvss.n1574 dvss.n1573 9.3005
R6229 dvss.n1584 dvss.n510 9.3005
R6230 dvss.n1746 dvss.n1745 9.3005
R6231 dvss.n1742 dvss.n511 9.3005
R6232 dvss.n1741 dvss.n1588 9.3005
R6233 dvss.n1740 dvss.n1589 9.3005
R6234 dvss.n1737 dvss.n1593 9.3005
R6235 dvss.n1736 dvss.n1594 9.3005
R6236 dvss.n1659 dvss.n1597 9.3005
R6237 dvss.n1732 dvss.n1598 9.3005
R6238 dvss.n1729 dvss.n1603 9.3005
R6239 dvss.n1667 dvss.n1666 9.3005
R6240 dvss.n1669 dvss.n1668 9.3005
R6241 dvss.n1723 dvss.n1609 9.3005
R6242 dvss.n1720 dvss.n1614 9.3005
R6243 dvss.n1719 dvss.n1615 9.3005
R6244 dvss.n1636 dvss.n1616 9.3005
R6245 dvss.n1712 dvss.n1618 9.3005
R6246 dvss.n1709 dvss.n1626 9.3005
R6247 dvss.n1708 dvss.n1627 9.3005
R6248 dvss.n1635 dvss.n1630 9.3005
R6249 dvss.n1698 dvss.n1631 9.3005
R6250 dvss.n1695 dvss.n459 9.3005
R6251 dvss.n3413 dvss.n3412 9.3005
R6252 dvss.n3417 dvss.n449 9.3005
R6253 dvss.n3439 dvss.n3438 9.3005
R6254 dvss.n3435 dvss.n450 9.3005
R6255 dvss.n3434 dvss.n3426 9.3005
R6256 dvss.n3433 dvss.n3432 9.3005
R6257 dvss.n3447 dvss.n440 9.3005
R6258 dvss.n439 dvss.n438 9.3005
R6259 dvss.n3454 dvss.n3453 9.3005
R6260 dvss.n3460 dvss.n434 9.3005
R6261 dvss.n3467 dvss.n3466 9.3005
R6262 dvss.n3473 dvss.n426 9.3005
R6263 dvss.n3482 dvss.n3481 9.3005
R6264 dvss.n3485 dvss.n3483 9.3005
R6265 dvss.n3484 dvss.n423 9.3005
R6266 dvss.n3497 dvss.n417 9.3005
R6267 dvss.n3503 dvss.n3502 9.3005
R6268 dvss.n3512 dvss.n3504 9.3005
R6269 dvss.n3511 dvss.n413 9.3005
R6270 dvss.n3530 dvss.n405 9.3005
R6271 dvss.n3527 dvss.n410 9.3005
R6272 dvss.n3526 dvss.n3525 9.3005
R6273 dvss.n3536 dvss.n391 9.3005
R6274 dvss.n3540 dvss.n3539 9.3005
R6275 dvss.n393 dvss.n385 9.3005
R6276 dvss.n3559 dvss.n3558 9.3005
R6277 dvss.n3555 dvss.n386 9.3005
R6278 dvss.n3554 dvss.n379 9.3005
R6279 dvss.n3566 dvss.n3565 9.3005
R6280 dvss.n3572 dvss.n374 9.3005
R6281 dvss.n3576 dvss.n3575 9.3005
R6282 dvss.n375 dvss.n369 9.3005
R6283 dvss.n3586 dvss.n3585 9.3005
R6284 dvss.n3598 dvss.n364 9.3005
R6285 dvss.n3602 dvss.n3601 9.3005
R6286 dvss.n3592 dvss.n357 9.3005
R6287 dvss.n3610 dvss.n3609 9.3005
R6288 dvss.n3613 dvss.n353 9.3005
R6289 dvss.n3619 dvss.n3618 9.3005
R6290 dvss.n3625 dvss.n348 9.3005
R6291 dvss.n3633 dvss.n3632 9.3005
R6292 dvss.n3647 dvss.n337 9.3005
R6293 dvss.n3644 dvss.n3642 9.3005
R6294 dvss.n3643 dvss.n331 9.3005
R6295 dvss.n3654 dvss.n3653 9.3005
R6296 dvss.n3657 dvss.n3655 9.3005
R6297 dvss.n3656 dvss.n326 9.3005
R6298 dvss.n3671 dvss.n319 9.3005
R6299 dvss.n3670 dvss.n320 9.3005
R6300 dvss.n3669 dvss.n3668 9.3005
R6301 dvss.n3679 dvss.n310 9.3005
R6302 dvss.n3686 dvss.n3685 9.3005
R6303 dvss.n3694 dvss.n3687 9.3005
R6304 dvss.n3689 dvss.n307 9.3005
R6305 dvss.n3704 dvss.n301 9.3005
R6306 dvss.n3705 dvss.n296 9.3005
R6307 dvss.n3718 dvss.n3717 9.3005
R6308 dvss.n3714 dvss.n297 9.3005
R6309 dvss.n3713 dvss.n292 9.3005
R6310 dvss.n3729 dvss.n286 9.3005
R6311 dvss.n3735 dvss.n3734 9.3005
R6312 dvss.n3744 dvss.n3736 9.3005
R6313 dvss.n3743 dvss.n282 9.3005
R6314 dvss.n3761 dvss.n274 9.3005
R6315 dvss.n3758 dvss.n279 9.3005
R6316 dvss.n3757 dvss.n3756 9.3005
R6317 dvss.n3767 dvss.n265 9.3005
R6318 dvss.n3877 dvss.n3876 9.3005
R6319 dvss.n3873 dvss.n266 9.3005
R6320 dvss.n3872 dvss.n3771 9.3005
R6321 dvss.n3871 dvss.n3772 9.3005
R6322 dvss.n3868 dvss.n3776 9.3005
R6323 dvss.n3867 dvss.n3777 9.3005
R6324 dvss.n3808 dvss.n3780 9.3005
R6325 dvss.n3863 dvss.n3781 9.3005
R6326 dvss.n3860 dvss.n3786 9.3005
R6327 dvss.n3805 dvss.n3804 9.3005
R6328 dvss.n3807 dvss.n3806 9.3005
R6329 dvss.n3854 dvss.n3792 9.3005
R6330 dvss.n3851 dvss.n3797 9.3005
R6331 dvss.n3850 dvss.n3841 9.3005
R6332 dvss.n3842 dvss.n125 9.3005
R6333 dvss.n4149 dvss.n4148 9.3005
R6334 dvss.n4145 dvss.n126 9.3005
R6335 dvss.n4144 dvss.n130 9.3005
R6336 dvss.n203 dvss.n133 9.3005
R6337 dvss.n205 dvss.n204 9.3005
R6338 dvss.n211 dvss.n192 9.3005
R6339 dvss.n213 dvss.n212 9.3005
R6340 dvss.n4132 dvss.n139 9.3005
R6341 dvss.n4129 dvss.n144 9.3005
R6342 dvss.n4128 dvss.n145 9.3005
R6343 dvss.n4127 dvss.n146 9.3005
R6344 dvss.n4124 dvss.n150 9.3005
R6345 dvss.n4123 dvss.n151 9.3005
R6346 dvss.n4075 dvss.n154 9.3005
R6347 dvss.n4119 dvss.n155 9.3005
R6348 dvss.n4116 dvss.n160 9.3005
R6349 dvss.n4083 dvss.n4082 9.3005
R6350 dvss.n4085 dvss.n4084 9.3005
R6351 dvss.n4110 dvss.n166 9.3005
R6352 dvss.n4107 dvss.n171 9.3005
R6353 dvss.n4106 dvss.n172 9.3005
R6354 dvss.n4098 dvss.n99 9.3005
R6355 dvss.n4191 dvss.n4190 9.3005
R6356 dvss.n4193 dvss.n93 9.3005
R6357 dvss.n4202 dvss.n4201 9.3005
R6358 dvss.n4212 dvss.n89 9.3005
R6359 dvss.n4209 dvss.n84 9.3005
R6360 dvss.n4220 dvss.n4219 9.3005
R6361 dvss.n4218 dvss.n74 9.3005
R6362 dvss.n4230 dvss.n4229 9.3005
R6363 dvss.n4233 dvss.n70 9.3005
R6364 dvss.n4235 dvss.n4234 9.3005
R6365 dvss.n4241 dvss.n64 9.3005
R6366 dvss.n1008 dvss.n841 9.3005
R6367 dvss.n1007 dvss.n842 9.3005
R6368 dvss.n847 dvss.n843 9.3005
R6369 dvss.n1001 dvss.n848 9.3005
R6370 dvss.n1000 dvss.n849 9.3005
R6371 dvss.n999 dvss.n850 9.3005
R6372 dvss.n855 dvss.n851 9.3005
R6373 dvss.n992 dvss.n859 9.3005
R6374 dvss.n991 dvss.n860 9.3005
R6375 dvss.n990 dvss.n861 9.3005
R6376 dvss.n871 dvss.n862 9.3005
R6377 dvss.n984 dvss.n872 9.3005
R6378 dvss.n983 dvss.n873 9.3005
R6379 dvss.n982 dvss.n874 9.3005
R6380 dvss.n884 dvss.n875 9.3005
R6381 dvss.n976 dvss.n885 9.3005
R6382 dvss.n975 dvss.n886 9.3005
R6383 dvss.n974 dvss.n887 9.3005
R6384 dvss.n891 dvss.n888 9.3005
R6385 dvss.n968 dvss.n892 9.3005
R6386 dvss.n967 dvss.n893 9.3005
R6387 dvss.n966 dvss.n894 9.3005
R6388 dvss.n913 dvss.n895 9.3005
R6389 dvss.n960 dvss.n899 9.3005
R6390 dvss.n959 dvss.n900 9.3005
R6391 dvss.n958 dvss.n901 9.3005
R6392 dvss.n921 dvss.n902 9.3005
R6393 dvss.n925 dvss.n906 9.3005
R6394 dvss.n949 dvss.n926 9.3005
R6395 dvss.n948 dvss.n927 9.3005
R6396 dvss.n947 dvss.n928 9.3005
R6397 dvss.n938 dvss.n929 9.3005
R6398 dvss.n941 dvss.n940 9.3005
R6399 dvss.n939 dvss.n622 9.3005
R6400 dvss.n1272 dvss.n1271 9.3005
R6401 dvss.n1273 dvss.n621 9.3005
R6402 dvss.n1276 dvss.n1275 9.3005
R6403 dvss.n1274 dvss.n618 9.3005
R6404 dvss.n1283 dvss.n1282 9.3005
R6405 dvss.n1284 dvss.n617 9.3005
R6406 dvss.n1288 dvss.n1287 9.3005
R6407 dvss.n1286 dvss.n613 9.3005
R6408 dvss.n1295 dvss.n1294 9.3005
R6409 dvss.n1296 dvss.n609 9.3005
R6410 dvss.n1303 dvss.n1302 9.3005
R6411 dvss.n610 dvss.n605 9.3005
R6412 dvss.n1311 dvss.n1310 9.3005
R6413 dvss.n604 dvss.n599 9.3005
R6414 dvss.n1318 dvss.n1317 9.3005
R6415 dvss.n601 dvss.n596 9.3005
R6416 dvss.n1326 dvss.n1325 9.3005
R6417 dvss.n1327 dvss.n591 9.3005
R6418 dvss.n1333 dvss.n1332 9.3005
R6419 dvss.n593 dvss.n588 9.3005
R6420 dvss.n1340 dvss.n1339 9.3005
R6421 dvss.n1346 dvss.n586 9.3005
R6422 dvss.n1456 dvss.n1455 9.3005
R6423 dvss.n1454 dvss.n587 9.3005
R6424 dvss.n1453 dvss.n1452 9.3005
R6425 dvss.n1451 dvss.n1450 9.3005
R6426 dvss.n1449 dvss.n1349 9.3005
R6427 dvss.n1448 dvss.n1447 9.3005
R6428 dvss.n1446 dvss.n1445 9.3005
R6429 dvss.n1444 dvss.n1352 9.3005
R6430 dvss.n1355 dvss.n1354 9.3005
R6431 dvss.n1439 dvss.n1438 9.3005
R6432 dvss.n1437 dvss.n1436 9.3005
R6433 dvss.n1361 dvss.n1358 9.3005
R6434 dvss.n1430 dvss.n1429 9.3005
R6435 dvss.n1428 dvss.n1427 9.3005
R6436 dvss.n1365 dvss.n1364 9.3005
R6437 dvss.n1422 dvss.n1421 9.3005
R6438 dvss.n1420 dvss.n1419 9.3005
R6439 dvss.n1418 dvss.n1368 9.3005
R6440 dvss.n1372 dvss.n1371 9.3005
R6441 dvss.n1412 dvss.n1411 9.3005
R6442 dvss.n1410 dvss.n1409 9.3005
R6443 dvss.n1403 dvss.n502 9.3005
R6444 dvss.n1755 dvss.n1754 9.3005
R6445 dvss.n1756 dvss.n501 9.3005
R6446 dvss.n1759 dvss.n1758 9.3005
R6447 dvss.n1757 dvss.n498 9.3005
R6448 dvss.n1766 dvss.n1765 9.3005
R6449 dvss.n1767 dvss.n497 9.3005
R6450 dvss.n1771 dvss.n1770 9.3005
R6451 dvss.n1769 dvss.n493 9.3005
R6452 dvss.n1778 dvss.n1777 9.3005
R6453 dvss.n1779 dvss.n489 9.3005
R6454 dvss.n1786 dvss.n1785 9.3005
R6455 dvss.n490 dvss.n485 9.3005
R6456 dvss.n1794 dvss.n1793 9.3005
R6457 dvss.n484 dvss.n479 9.3005
R6458 dvss.n1801 dvss.n1800 9.3005
R6459 dvss.n481 dvss.n476 9.3005
R6460 dvss.n1809 dvss.n1808 9.3005
R6461 dvss.n1810 dvss.n471 9.3005
R6462 dvss.n1816 dvss.n1815 9.3005
R6463 dvss.n473 dvss.n468 9.3005
R6464 dvss.n1823 dvss.n1822 9.3005
R6465 dvss.n1829 dvss.n466 9.3005
R6466 dvss.n3405 dvss.n3404 9.3005
R6467 dvss.n3403 dvss.n467 9.3005
R6468 dvss.n3402 dvss.n3401 9.3005
R6469 dvss.n3400 dvss.n3399 9.3005
R6470 dvss.n3398 dvss.n1832 9.3005
R6471 dvss.n3397 dvss.n3396 9.3005
R6472 dvss.n3395 dvss.n3394 9.3005
R6473 dvss.n3393 dvss.n1835 9.3005
R6474 dvss.n1838 dvss.n1837 9.3005
R6475 dvss.n3388 dvss.n3387 9.3005
R6476 dvss.n3386 dvss.n3385 9.3005
R6477 dvss.n1844 dvss.n1841 9.3005
R6478 dvss.n3379 dvss.n3378 9.3005
R6479 dvss.n3377 dvss.n3376 9.3005
R6480 dvss.n1848 dvss.n1847 9.3005
R6481 dvss.n3371 dvss.n3370 9.3005
R6482 dvss.n3369 dvss.n3368 9.3005
R6483 dvss.n3367 dvss.n1851 9.3005
R6484 dvss.n1855 dvss.n1854 9.3005
R6485 dvss.n3361 dvss.n3360 9.3005
R6486 dvss.n3359 dvss.n3358 9.3005
R6487 dvss.n3352 dvss.n1858 9.3005
R6488 dvss.n3351 dvss.n3350 9.3005
R6489 dvss.n3349 dvss.n3348 9.3005
R6490 dvss.n3347 dvss.n1861 9.3005
R6491 dvss.n3346 dvss.n3345 9.3005
R6492 dvss.n3344 dvss.n3343 9.3005
R6493 dvss.n3342 dvss.n1864 9.3005
R6494 dvss.n3341 dvss.n3340 9.3005
R6495 dvss.n3339 dvss.n3338 9.3005
R6496 dvss.n1869 dvss.n1867 9.3005
R6497 dvss.n3333 dvss.n3332 9.3005
R6498 dvss.n3331 dvss.n3330 9.3005
R6499 dvss.n1875 dvss.n1872 9.3005
R6500 dvss.n3324 dvss.n3323 9.3005
R6501 dvss.n3322 dvss.n3321 9.3005
R6502 dvss.n1879 dvss.n1878 9.3005
R6503 dvss.n3316 dvss.n3315 9.3005
R6504 dvss.n3314 dvss.n3313 9.3005
R6505 dvss.n3312 dvss.n1882 9.3005
R6506 dvss.n1886 dvss.n1885 9.3005
R6507 dvss.n3306 dvss.n3305 9.3005
R6508 dvss.n3304 dvss.n3303 9.3005
R6509 dvss.n3302 dvss.n1889 9.3005
R6510 dvss.n3301 dvss.n3300 9.3005
R6511 dvss.n3299 dvss.n3298 9.3005
R6512 dvss.n3297 dvss.n1892 9.3005
R6513 dvss.n3296 dvss.n3295 9.3005
R6514 dvss.n3294 dvss.n3293 9.3005
R6515 dvss.n3292 dvss.n1895 9.3005
R6516 dvss.n3291 dvss.n3290 9.3005
R6517 dvss.n3289 dvss.n3288 9.3005
R6518 dvss.n1900 dvss.n1898 9.3005
R6519 dvss.n3283 dvss.n3282 9.3005
R6520 dvss.n3281 dvss.n3280 9.3005
R6521 dvss.n1906 dvss.n1903 9.3005
R6522 dvss.n3274 dvss.n3273 9.3005
R6523 dvss.n3272 dvss.n3271 9.3005
R6524 dvss.n1910 dvss.n1909 9.3005
R6525 dvss.n3266 dvss.n3265 9.3005
R6526 dvss.n3264 dvss.n3263 9.3005
R6527 dvss.n3262 dvss.n1913 9.3005
R6528 dvss.n1917 dvss.n1916 9.3005
R6529 dvss.n3256 dvss.n3255 9.3005
R6530 dvss.n3254 dvss.n3253 9.3005
R6531 dvss.n3252 dvss.n256 9.3005
R6532 dvss.n3886 dvss.n3885 9.3005
R6533 dvss.n3887 dvss.n255 9.3005
R6534 dvss.n3890 dvss.n3889 9.3005
R6535 dvss.n3888 dvss.n252 9.3005
R6536 dvss.n3897 dvss.n3896 9.3005
R6537 dvss.n3898 dvss.n251 9.3005
R6538 dvss.n3902 dvss.n3901 9.3005
R6539 dvss.n3900 dvss.n247 9.3005
R6540 dvss.n3909 dvss.n3908 9.3005
R6541 dvss.n3910 dvss.n243 9.3005
R6542 dvss.n3917 dvss.n3916 9.3005
R6543 dvss.n244 dvss.n239 9.3005
R6544 dvss.n3925 dvss.n3924 9.3005
R6545 dvss.n238 dvss.n233 9.3005
R6546 dvss.n3932 dvss.n3931 9.3005
R6547 dvss.n235 dvss.n230 9.3005
R6548 dvss.n3940 dvss.n3939 9.3005
R6549 dvss.n3941 dvss.n225 9.3005
R6550 dvss.n3947 dvss.n3946 9.3005
R6551 dvss.n227 dvss.n222 9.3005
R6552 dvss.n3954 dvss.n3953 9.3005
R6553 dvss.n3955 dvss.n220 9.3005
R6554 dvss.n4062 dvss.n4061 9.3005
R6555 dvss.n4060 dvss.n221 9.3005
R6556 dvss.n4059 dvss.n4058 9.3005
R6557 dvss.n4057 dvss.n4056 9.3005
R6558 dvss.n4055 dvss.n3958 9.3005
R6559 dvss.n4054 dvss.n4053 9.3005
R6560 dvss.n4052 dvss.n4051 9.3005
R6561 dvss.n4050 dvss.n3961 9.3005
R6562 dvss.n3964 dvss.n3963 9.3005
R6563 dvss.n4045 dvss.n4044 9.3005
R6564 dvss.n4043 dvss.n4042 9.3005
R6565 dvss.n3970 dvss.n3967 9.3005
R6566 dvss.n4036 dvss.n4035 9.3005
R6567 dvss.n4034 dvss.n4033 9.3005
R6568 dvss.n3990 dvss.n3989 9.3005
R6569 dvss.n4028 dvss.n4027 9.3005
R6570 dvss.n4026 dvss.n4025 9.3005
R6571 dvss.n4024 dvss.n3993 9.3005
R6572 dvss.n3997 dvss.n3996 9.3005
R6573 dvss.n4018 dvss.n4017 9.3005
R6574 dvss.n4016 dvss.n4015 9.3005
R6575 dvss.n4014 dvss.n4012 9.3005
R6576 dvss.n4013 dvss.n62 9.3005
R6577 dvss.n4307 dvss.n4306 9.3005
R6578 dvss.n4305 dvss.n63 9.3005
R6579 dvss.n4304 dvss.n4303 9.3005
R6580 dvss.n1020 dvss.n1019 9.3005
R6581 dvss.n1022 dvss.n804 9.3005
R6582 dvss.n1088 dvss.n805 9.3005
R6583 dvss.n1087 dvss.n806 9.3005
R6584 dvss.n1086 dvss.n807 9.3005
R6585 dvss.n1085 dvss.n808 9.3005
R6586 dvss.n1083 dvss.n809 9.3005
R6587 dvss.n1080 dvss.n810 9.3005
R6588 dvss.n1079 dvss.n811 9.3005
R6589 dvss.n1076 dvss.n812 9.3005
R6590 dvss.n1075 dvss.n813 9.3005
R6591 dvss.n1072 dvss.n814 9.3005
R6592 dvss.n1071 dvss.n1070 9.3005
R6593 dvss.n1068 dvss.n795 9.3005
R6594 dvss.n1059 dvss.n786 9.3005
R6595 dvss.n1097 dvss.n1096 9.3005
R6596 dvss.n789 dvss.n788 9.3005
R6597 dvss.n1107 dvss.n779 9.3005
R6598 dvss.n1114 dvss.n1113 9.3005
R6599 dvss.n1115 dvss.n774 9.3005
R6600 dvss.n1121 dvss.n772 9.3005
R6601 dvss.n1124 dvss.n1123 9.3005
R6602 dvss.n1130 dvss.n764 9.3005
R6603 dvss.n1137 dvss.n1136 9.3005
R6604 dvss.n766 dvss.n757 9.3005
R6605 dvss.n1151 dvss.n1150 9.3005
R6606 dvss.n1142 dvss.n752 9.3005
R6607 dvss.n1159 dvss.n1158 9.3005
R6608 dvss.n749 dvss.n746 9.3005
R6609 dvss.n1175 dvss.n1174 9.3005
R6610 dvss.n1173 dvss.n737 9.3005
R6611 dvss.n1191 dvss.n1190 9.3005
R6612 dvss.n1189 dvss.n1188 9.3005
R6613 dvss.n1187 dvss.n729 9.3005
R6614 dvss.n1199 dvss.n1198 9.3005
R6615 dvss.n1200 dvss.n631 9.3005
R6616 dvss.n1201 dvss.n632 9.3005
R6617 dvss.n725 dvss.n633 9.3005
R6618 dvss.n1207 dvss.n1206 9.3005
R6619 dvss.n1210 dvss.n723 9.3005
R6620 dvss.n1217 dvss.n1216 9.3005
R6621 dvss.n1218 dvss.n642 9.3005
R6622 dvss.n1221 dvss.n643 9.3005
R6623 dvss.n1222 dvss.n644 9.3005
R6624 dvss.n1225 dvss.n1224 9.3005
R6625 dvss.n1223 dvss.n651 9.3005
R6626 dvss.n660 dvss.n652 9.3005
R6627 dvss.n1240 dvss.n653 9.3005
R6628 dvss.n1239 dvss.n1238 9.3005
R6629 dvss.n662 dvss.n661 9.3005
R6630 dvss.n718 dvss.n717 9.3005
R6631 dvss.n716 dvss.n715 9.3005
R6632 dvss.n714 dvss.n667 9.3005
R6633 dvss.n677 dvss.n675 9.3005
R6634 dvss.n704 dvss.n703 9.3005
R6635 dvss.n702 dvss.n701 9.3005
R6636 dvss.n1464 dvss.n571 9.3005
R6637 dvss.n1469 dvss.n1468 9.3005
R6638 dvss.n1470 dvss.n569 9.3005
R6639 dvss.n1486 dvss.n1485 9.3005
R6640 dvss.n1484 dvss.n1483 9.3005
R6641 dvss.n1482 dvss.n560 9.3005
R6642 dvss.n1496 dvss.n1495 9.3005
R6643 dvss.n1494 dvss.n558 9.3005
R6644 dvss.n1502 dvss.n554 9.3005
R6645 dvss.n1509 dvss.n1508 9.3005
R6646 dvss.n1515 dvss.n548 9.3005
R6647 dvss.n1522 dvss.n1521 9.3005
R6648 dvss.n1530 dvss.n544 9.3005
R6649 dvss.n1535 dvss.n1534 9.3005
R6650 dvss.n1533 dvss.n539 9.3005
R6651 dvss.n1546 dvss.n1545 9.3005
R6652 dvss.n1551 dvss.n535 9.3005
R6653 dvss.n1562 dvss.n1561 9.3005
R6654 dvss.n1560 dvss.n526 9.3005
R6655 dvss.n1578 dvss.n1577 9.3005
R6656 dvss.n1576 dvss.n1575 9.3005
R6657 dvss.n1574 dvss.n513 9.3005
R6658 dvss.n1585 dvss.n1584 9.3005
R6659 dvss.n1745 dvss.n1744 9.3005
R6660 dvss.n1743 dvss.n1742 9.3005
R6661 dvss.n1741 dvss.n1587 9.3005
R6662 dvss.n1740 dvss.n1739 9.3005
R6663 dvss.n1738 dvss.n1737 9.3005
R6664 dvss.n1736 dvss.n1592 9.3005
R6665 dvss.n1599 dvss.n1597 9.3005
R6666 dvss.n1732 dvss.n1731 9.3005
R6667 dvss.n1730 dvss.n1729 9.3005
R6668 dvss.n1667 dvss.n1602 9.3005
R6669 dvss.n1668 dvss.n1610 9.3005
R6670 dvss.n1723 dvss.n1722 9.3005
R6671 dvss.n1721 dvss.n1720 9.3005
R6672 dvss.n1719 dvss.n1613 9.3005
R6673 dvss.n1619 dvss.n1616 9.3005
R6674 dvss.n1712 dvss.n1711 9.3005
R6675 dvss.n1710 dvss.n1709 9.3005
R6676 dvss.n1708 dvss.n1622 9.3005
R6677 dvss.n1632 dvss.n1630 9.3005
R6678 dvss.n1698 dvss.n1697 9.3005
R6679 dvss.n1696 dvss.n1695 9.3005
R6680 dvss.n3413 dvss.n451 9.3005
R6681 dvss.n3418 dvss.n3417 9.3005
R6682 dvss.n3438 dvss.n3437 9.3005
R6683 dvss.n3436 dvss.n3435 9.3005
R6684 dvss.n3434 dvss.n3425 9.3005
R6685 dvss.n3433 dvss.n441 9.3005
R6686 dvss.n3447 dvss.n3446 9.3005
R6687 dvss.n3445 dvss.n439 9.3005
R6688 dvss.n3453 dvss.n435 9.3005
R6689 dvss.n3460 dvss.n3459 9.3005
R6690 dvss.n3466 dvss.n429 9.3005
R6691 dvss.n3473 dvss.n3472 9.3005
R6692 dvss.n3481 dvss.n425 9.3005
R6693 dvss.n3486 dvss.n3485 9.3005
R6694 dvss.n3484 dvss.n420 9.3005
R6695 dvss.n3497 dvss.n3496 9.3005
R6696 dvss.n3502 dvss.n416 9.3005
R6697 dvss.n3513 dvss.n3512 9.3005
R6698 dvss.n3511 dvss.n407 9.3005
R6699 dvss.n3530 dvss.n3529 9.3005
R6700 dvss.n3528 dvss.n3527 9.3005
R6701 dvss.n3526 dvss.n394 9.3005
R6702 dvss.n3537 dvss.n3536 9.3005
R6703 dvss.n3539 dvss.n3538 9.3005
R6704 dvss.n393 dvss.n387 9.3005
R6705 dvss.n3558 dvss.n3557 9.3005
R6706 dvss.n3556 dvss.n3555 9.3005
R6707 dvss.n3554 dvss.n3553 9.3005
R6708 dvss.n3566 dvss.n377 9.3005
R6709 dvss.n3573 dvss.n3572 9.3005
R6710 dvss.n3575 dvss.n3574 9.3005
R6711 dvss.n375 dvss.n372 9.3005
R6712 dvss.n3586 dvss.n365 9.3005
R6713 dvss.n3599 dvss.n3598 9.3005
R6714 dvss.n3601 dvss.n3600 9.3005
R6715 dvss.n3592 dvss.n355 9.3005
R6716 dvss.n3611 dvss.n3610 9.3005
R6717 dvss.n3613 dvss.n3612 9.3005
R6718 dvss.n3618 dvss.n349 9.3005
R6719 dvss.n3625 dvss.n3624 9.3005
R6720 dvss.n3632 dvss.n339 9.3005
R6721 dvss.n3647 dvss.n3646 9.3005
R6722 dvss.n3645 dvss.n3644 9.3005
R6723 dvss.n3643 dvss.n342 9.3005
R6724 dvss.n3653 dvss.n329 9.3005
R6725 dvss.n3658 dvss.n3657 9.3005
R6726 dvss.n3656 dvss.n317 9.3005
R6727 dvss.n3672 dvss.n3671 9.3005
R6728 dvss.n3670 dvss.n318 9.3005
R6729 dvss.n3669 dvss.n312 9.3005
R6730 dvss.n3679 dvss.n3678 9.3005
R6731 dvss.n3685 dvss.n309 9.3005
R6732 dvss.n3695 dvss.n3694 9.3005
R6733 dvss.n3689 dvss.n302 9.3005
R6734 dvss.n3704 dvss.n3703 9.3005
R6735 dvss.n3705 dvss.n298 9.3005
R6736 dvss.n3717 dvss.n3716 9.3005
R6737 dvss.n3715 dvss.n3714 9.3005
R6738 dvss.n3713 dvss.n289 9.3005
R6739 dvss.n3729 dvss.n3728 9.3005
R6740 dvss.n3734 dvss.n285 9.3005
R6741 dvss.n3745 dvss.n3744 9.3005
R6742 dvss.n3743 dvss.n276 9.3005
R6743 dvss.n3761 dvss.n3760 9.3005
R6744 dvss.n3759 dvss.n3758 9.3005
R6745 dvss.n3757 dvss.n268 9.3005
R6746 dvss.n3768 dvss.n3767 9.3005
R6747 dvss.n3876 dvss.n3875 9.3005
R6748 dvss.n3874 dvss.n3873 9.3005
R6749 dvss.n3872 dvss.n3770 9.3005
R6750 dvss.n3871 dvss.n3870 9.3005
R6751 dvss.n3869 dvss.n3868 9.3005
R6752 dvss.n3867 dvss.n3775 9.3005
R6753 dvss.n3782 dvss.n3780 9.3005
R6754 dvss.n3863 dvss.n3862 9.3005
R6755 dvss.n3861 dvss.n3860 9.3005
R6756 dvss.n3805 dvss.n3785 9.3005
R6757 dvss.n3806 dvss.n3793 9.3005
R6758 dvss.n3854 dvss.n3853 9.3005
R6759 dvss.n3852 dvss.n3851 9.3005
R6760 dvss.n3850 dvss.n3796 9.3005
R6761 dvss.n3842 dvss.n127 9.3005
R6762 dvss.n4148 dvss.n4147 9.3005
R6763 dvss.n4146 dvss.n4145 9.3005
R6764 dvss.n4144 dvss.n129 9.3005
R6765 dvss.n199 dvss.n133 9.3005
R6766 dvss.n204 dvss.n193 9.3005
R6767 dvss.n211 dvss.n210 9.3005
R6768 dvss.n212 dvss.n140 9.3005
R6769 dvss.n4132 dvss.n4131 9.3005
R6770 dvss.n4130 dvss.n4129 9.3005
R6771 dvss.n4128 dvss.n143 9.3005
R6772 dvss.n4127 dvss.n4126 9.3005
R6773 dvss.n4125 dvss.n4124 9.3005
R6774 dvss.n4123 dvss.n149 9.3005
R6775 dvss.n156 dvss.n154 9.3005
R6776 dvss.n4119 dvss.n4118 9.3005
R6777 dvss.n4117 dvss.n4116 9.3005
R6778 dvss.n4083 dvss.n159 9.3005
R6779 dvss.n4084 dvss.n167 9.3005
R6780 dvss.n4110 dvss.n4109 9.3005
R6781 dvss.n4108 dvss.n4107 9.3005
R6782 dvss.n4106 dvss.n170 9.3005
R6783 dvss.n4098 dvss.n4097 9.3005
R6784 dvss.n4191 dvss.n98 9.3005
R6785 dvss.n4194 dvss.n4193 9.3005
R6786 dvss.n4202 dvss.n91 9.3005
R6787 dvss.n4212 dvss.n4211 9.3005
R6788 dvss.n4210 dvss.n4209 9.3005
R6789 dvss.n4219 dvss.n82 9.3005
R6790 dvss.n4218 dvss.n71 9.3005
R6791 dvss.n4231 dvss.n4230 9.3005
R6792 dvss.n4233 dvss.n4232 9.3005
R6793 dvss.n4234 dvss.n65 9.3005
R6794 dvss.n4241 dvss.n4240 9.3005
R6795 dvss.n2537 dvss.n2536 9.3005
R6796 dvss.n2535 dvss.n2133 9.3005
R6797 dvss.n2548 dvss.n2547 9.3005
R6798 dvss.n2563 dvss.n2562 9.3005
R6799 dvss.n2557 dvss.n2556 9.3005
R6800 dvss.n2554 dvss.n2553 9.3005
R6801 dvss.n2547 dvss.n2545 9.3005
R6802 dvss.n2570 dvss.n2114 9.3005
R6803 dvss.n2569 dvss.n2568 9.3005
R6804 dvss.n2567 dvss.n2566 9.3005
R6805 dvss.n2119 dvss.n2117 9.3005
R6806 dvss.n2561 dvss.n2560 9.3005
R6807 dvss.n2559 dvss.n2558 9.3005
R6808 dvss.n2125 dvss.n2122 9.3005
R6809 dvss.n2552 dvss.n2551 9.3005
R6810 dvss.n2550 dvss.n2549 9.3005
R6811 dvss.n2129 dvss.n2128 9.3005
R6812 dvss.n2544 dvss.n2543 9.3005
R6813 dvss.n2542 dvss.n2541 9.3005
R6814 dvss.n2540 dvss.n2132 9.3005
R6815 dvss.n2136 dvss.n2135 9.3005
R6816 dvss.n2534 dvss.n2533 9.3005
R6817 dvss.n2532 dvss.n2531 9.3005
R6818 dvss.n2530 dvss.n2139 9.3005
R6819 dvss.n2529 dvss.n2528 9.3005
R6820 dvss.n2527 dvss.n2526 9.3005
R6821 dvss.n2525 dvss.n2142 9.3005
R6822 dvss.n2524 dvss.n2523 9.3005
R6823 dvss.n2354 dvss.n2353 9.3005
R6824 dvss.n2352 dvss.n2351 9.3005
R6825 dvss.n2350 dvss.n2349 9.3005
R6826 dvss.n2348 dvss.n2342 9.3005
R6827 dvss.n2347 dvss.n2346 9.3005
R6828 dvss.n2321 dvss.n2320 9.3005
R6829 dvss.n2323 dvss.n2315 9.3005
R6830 dvss.n2327 dvss.n2326 9.3005
R6831 dvss.n2328 dvss.n2314 9.3005
R6832 dvss.n2330 dvss.n2329 9.3005
R6833 dvss.n2332 dvss.n2312 9.3005
R6834 dvss.n2336 dvss.n2335 9.3005
R6835 dvss.n2337 dvss.n2309 9.3005
R6836 dvss.n2362 dvss.n2361 9.3005
R6837 dvss.n2360 dvss.n2359 9.3005
R6838 dvss.n2357 dvss.n2338 9.3005
R6839 dvss.n2356 dvss.n2355 9.3005
R6840 dvss.n2429 dvss.n2376 9.3005
R6841 dvss.n2428 dvss.n2427 9.3005
R6842 dvss.n2426 dvss.n2378 9.3005
R6843 dvss.n2425 dvss.n2424 9.3005
R6844 dvss.n2422 dvss.n2421 9.3005
R6845 dvss.n2396 dvss.n2395 9.3005
R6846 dvss.n2397 dvss.n2389 9.3005
R6847 dvss.n2399 dvss.n2398 9.3005
R6848 dvss.n2401 dvss.n2387 9.3005
R6849 dvss.n2405 dvss.n2404 9.3005
R6850 dvss.n2406 dvss.n2386 9.3005
R6851 dvss.n2408 dvss.n2407 9.3005
R6852 dvss.n2410 dvss.n2384 9.3005
R6853 dvss.n2414 dvss.n2413 9.3005
R6854 dvss.n2416 dvss.n2415 9.3005
R6855 dvss.n2418 dvss.n2380 9.3005
R6856 dvss.n2420 dvss.n2419 9.3005
R6857 dvss.n2503 dvss.n2502 9.3005
R6858 dvss.n2506 dvss.n2505 9.3005
R6859 dvss.n2507 dvss.n2275 9.3005
R6860 dvss.n2509 dvss.n2508 9.3005
R6861 dvss.n2510 dvss.n2273 9.3005
R6862 dvss.n2293 dvss.n2292 9.3005
R6863 dvss.n2294 dvss.n2286 9.3005
R6864 dvss.n2296 dvss.n2295 9.3005
R6865 dvss.n2298 dvss.n2284 9.3005
R6866 dvss.n2302 dvss.n2301 9.3005
R6867 dvss.n2303 dvss.n2283 9.3005
R6868 dvss.n2305 dvss.n2304 9.3005
R6869 dvss.n2307 dvss.n2281 9.3005
R6870 dvss.n2495 dvss.n2494 9.3005
R6871 dvss.n2497 dvss.n2496 9.3005
R6872 dvss.n2499 dvss.n2277 9.3005
R6873 dvss.n2501 dvss.n2500 9.3005
R6874 dvss.n2480 dvss.n1 9.3005
R6875 dvss.n4407 dvss.n4406 9.3005
R6876 dvss.n4404 dvss.n0 9.3005
R6877 dvss.n4403 dvss.n4402 9.3005
R6878 dvss.n4401 dvss.n3 9.3005
R6879 dvss.n4400 dvss.n4399 9.3005
R6880 dvss.n4398 dvss.n4397 9.3005
R6881 dvss.n4396 dvss.n4395 9.3005
R6882 dvss.n4394 dvss.n6 9.3005
R6883 dvss.n4393 dvss.n4392 9.3005
R6884 dvss.n2460 dvss.n2459 9.3005
R6885 dvss.n2461 dvss.n2453 9.3005
R6886 dvss.n2463 dvss.n2462 9.3005
R6887 dvss.n2465 dvss.n2451 9.3005
R6888 dvss.n2469 dvss.n2468 9.3005
R6889 dvss.n2470 dvss.n2450 9.3005
R6890 dvss.n2472 dvss.n2471 9.3005
R6891 dvss.n2474 dvss.n2448 9.3005
R6892 dvss.n2478 dvss.n2477 9.3005
R6893 dvss.n2479 dvss.n2444 9.3005
R6894 dvss.n2483 dvss.n2482 9.3005
R6895 dvss.n2481 dvss.n2447 9.3005
R6896 dvss.n1062 dvss.n1060 8.56999
R6897 dvss.n2670 dvss.n2668 8.56999
R6898 dvss.n4121 dvss.n153 8.54791
R6899 dvss.n3865 dvss.n3779 8.54791
R6900 dvss.n3683 dvss.n3682 8.54791
R6901 dvss.n3570 dvss.n3569 8.54791
R6902 dvss.n3451 dvss.n3450 8.54791
R6903 dvss.n1734 dvss.n1596 8.54791
R6904 dvss.n1500 dvss.n1499 8.54791
R6905 dvss.n1214 dvss.n1212 8.54791
R6906 dvss.n1111 dvss.n1109 8.54791
R6907 dvss.n4356 dvss.n31 8.54791
R6908 dvss.n2061 dvss.n2036 8.54791
R6909 dvss.n3206 dvss.n3205 8.54791
R6910 dvss.n2876 dvss.n2875 8.54791
R6911 dvss.n2837 dvss.n2836 8.54791
R6912 dvss.n2798 dvss.n2797 8.54791
R6913 dvss.n2759 dvss.n2758 8.54791
R6914 dvss.n2720 dvss.n2719 8.54791
R6915 dvss.n2681 dvss.n2680 8.54791
R6916 dvss.n2188 dvss.n2187 8.54791
R6917 dvss.n821 dvss 8.48432
R6918 dvss.n2658 dvss 8.48432
R6919 dvss.n153 dvss 8.43944
R6920 dvss.n3779 dvss 8.43944
R6921 dvss.n3682 dvss 8.43944
R6922 dvss.n3569 dvss 8.43944
R6923 dvss.n3450 dvss 8.43944
R6924 dvss.n1596 dvss 8.43944
R6925 dvss.n1499 dvss 8.43944
R6926 dvss.n1212 dvss 8.43944
R6927 dvss.n1109 dvss 8.43944
R6928 dvss.n31 dvss 8.43944
R6929 dvss.n2036 dvss 8.43944
R6930 dvss.n3205 dvss 8.43944
R6931 dvss.n2875 dvss 8.43944
R6932 dvss.n2836 dvss 8.43944
R6933 dvss.n2797 dvss 8.43944
R6934 dvss.n2758 dvss 8.43944
R6935 dvss.n2719 dvss 8.43944
R6936 dvss.n2680 dvss 8.43944
R6937 dvss.n2187 dvss 8.43944
R6938 dvss.n2332 dvss.n2331 8.35606
R6939 dvss.n2300 dvss.n2283 8.35606
R6940 dvss.n2403 dvss.n2386 8.2416
R6941 dvss.n2331 dvss.n2330 8.0005
R6942 dvss.n2301 dvss.n2300 8.0005
R6943 dvss.n877 dvss.t265 7.99565
R6944 dvss.n2404 dvss.n2403 7.89091
R6945 dvss.n2467 dvss.n2450 7.5205
R6946 dvss.n1063 dvss.n1062 7.37677
R6947 dvss.n2671 dvss.n2670 7.37677
R6948 dvss.n4293 dvss.n4247 7.3244
R6949 dvss.n4301 dvss.n4300 7.25358
R6950 dvss.n2468 dvss.n2467 7.2005
R6951 dvss.n2485 dvss.n2484 7.2005
R6952 dvss.n2485 dvss.n2444 7.0405
R6953 dvss.n4207 dvss 6.4005
R6954 dvss.n131 dvss 6.4005
R6955 dvss.n3738 dvss 6.4005
R6956 dvss.n3627 dvss 6.4005
R6957 dvss.n3506 dvss 6.4005
R6958 dvss.n1628 dvss 6.4005
R6959 dvss.n1555 dvss 6.4005
R6960 dvss.n673 dvss 6.4005
R6961 dvss.n1168 dvss 6.4005
R6962 dvss.n3994 dvss 6.4005
R6963 dvss.n229 dvss 6.4005
R6964 dvss.n1914 dvss 6.4005
R6965 dvss.n1883 dvss 6.4005
R6966 dvss.n1852 dvss 6.4005
R6967 dvss.n475 dvss 6.4005
R6968 dvss.n1369 dvss 6.4005
R6969 dvss.n595 dvss 6.4005
R6970 dvss.n936 dvss 6.4005
R6971 dvss.n2133 dvss 6.4005
R6972 dvss.n2319 dvss.n2318 5.90523
R6973 dvss.n2289 dvss.n2287 5.90523
R6974 dvss.n2392 dvss.n2390 5.87299
R6975 dvss.n2456 dvss.n2454 5.65757
R6976 dvss.n2325 dvss.n2314 5.51161
R6977 dvss.n2298 dvss.n2297 5.51161
R6978 dvss.n4206 dvss 5.45235
R6979 dvss.n4142 dvss 5.45235
R6980 dvss.n3741 dvss 5.45235
R6981 dvss.n3630 dvss 5.45235
R6982 dvss.n3509 dvss 5.45235
R6983 dvss.n1706 dvss 5.45235
R6984 dvss.n1558 dvss 5.45235
R6985 dvss.n712 dvss 5.45235
R6986 dvss.n1171 dvss 5.45235
R6987 dvss.n4022 dvss 5.45235
R6988 dvss.n3943 dvss 5.45235
R6989 dvss.n3260 dvss 5.45235
R6990 dvss.n3310 dvss 5.45235
R6991 dvss.n3365 dvss 5.45235
R6992 dvss.n1812 dvss 5.45235
R6993 dvss.n1416 dvss 5.45235
R6994 dvss.n1329 dvss 5.45235
R6995 dvss.n935 dvss 5.45235
R6996 dvss.n2538 dvss 5.45235
R6997 dvss.n2401 dvss.n2400 5.43612
R6998 dvss.n2335 dvss.n2334 5.15606
R6999 dvss.n2306 dvss.n2305 5.15606
R7000 dvss.n1017 dvss.n1014 5.11678
R7001 dvss.n1016 dvss.n1015 5.11678
R7002 dvss.n2409 dvss.n2408 5.08543
R7003 dvss.n399 dvss.n398 4.96991
R7004 dvss.n457 dvss.n456 4.96991
R7005 dvss.n577 dvss.n576 4.96991
R7006 dvss.n518 dvss.n517 4.96991
R7007 dvss.n3356 dvss.n3355 4.96991
R7008 dvss.n1827 dvss.n1826 4.96991
R7009 dvss.n1407 dvss.n1406 4.96991
R7010 dvss.n1344 dvss.n1343 4.96991
R7011 dvss.n2465 dvss.n2464 4.9605
R7012 dvss dvss.n4390 4.88722
R7013 dvss.n2432 dvss 4.88201
R7014 dvss dvss.n2272 4.8781
R7015 dvss.n2513 dvss 4.8729
R7016 dvss.n4302 dvss.n4301 4.80519
R7017 dvss.n2473 dvss.n2472 4.6405
R7018 dvss.n4288 dvss.n4264 4.3437
R7019 dvss.n4294 dvss.n4293 4.25273
R7020 dvss.n4279 dvss.n4278 3.72777
R7021 dvss.n4215 dvss.n4214 3.68864
R7022 dvss.n4138 dvss.n4135 3.68864
R7023 dvss.n3764 dvss.n3763 3.68864
R7024 dvss.n3650 dvss.n3649 3.68864
R7025 dvss.n3533 dvss.n3532 3.68864
R7026 dvss.n1702 dvss.n453 3.68864
R7027 dvss.n1581 dvss.n1580 3.68864
R7028 dvss.n708 dvss.n573 3.68864
R7029 dvss.n1194 dvss.n1193 3.68864
R7030 dvss.n4331 dvss.n43 3.68864
R7031 dvss.n4370 dvss.n21 3.68864
R7032 dvss.n2075 dvss.n2003 3.68864
R7033 dvss.n3176 dvss.n3175 3.68864
R7034 dvss.n2862 dvss.n2861 3.68864
R7035 dvss.n2823 dvss.n2822 3.68864
R7036 dvss.n2784 dvss.n2783 3.68864
R7037 dvss.n2745 dvss.n2744 3.68864
R7038 dvss.n2706 dvss.n2705 3.68864
R7039 dvss.n2257 dvss.n2256 3.68864
R7040 dvss.n398 dvss 3.46403
R7041 dvss.n456 dvss 3.46403
R7042 dvss.n576 dvss 3.46403
R7043 dvss.n517 dvss 3.46403
R7044 dvss.n3355 dvss 3.46403
R7045 dvss.n1826 dvss 3.46403
R7046 dvss.n1406 dvss 3.46403
R7047 dvss.n1343 dvss 3.46403
R7048 dvss.n1060 dvss 3.25474
R7049 dvss.n2668 dvss 3.25474
R7050 dvss dvss.n2514 2.98292
R7051 dvss.n4390 dvss.n4389 2.94679
R7052 dvss.n4242 dvss 2.94111
R7053 dvss.n105 dvss.n103 2.87444
R7054 dvss.n4206 dvss.n4205 2.84494
R7055 dvss.n4142 dvss.n4141 2.84494
R7056 dvss.n3741 dvss.n3740 2.84494
R7057 dvss.n3630 dvss.n3629 2.84494
R7058 dvss.n3509 dvss.n3508 2.84494
R7059 dvss.n1706 dvss.n1705 2.84494
R7060 dvss.n1558 dvss.n1557 2.84494
R7061 dvss.n712 dvss.n711 2.84494
R7062 dvss.n1171 dvss.n1170 2.84494
R7063 dvss.n4022 dvss.n4021 2.84494
R7064 dvss.n3944 dvss.n3943 2.84494
R7065 dvss.n3260 dvss.n3259 2.84494
R7066 dvss.n3310 dvss.n3309 2.84494
R7067 dvss.n3365 dvss.n3364 2.84494
R7068 dvss.n1813 dvss.n1812 2.84494
R7069 dvss.n1416 dvss.n1415 2.84494
R7070 dvss.n1330 dvss.n1329 2.84494
R7071 dvss.n935 dvss.n934 2.84494
R7072 dvss.n2538 dvss.n2537 2.84494
R7073 dvss.n399 dvss 2.71109
R7074 dvss.n457 dvss 2.71109
R7075 dvss.n577 dvss 2.71109
R7076 dvss.n518 dvss 2.71109
R7077 dvss.n3356 dvss 2.71109
R7078 dvss.n1827 dvss 2.71109
R7079 dvss.n1407 dvss 2.71109
R7080 dvss.n1344 dvss 2.71109
R7081 dvss.n2323 dvss.n2322 2.66717
R7082 dvss.n2291 dvss.n2286 2.66717
R7083 dvss.n2394 dvss.n2389 2.63064
R7084 dvss.n4205 dvss 2.60791
R7085 dvss.n4141 dvss 2.60791
R7086 dvss.n3740 dvss 2.60791
R7087 dvss.n3629 dvss 2.60791
R7088 dvss.n3508 dvss 2.60791
R7089 dvss.n1705 dvss 2.60791
R7090 dvss.n1557 dvss 2.60791
R7091 dvss.n711 dvss 2.60791
R7092 dvss.n1170 dvss 2.60791
R7093 dvss.n4021 dvss 2.60791
R7094 dvss.n3944 dvss 2.60791
R7095 dvss.n3259 dvss 2.60791
R7096 dvss.n3309 dvss 2.60791
R7097 dvss.n3364 dvss 2.60791
R7098 dvss.n1813 dvss 2.60791
R7099 dvss.n1415 dvss 2.60791
R7100 dvss.n1330 dvss 2.60791
R7101 dvss.n934 dvss 2.60791
R7102 dvss.n2537 dvss 2.60791
R7103 dvss.n818 dvss 2.49542
R7104 dvss.n1030 dvss 2.49542
R7105 dvss.n869 dvss 2.49542
R7106 dvss.n857 dvss 2.49542
R7107 dvss.t115 dvss.t47 2.48392
R7108 dvss.n2434 dvss.n2433 2.43615
R7109 dvss.n2458 dvss.n2453 2.4005
R7110 dvss.n2362 dvss.n2311 2.31161
R7111 dvss.n2353 dvss.n2340 2.31161
R7112 dvss.n2494 dvss.n2280 2.31161
R7113 dvss.n2503 dvss.n2276 2.31161
R7114 dvss.n2413 dvss.n2383 2.27995
R7115 dvss.n2422 dvss.n2379 2.27995
R7116 dvss.n2374 dvss.n2372 2.17238
R7117 dvss.n2477 dvss.n2476 2.0805
R7118 dvss.n2446 dvss.n1 2.0805
R7119 dvss.n2514 dvss.n2513 1.87648
R7120 dvss.n4104 dvss 1.84457
R7121 dvss dvss.n4103 1.84457
R7122 dvss.n4103 dvss 1.84457
R7123 dvss.n3848 dvss 1.84457
R7124 dvss dvss.n3847 1.84457
R7125 dvss.n3847 dvss 1.84457
R7126 dvss.n3731 dvss 1.84457
R7127 dvss.n3710 dvss 1.84457
R7128 dvss.n3710 dvss 1.84457
R7129 dvss.n3615 dvss 1.84457
R7130 dvss.n3591 dvss 1.84457
R7131 dvss.n3591 dvss 1.84457
R7132 dvss.n3499 dvss 1.84457
R7133 dvss.n3478 dvss 1.84457
R7134 dvss.n3478 dvss 1.84457
R7135 dvss.n1717 dvss 1.84457
R7136 dvss dvss.n1716 1.84457
R7137 dvss.n1716 dvss 1.84457
R7138 dvss.n1548 dvss 1.84457
R7139 dvss.n1527 dvss 1.84457
R7140 dvss.n1527 dvss 1.84457
R7141 dvss.n1236 dvss 1.84457
R7142 dvss dvss.n1235 1.84457
R7143 dvss.n1235 dvss 1.84457
R7144 dvss.n1155 dvss 1.84457
R7145 dvss dvss.n1154 1.84457
R7146 dvss.n1154 dvss 1.84457
R7147 dvss.n4031 dvss 1.84457
R7148 dvss dvss.n4030 1.84457
R7149 dvss.n4030 dvss 1.84457
R7150 dvss.n3929 dvss 1.84457
R7151 dvss dvss.n3928 1.84457
R7152 dvss.n3928 dvss 1.84457
R7153 dvss.n3269 dvss 1.84457
R7154 dvss dvss.n3268 1.84457
R7155 dvss.n3268 dvss 1.84457
R7156 dvss.n3319 dvss 1.84457
R7157 dvss dvss.n3318 1.84457
R7158 dvss.n3318 dvss 1.84457
R7159 dvss.n3374 dvss 1.84457
R7160 dvss dvss.n3373 1.84457
R7161 dvss.n3373 dvss 1.84457
R7162 dvss.n1798 dvss 1.84457
R7163 dvss dvss.n1797 1.84457
R7164 dvss.n1797 dvss 1.84457
R7165 dvss.n1425 dvss 1.84457
R7166 dvss dvss.n1424 1.84457
R7167 dvss.n1424 dvss 1.84457
R7168 dvss.n1315 dvss 1.84457
R7169 dvss dvss.n1314 1.84457
R7170 dvss.n1314 dvss 1.84457
R7171 dvss.n923 dvss 1.84457
R7172 dvss dvss.n920 1.84457
R7173 dvss.n920 dvss 1.84457
R7174 dvss.n2547 dvss 1.84457
R7175 dvss dvss.n2546 1.84457
R7176 dvss.n2546 dvss 1.84457
R7177 dvss.n4284 dvss.n4270 1.72109
R7178 dvss.n4271 dvss.n4264 1.72109
R7179 dvss.n4302 dvss.n4242 1.5923
R7180 dvss.n2412 dvss.n2410 1.57858
R7181 dvss.n2514 dvss 1.47268
R7182 dvss.n2352 dvss.n2341 1.42272
R7183 dvss.n2505 dvss.n2504 1.42272
R7184 dvss.n2424 dvss.n2423 1.40324
R7185 dvss.n4253 dvss.n4244 1.35909
R7186 dvss.n4114 dvss.n163 1.34003
R7187 dvss.n4112 dvss.n165 1.34003
R7188 dvss.n4102 dvss.n165 1.34003
R7189 dvss.n3858 dvss.n3789 1.34003
R7190 dvss.n3856 dvss.n3791 1.34003
R7191 dvss.n3846 dvss.n3791 1.34003
R7192 dvss.n3692 dvss.n3691 1.34003
R7193 dvss.n3709 dvss.n3707 1.34003
R7194 dvss.n3711 dvss.n3709 1.34003
R7195 dvss.n3588 dvss.n368 1.34003
R7196 dvss.n3596 dvss.n3595 1.34003
R7197 dvss.n3595 dvss.n3594 1.34003
R7198 dvss.n3464 dvss.n3463 1.34003
R7199 dvss.n3477 dvss.n3475 1.34003
R7200 dvss.n3479 dvss.n3477 1.34003
R7201 dvss.n1727 dvss.n1606 1.34003
R7202 dvss.n1725 dvss.n1608 1.34003
R7203 dvss.n1715 dvss.n1608 1.34003
R7204 dvss.n1513 dvss.n1512 1.34003
R7205 dvss.n1526 dvss.n1524 1.34003
R7206 dvss.n1528 dvss.n1526 1.34003
R7207 dvss.n1227 dvss.n722 1.34003
R7208 dvss.n1232 dvss.n1230 1.34003
R7209 dvss.n1234 dvss.n1232 1.34003
R7210 dvss.n1132 dvss.n768 1.34003
R7211 dvss.n1134 dvss.n755 1.34003
R7212 dvss.n1153 dvss.n755 1.34003
R7213 dvss.n4048 dvss.n4047 1.34003
R7214 dvss.n4040 dvss.n4039 1.34003
R7215 dvss.n4039 dvss.n4038 1.34003
R7216 dvss.n3912 dvss.n246 1.34003
R7217 dvss.n3914 dvss.n237 1.34003
R7218 dvss.n3927 dvss.n237 1.34003
R7219 dvss.n3286 dvss.n3285 1.34003
R7220 dvss.n3278 dvss.n3277 1.34003
R7221 dvss.n3277 dvss.n3276 1.34003
R7222 dvss.n3336 dvss.n3335 1.34003
R7223 dvss.n3328 dvss.n3327 1.34003
R7224 dvss.n3327 dvss.n3326 1.34003
R7225 dvss.n3391 dvss.n3390 1.34003
R7226 dvss.n3383 dvss.n3382 1.34003
R7227 dvss.n3382 dvss.n3381 1.34003
R7228 dvss.n1781 dvss.n492 1.34003
R7229 dvss.n1783 dvss.n483 1.34003
R7230 dvss.n1796 dvss.n483 1.34003
R7231 dvss.n1442 dvss.n1441 1.34003
R7232 dvss.n1434 dvss.n1433 1.34003
R7233 dvss.n1433 dvss.n1432 1.34003
R7234 dvss.n1298 dvss.n612 1.34003
R7235 dvss.n1300 dvss.n603 1.34003
R7236 dvss.n1313 dvss.n603 1.34003
R7237 dvss.n911 dvss.n909 1.34003
R7238 dvss.n917 dvss.n915 1.34003
R7239 dvss.n919 dvss.n917 1.34003
R7240 dvss.n2564 dvss.n2563 1.34003
R7241 dvss.n2556 dvss.n2555 1.34003
R7242 dvss.n2555 dvss.n2554 1.34003
R7243 dvss.n4406 dvss.n4405 1.2805
R7244 dvss.n4398 dvss.n5 1.2805
R7245 dvss dvss.n4302 1.23235
R7246 dvss.n2433 dvss.n2432 1.16554
R7247 dvss.n2460 dvss.n2454 1.12105
R7248 dvss.n4294 dvss.n4244 1.09648
R7249 dvss.n2434 dvss.n2375 1.09487
R7250 dvss.n2396 dvss.n2390 1.05227
R7251 dvss.n2320 dvss.n2319 1.04213
R7252 dvss.n2293 dvss.n2287 1.04213
R7253 dvss.n4399 dvss.n4 0.9605
R7254 dvss.n2433 dvss.n2272 0.934094
R7255 dvss.n2435 dvss.n2434 0.886661
R7256 dvss.n4114 dvss 0.856314
R7257 dvss.n4113 dvss.n4112 0.856314
R7258 dvss dvss.n4102 0.856314
R7259 dvss.n3858 dvss 0.856314
R7260 dvss.n3857 dvss.n3856 0.856314
R7261 dvss dvss.n3846 0.856314
R7262 dvss.n3691 dvss 0.856314
R7263 dvss.n3707 dvss.n300 0.856314
R7264 dvss.n3711 dvss 0.856314
R7265 dvss dvss.n3588 0.856314
R7266 dvss.n3596 dvss.n3589 0.856314
R7267 dvss.n3594 dvss 0.856314
R7268 dvss.n3464 dvss 0.856314
R7269 dvss.n3475 dvss.n428 0.856314
R7270 dvss.n3479 dvss 0.856314
R7271 dvss.n1727 dvss 0.856314
R7272 dvss.n1726 dvss.n1725 0.856314
R7273 dvss dvss.n1715 0.856314
R7274 dvss.n1513 dvss 0.856314
R7275 dvss.n1524 dvss.n547 0.856314
R7276 dvss.n1528 dvss 0.856314
R7277 dvss dvss.n1227 0.856314
R7278 dvss.n1230 dvss.n1228 0.856314
R7279 dvss dvss.n1234 0.856314
R7280 dvss dvss.n1132 0.856314
R7281 dvss.n1134 dvss.n1133 0.856314
R7282 dvss dvss.n1153 0.856314
R7283 dvss.n4047 dvss 0.856314
R7284 dvss.n4040 dvss.n3968 0.856314
R7285 dvss.n4038 dvss 0.856314
R7286 dvss dvss.n3912 0.856314
R7287 dvss.n3914 dvss.n3913 0.856314
R7288 dvss dvss.n3927 0.856314
R7289 dvss.n3285 dvss 0.856314
R7290 dvss.n3278 dvss.n1904 0.856314
R7291 dvss.n3276 dvss 0.856314
R7292 dvss.n3335 dvss 0.856314
R7293 dvss.n3328 dvss.n1873 0.856314
R7294 dvss.n3326 dvss 0.856314
R7295 dvss.n3390 dvss 0.856314
R7296 dvss.n3383 dvss.n1842 0.856314
R7297 dvss.n3381 dvss 0.856314
R7298 dvss dvss.n1781 0.856314
R7299 dvss.n1783 dvss.n1782 0.856314
R7300 dvss dvss.n1796 0.856314
R7301 dvss.n1441 dvss 0.856314
R7302 dvss.n1434 dvss.n1359 0.856314
R7303 dvss.n1432 dvss 0.856314
R7304 dvss dvss.n1298 0.856314
R7305 dvss.n1300 dvss.n1299 0.856314
R7306 dvss dvss.n1313 0.856314
R7307 dvss dvss.n911 0.856314
R7308 dvss.n915 dvss.n912 0.856314
R7309 dvss dvss.n919 0.856314
R7310 dvss.n2563 dvss 0.856314
R7311 dvss.n2556 dvss.n2123 0.856314
R7312 dvss.n2554 dvss 0.856314
R7313 dvss.n2513 dvss.n2272 0.808117
R7314 dvss.n2375 dvss.n2368 0.7755
R7315 dvss.n2438 dvss.n2437 0.7755
R7316 dvss.n2363 dvss.n2309 0.711611
R7317 dvss.n2493 dvss.n2307 0.711611
R7318 dvss.n2436 dvss.n2435 0.705857
R7319 dvss.n4298 dvss.t171 0.627052
R7320 dvss.n4296 dvss.t170 0.627052
R7321 dvss.n4273 dvss.t573 0.627052
R7322 dvss.n4297 dvss.n4296 0.5805
R7323 dvss.n4299 dvss.n4298 0.5805
R7324 dvss.n4277 dvss.n4276 0.5805
R7325 dvss.n4276 dvss.n4275 0.5805
R7326 dvss.n4275 dvss.n4274 0.5805
R7327 dvss.n4274 dvss.n4273 0.5805
R7328 dvss.n4282 dvss.n4243 0.54848
R7329 dvss.n4242 dvss 0.543548
R7330 dvss.n2358 dvss.n2357 0.533833
R7331 dvss.n2499 dvss.n2498 0.533833
R7332 dvss.n2437 dvss.n2372 0.529518
R7333 dvss.n2418 dvss.n2417 0.526527
R7334 dvss.n4390 dvss 0.506359
R7335 dvss.n2484 dvss.n2483 0.4805
R7336 dvss.n4257 dvss.n4256 0.427268
R7337 dvss.n4260 dvss.n4247 0.312562
R7338 dvss.n4255 dvss.n4254 0.299742
R7339 dvss.n4300 dvss.n4297 0.279444
R7340 dvss.n4300 dvss.n4299 0.268206
R7341 dvss.n4261 dvss.n4260 0.254288
R7342 dvss.n2375 dvss.n2374 0.2505
R7343 dvss.n2432 dvss 0.187023
R7344 dvss.n4285 dvss.n4279 0.179346
R7345 dvss.n4283 dvss.n4282 0.179346
R7346 dvss.n4293 dvss.n4292 0.179346
R7347 dvss.n4262 dvss.n4261 0.179346
R7348 dvss.n2437 dvss.n2436 0.176839
R7349 dvss.n4247 dvss.n4246 0.174082
R7350 dvss.n4261 dvss.n4257 0.145702
R7351 dvss.n4282 dvss.n4281 0.129288
R7352 dvss.n2320 dvss.n2315 0.120292
R7353 dvss.n2327 dvss.n2315 0.120292
R7354 dvss.n2328 dvss.n2327 0.120292
R7355 dvss.n2329 dvss.n2328 0.120292
R7356 dvss.n2329 dvss.n2312 0.120292
R7357 dvss.n2336 dvss.n2312 0.120292
R7358 dvss.n2337 dvss.n2336 0.120292
R7359 dvss.n2361 dvss.n2337 0.120292
R7360 dvss.n2361 dvss.n2360 0.120292
R7361 dvss.n2360 dvss.n2338 0.120292
R7362 dvss.n2355 dvss.n2338 0.120292
R7363 dvss.n2355 dvss.n2354 0.120292
R7364 dvss.n2351 dvss.n2350 0.120292
R7365 dvss.n2350 dvss.n2342 0.120292
R7366 dvss.n2346 dvss.n2342 0.120292
R7367 dvss.n2346 dvss.n2345 0.120292
R7368 dvss.n2397 dvss.n2396 0.120292
R7369 dvss.n2398 dvss.n2397 0.120292
R7370 dvss.n2398 dvss.n2387 0.120292
R7371 dvss.n2405 dvss.n2387 0.120292
R7372 dvss.n2406 dvss.n2405 0.120292
R7373 dvss.n2407 dvss.n2406 0.120292
R7374 dvss.n2407 dvss.n2384 0.120292
R7375 dvss.n2414 dvss.n2384 0.120292
R7376 dvss.n2415 dvss.n2414 0.120292
R7377 dvss.n2415 dvss.n2380 0.120292
R7378 dvss.n2420 dvss.n2380 0.120292
R7379 dvss.n2421 dvss.n2420 0.120292
R7380 dvss.n2426 dvss.n2425 0.120292
R7381 dvss.n2427 dvss.n2426 0.120292
R7382 dvss.n2427 dvss.n2376 0.120292
R7383 dvss.n2431 dvss.n2376 0.120292
R7384 dvss.n2294 dvss.n2293 0.120292
R7385 dvss.n2295 dvss.n2294 0.120292
R7386 dvss.n2295 dvss.n2284 0.120292
R7387 dvss.n2302 dvss.n2284 0.120292
R7388 dvss.n2303 dvss.n2302 0.120292
R7389 dvss.n2304 dvss.n2303 0.120292
R7390 dvss.n2304 dvss.n2281 0.120292
R7391 dvss.n2495 dvss.n2281 0.120292
R7392 dvss.n2496 dvss.n2495 0.120292
R7393 dvss.n2496 dvss.n2277 0.120292
R7394 dvss.n2501 dvss.n2277 0.120292
R7395 dvss.n2502 dvss.n2501 0.120292
R7396 dvss.n2507 dvss.n2506 0.120292
R7397 dvss.n2508 dvss.n2507 0.120292
R7398 dvss.n2508 dvss.n2273 0.120292
R7399 dvss.n2512 dvss.n2273 0.120292
R7400 dvss.n2461 dvss.n2460 0.120292
R7401 dvss.n2462 dvss.n2461 0.120292
R7402 dvss.n2462 dvss.n2451 0.120292
R7403 dvss.n2469 dvss.n2451 0.120292
R7404 dvss.n2470 dvss.n2469 0.120292
R7405 dvss.n2471 dvss.n2470 0.120292
R7406 dvss.n2471 dvss.n2448 0.120292
R7407 dvss.n2478 dvss.n2448 0.120292
R7408 dvss.n2479 dvss.n2478 0.120292
R7409 dvss.n2482 dvss.n2479 0.120292
R7410 dvss.n2482 dvss.n2481 0.120292
R7411 dvss.n2481 dvss.n2480 0.120292
R7412 dvss.n4407 dvss.n0 0.120292
R7413 dvss.n4402 dvss.n0 0.120292
R7414 dvss.n4402 dvss.n4401 0.120292
R7415 dvss.n4401 dvss.n4400 0.120292
R7416 dvss.n4397 dvss.n4396 0.120292
R7417 dvss.n4396 dvss.n6 0.120292
R7418 dvss.n4392 dvss.n6 0.120292
R7419 dvss.n4392 dvss.n4391 0.120292
R7420 dvss.n4260 dvss.n4259 0.101043
R7421 dvss.n4254 dvss.n4253 0.100247
R7422 dvss.n4256 dvss.n4255 0.0989849
R7423 dvss.n4281 dvss.n4244 0.0888838
R7424 dvss.n4295 dvss.n4243 0.0808571
R7425 dvss.n2647 dvss 0.067223
R7426 dvss.n2648 dvss 0.067223
R7427 dvss.n2649 dvss 0.067223
R7428 dvss.n2650 dvss 0.067223
R7429 dvss.n2651 dvss 0.067223
R7430 dvss.n2652 dvss 0.067223
R7431 dvss.n2653 dvss 0.067223
R7432 dvss.n2654 dvss 0.067223
R7433 dvss.n2655 dvss 0.067223
R7434 dvss.n2656 dvss 0.067223
R7435 dvss.n2664 dvss 0.067223
R7436 dvss.n2665 dvss 0.067223
R7437 dvss.n2674 dvss 0.067223
R7438 dvss.n2676 dvss 0.067223
R7439 dvss.n2684 dvss 0.067223
R7440 dvss.n2685 dvss 0.067223
R7441 dvss.n2686 dvss 0.067223
R7442 dvss.n2687 dvss 0.067223
R7443 dvss.n2688 dvss 0.067223
R7444 dvss.n2689 dvss 0.067223
R7445 dvss.n2690 dvss 0.067223
R7446 dvss.n2693 dvss 0.067223
R7447 dvss.n2696 dvss 0.067223
R7448 dvss.n2697 dvss 0.067223
R7449 dvss.n2711 dvss 0.067223
R7450 dvss.n2712 dvss 0.067223
R7451 dvss.n2713 dvss 0.067223
R7452 dvss.n2715 dvss 0.067223
R7453 dvss.n2723 dvss 0.067223
R7454 dvss.n2724 dvss 0.067223
R7455 dvss.n2725 dvss 0.067223
R7456 dvss.n2726 dvss 0.067223
R7457 dvss.n2727 dvss 0.067223
R7458 dvss.n2728 dvss 0.067223
R7459 dvss.n2729 dvss 0.067223
R7460 dvss.n2732 dvss 0.067223
R7461 dvss.n2735 dvss 0.067223
R7462 dvss.n2736 dvss 0.067223
R7463 dvss.n2750 dvss 0.067223
R7464 dvss.n2751 dvss 0.067223
R7465 dvss.n2752 dvss 0.067223
R7466 dvss.n2754 dvss 0.067223
R7467 dvss.n2762 dvss 0.067223
R7468 dvss.n2763 dvss 0.067223
R7469 dvss.n2764 dvss 0.067223
R7470 dvss.n2765 dvss 0.067223
R7471 dvss.n2766 dvss 0.067223
R7472 dvss.n2767 dvss 0.067223
R7473 dvss.n2768 dvss 0.067223
R7474 dvss.n2771 dvss 0.067223
R7475 dvss.n2774 dvss 0.067223
R7476 dvss.n2775 dvss 0.067223
R7477 dvss.n2789 dvss 0.067223
R7478 dvss.n2790 dvss 0.067223
R7479 dvss.n2791 dvss 0.067223
R7480 dvss.n2793 dvss 0.067223
R7481 dvss.n2801 dvss 0.067223
R7482 dvss.n2802 dvss 0.067223
R7483 dvss.n2803 dvss 0.067223
R7484 dvss.n2804 dvss 0.067223
R7485 dvss.n2805 dvss 0.067223
R7486 dvss.n2806 dvss 0.067223
R7487 dvss.n2807 dvss 0.067223
R7488 dvss.n2810 dvss 0.067223
R7489 dvss.n2813 dvss 0.067223
R7490 dvss.n2814 dvss 0.067223
R7491 dvss.n2828 dvss 0.067223
R7492 dvss.n2829 dvss 0.067223
R7493 dvss.n2830 dvss 0.067223
R7494 dvss.n2832 dvss 0.067223
R7495 dvss.n2840 dvss 0.067223
R7496 dvss.n2841 dvss 0.067223
R7497 dvss.n2842 dvss 0.067223
R7498 dvss.n2843 dvss 0.067223
R7499 dvss.n2844 dvss 0.067223
R7500 dvss.n2845 dvss 0.067223
R7501 dvss.n2846 dvss 0.067223
R7502 dvss.n2849 dvss 0.067223
R7503 dvss.n2852 dvss 0.067223
R7504 dvss.n2853 dvss 0.067223
R7505 dvss.n2867 dvss 0.067223
R7506 dvss.n2868 dvss 0.067223
R7507 dvss.n2869 dvss 0.067223
R7508 dvss.n2871 dvss 0.067223
R7509 dvss.n2880 dvss 0.067223
R7510 dvss dvss.n2879 0.067223
R7511 dvss.n3147 dvss 0.067223
R7512 dvss.n3148 dvss 0.067223
R7513 dvss.n3150 dvss 0.067223
R7514 dvss dvss.n3149 0.067223
R7515 dvss.n3158 dvss 0.067223
R7516 dvss dvss.n3162 0.067223
R7517 dvss dvss.n2101 0.067223
R7518 dvss.n3181 dvss 0.067223
R7519 dvss.n3190 dvss 0.067223
R7520 dvss.n3191 dvss 0.067223
R7521 dvss.n3193 dvss 0.067223
R7522 dvss.n3202 dvss 0.067223
R7523 dvss dvss.n3208 0.067223
R7524 dvss.n3217 dvss 0.067223
R7525 dvss.n3218 dvss 0.067223
R7526 dvss.n3220 dvss 0.067223
R7527 dvss dvss.n3219 0.067223
R7528 dvss.n3229 dvss 0.067223
R7529 dvss.n3230 dvss 0.067223
R7530 dvss.n2016 dvss 0.067223
R7531 dvss dvss.n2021 0.067223
R7532 dvss dvss.n2020 0.067223
R7533 dvss.n2069 dvss 0.067223
R7534 dvss dvss.n2068 0.067223
R7535 dvss dvss.n2067 0.067223
R7536 dvss dvss.n2063 0.067223
R7537 dvss dvss.n4388 0.067223
R7538 dvss.n4385 dvss 0.067223
R7539 dvss dvss.n4384 0.067223
R7540 dvss dvss.n4383 0.067223
R7541 dvss.n4380 dvss 0.067223
R7542 dvss dvss.n4379 0.067223
R7543 dvss dvss.n4378 0.067223
R7544 dvss.n117 dvss 0.067223
R7545 dvss dvss.n111 0.067223
R7546 dvss dvss.n110 0.067223
R7547 dvss.n4364 dvss 0.067223
R7548 dvss dvss.n4363 0.067223
R7549 dvss dvss.n4362 0.067223
R7550 dvss dvss.n4358 0.067223
R7551 dvss.n4351 dvss 0.067223
R7552 dvss dvss.n4350 0.067223
R7553 dvss dvss.n4349 0.067223
R7554 dvss.n4346 dvss 0.067223
R7555 dvss dvss.n4345 0.067223
R7556 dvss dvss.n4344 0.067223
R7557 dvss.n4341 dvss 0.067223
R7558 dvss.n4333 dvss 0.067223
R7559 dvss.n4325 dvss 0.067223
R7560 dvss dvss.n4324 0.067223
R7561 dvss.n4317 dvss 0.067223
R7562 dvss dvss.n4316 0.067223
R7563 dvss dvss.n4315 0.067223
R7564 dvss.n2184 dvss 0.067223
R7565 dvss.n2192 dvss 0.067223
R7566 dvss dvss.n2191 0.067223
R7567 dvss.n2200 dvss 0.067223
R7568 dvss.n2201 dvss 0.067223
R7569 dvss.n2203 dvss 0.067223
R7570 dvss dvss.n2202 0.067223
R7571 dvss.n2239 dvss 0.067223
R7572 dvss dvss.n2243 0.067223
R7573 dvss dvss.n2157 0.067223
R7574 dvss.n2262 dvss 0.067223
R7575 dvss.n2270 dvss 0.067223
R7576 dvss.n2271 dvss 0.067223
R7577 dvss.n2515 dvss 0.067223
R7578 dvss dvss.n2570 0.067223
R7579 dvss dvss.n2569 0.067223
R7580 dvss.n2566 dvss 0.067223
R7581 dvss.n2558 dvss 0.067223
R7582 dvss.n2549 dvss 0.067223
R7583 dvss.n2541 dvss 0.067223
R7584 dvss dvss.n2540 0.067223
R7585 dvss.n2531 dvss 0.067223
R7586 dvss dvss.n2530 0.067223
R7587 dvss dvss.n2529 0.067223
R7588 dvss.n2526 dvss 0.067223
R7589 dvss dvss.n2525 0.067223
R7590 dvss dvss.n2524 0.067223
R7591 dvss dvss.n2548 0.0663784
R7592 dvss.n2704 dvss 0.0638446
R7593 dvss.n2743 dvss 0.0638446
R7594 dvss.n2782 dvss 0.0638446
R7595 dvss.n2821 dvss 0.0638446
R7596 dvss.n2860 dvss 0.0638446
R7597 dvss.n3174 dvss 0.0638446
R7598 dvss.n2017 dvss 0.0638446
R7599 dvss dvss.n116 0.0638446
R7600 dvss dvss.n4332 0.0638446
R7601 dvss.n2255 dvss 0.0638446
R7602 dvss.n2683 dvss 0.0613108
R7603 dvss.n2722 dvss 0.0613108
R7604 dvss.n2761 dvss 0.0613108
R7605 dvss.n2800 dvss 0.0613108
R7606 dvss.n2839 dvss 0.0613108
R7607 dvss.n2878 dvss 0.0613108
R7608 dvss.n3209 dvss 0.0613108
R7609 dvss dvss.n9 0.0613108
R7610 dvss dvss.n4354 0.0613108
R7611 dvss.n2190 dvss 0.0613108
R7612 dvss.n2351 dvss 0.0603958
R7613 dvss.n2425 dvss 0.0603958
R7614 dvss.n2506 dvss 0.0603958
R7615 dvss dvss.n4407 0.0603958
R7616 dvss.n4397 dvss 0.0603958
R7617 dvss dvss.n2561 0.0477973
R7618 dvss.n4299 dvss.t169 0.047052
R7619 dvss.n4298 dvss.t173 0.047052
R7620 dvss.n4296 dvss.t174 0.047052
R7621 dvss.n4297 dvss.t172 0.047052
R7622 dvss.n4273 dvss.t572 0.047052
R7623 dvss.n4274 dvss.t581 0.047052
R7624 dvss.n4275 dvss.t576 0.047052
R7625 dvss.n4276 dvss.t578 0.047052
R7626 dvss.n4277 dvss.t577 0.047052
R7627 dvss.n2662 dvss 0.0469527
R7628 dvss.n2709 dvss 0.0469527
R7629 dvss.n2748 dvss 0.0469527
R7630 dvss.n2787 dvss 0.0469527
R7631 dvss.n2826 dvss 0.0469527
R7632 dvss.n2865 dvss 0.0469527
R7633 dvss.n3178 dvss 0.0469527
R7634 dvss.n2073 dvss 0.0469527
R7635 dvss.n4368 dvss 0.0469527
R7636 dvss.n4321 dvss 0.0469527
R7637 dvss.n2259 dvss 0.0469527
R7638 dvss dvss.n2535 0.0469527
R7639 dvss dvss.n2557 0.0461081
R7640 dvss.n2545 dvss 0.0461081
R7641 dvss.n2700 dvss 0.0435743
R7642 dvss.n2702 dvss 0.0435743
R7643 dvss.n2739 dvss 0.0435743
R7644 dvss.n2741 dvss 0.0435743
R7645 dvss.n2778 dvss 0.0435743
R7646 dvss.n2780 dvss 0.0435743
R7647 dvss.n2817 dvss 0.0435743
R7648 dvss.n2819 dvss 0.0435743
R7649 dvss.n2856 dvss 0.0435743
R7650 dvss.n2858 dvss 0.0435743
R7651 dvss.n3159 dvss 0.0435743
R7652 dvss dvss.n2098 0.0435743
R7653 dvss.n3231 dvss 0.0435743
R7654 dvss.n2019 dvss 0.0435743
R7655 dvss.n4372 dvss 0.0435743
R7656 dvss dvss.n114 0.0435743
R7657 dvss dvss.n4340 0.0435743
R7658 dvss.n4329 dvss 0.0435743
R7659 dvss.n2240 dvss 0.0435743
R7660 dvss dvss.n2154 0.0435743
R7661 dvss.n2135 dvss 0.0418851
R7662 dvss.n2675 dvss 0.0410405
R7663 dvss dvss.n2677 0.0410405
R7664 dvss.n2714 dvss 0.0410405
R7665 dvss dvss.n2716 0.0410405
R7666 dvss.n2753 dvss 0.0410405
R7667 dvss dvss.n2755 0.0410405
R7668 dvss.n2792 dvss 0.0410405
R7669 dvss dvss.n2794 0.0410405
R7670 dvss.n2831 dvss 0.0410405
R7671 dvss dvss.n2833 0.0410405
R7672 dvss.n2870 dvss 0.0410405
R7673 dvss dvss.n2872 0.0410405
R7674 dvss dvss.n3192 0.0410405
R7675 dvss dvss.n2086 0.0410405
R7676 dvss.n2064 dvss 0.0410405
R7677 dvss.n2059 dvss 0.0410405
R7678 dvss.n4359 dvss 0.0410405
R7679 dvss.n32 dvss 0.0410405
R7680 dvss dvss.n2174 0.0410405
R7681 dvss.n2667 dvss 0.0385068
R7682 dvss.n4295 dvss.n4294 0.0362143
R7683 dvss.n2673 dvss 0.0351284
R7684 dvss.n841 dvss 0.0323548
R7685 dvss.n842 dvss 0.0323548
R7686 dvss.n847 dvss 0.0323548
R7687 dvss.n848 dvss 0.0323548
R7688 dvss.n849 dvss 0.0323548
R7689 dvss.n850 dvss 0.0323548
R7690 dvss.n860 dvss 0.0323548
R7691 dvss.n861 dvss 0.0323548
R7692 dvss.n872 dvss 0.0323548
R7693 dvss.n873 dvss 0.0323548
R7694 dvss.n885 dvss 0.0323548
R7695 dvss.n887 dvss 0.0323548
R7696 dvss.n891 dvss 0.0323548
R7697 dvss.n892 dvss 0.0323548
R7698 dvss.n913 dvss 0.0323548
R7699 dvss.n901 dvss 0.0323548
R7700 dvss.n926 dvss 0.0323548
R7701 dvss.n927 dvss 0.0323548
R7702 dvss.n940 dvss 0.0323548
R7703 dvss dvss.n939 0.0323548
R7704 dvss.n1272 dvss 0.0323548
R7705 dvss.n1273 dvss 0.0323548
R7706 dvss.n1275 dvss 0.0323548
R7707 dvss dvss.n1274 0.0323548
R7708 dvss.n1284 dvss 0.0323548
R7709 dvss.n1287 dvss 0.0323548
R7710 dvss dvss.n1286 0.0323548
R7711 dvss.n1302 dvss 0.0323548
R7712 dvss dvss.n604 0.0323548
R7713 dvss.n1326 dvss 0.0323548
R7714 dvss.n1327 dvss 0.0323548
R7715 dvss.n1340 dvss 0.0323548
R7716 dvss.n1455 dvss 0.0323548
R7717 dvss dvss.n1454 0.0323548
R7718 dvss dvss.n1453 0.0323548
R7719 dvss.n1450 dvss 0.0323548
R7720 dvss dvss.n1448 0.0323548
R7721 dvss.n1445 dvss 0.0323548
R7722 dvss dvss.n1444 0.0323548
R7723 dvss.n1436 dvss 0.0323548
R7724 dvss.n1427 dvss 0.0323548
R7725 dvss.n1419 dvss 0.0323548
R7726 dvss dvss.n1418 0.0323548
R7727 dvss.n1409 dvss 0.0323548
R7728 dvss.n1755 dvss 0.0323548
R7729 dvss.n1756 dvss 0.0323548
R7730 dvss.n1758 dvss 0.0323548
R7731 dvss dvss.n1757 0.0323548
R7732 dvss.n1767 dvss 0.0323548
R7733 dvss.n1770 dvss 0.0323548
R7734 dvss dvss.n1769 0.0323548
R7735 dvss.n1785 dvss 0.0323548
R7736 dvss dvss.n484 0.0323548
R7737 dvss.n1809 dvss 0.0323548
R7738 dvss.n1810 dvss 0.0323548
R7739 dvss.n1823 dvss 0.0323548
R7740 dvss.n3404 dvss 0.0323548
R7741 dvss dvss.n3403 0.0323548
R7742 dvss dvss.n3402 0.0323548
R7743 dvss.n3399 dvss 0.0323548
R7744 dvss dvss.n3397 0.0323548
R7745 dvss.n3394 dvss 0.0323548
R7746 dvss dvss.n3393 0.0323548
R7747 dvss.n3385 dvss 0.0323548
R7748 dvss.n3376 dvss 0.0323548
R7749 dvss.n3368 dvss 0.0323548
R7750 dvss dvss.n3367 0.0323548
R7751 dvss.n3358 dvss 0.0323548
R7752 dvss dvss.n3351 0.0323548
R7753 dvss.n3348 dvss 0.0323548
R7754 dvss dvss.n3347 0.0323548
R7755 dvss dvss.n3346 0.0323548
R7756 dvss dvss.n3342 0.0323548
R7757 dvss dvss.n3341 0.0323548
R7758 dvss.n3338 dvss 0.0323548
R7759 dvss.n3330 dvss 0.0323548
R7760 dvss.n3321 dvss 0.0323548
R7761 dvss.n3313 dvss 0.0323548
R7762 dvss dvss.n3312 0.0323548
R7763 dvss.n3303 dvss 0.0323548
R7764 dvss dvss.n3302 0.0323548
R7765 dvss dvss.n3301 0.0323548
R7766 dvss.n3298 dvss 0.0323548
R7767 dvss dvss.n3297 0.0323548
R7768 dvss dvss.n3296 0.0323548
R7769 dvss dvss.n3292 0.0323548
R7770 dvss dvss.n3291 0.0323548
R7771 dvss.n3288 dvss 0.0323548
R7772 dvss.n3280 dvss 0.0323548
R7773 dvss.n3271 dvss 0.0323548
R7774 dvss.n3263 dvss 0.0323548
R7775 dvss dvss.n3262 0.0323548
R7776 dvss.n3253 dvss 0.0323548
R7777 dvss dvss.n3252 0.0323548
R7778 dvss.n3886 dvss 0.0323548
R7779 dvss.n3887 dvss 0.0323548
R7780 dvss.n3889 dvss 0.0323548
R7781 dvss dvss.n3888 0.0323548
R7782 dvss.n3898 dvss 0.0323548
R7783 dvss.n3901 dvss 0.0323548
R7784 dvss dvss.n3900 0.0323548
R7785 dvss.n3916 dvss 0.0323548
R7786 dvss dvss.n238 0.0323548
R7787 dvss.n3940 dvss 0.0323548
R7788 dvss.n3941 dvss 0.0323548
R7789 dvss.n3954 dvss 0.0323548
R7790 dvss.n3955 dvss 0.0323548
R7791 dvss.n4061 dvss 0.0323548
R7792 dvss dvss.n4060 0.0323548
R7793 dvss dvss.n4059 0.0323548
R7794 dvss.n4056 dvss 0.0323548
R7795 dvss dvss.n4054 0.0323548
R7796 dvss.n4051 dvss 0.0323548
R7797 dvss dvss.n4050 0.0323548
R7798 dvss.n4042 dvss 0.0323548
R7799 dvss.n4033 dvss 0.0323548
R7800 dvss.n4025 dvss 0.0323548
R7801 dvss dvss.n4024 0.0323548
R7802 dvss.n4015 dvss 0.0323548
R7803 dvss dvss.n4014 0.0323548
R7804 dvss dvss.n4013 0.0323548
R7805 dvss.n4306 dvss 0.0323548
R7806 dvss dvss.n4305 0.0323548
R7807 dvss dvss.n4304 0.0323548
R7808 dvss.n922 dvss 0.0319516
R7809 dvss dvss.n600 0.0319516
R7810 dvss dvss.n1426 0.0319516
R7811 dvss dvss.n480 0.0319516
R7812 dvss dvss.n3375 0.0319516
R7813 dvss dvss.n3320 0.0319516
R7814 dvss dvss.n3270 0.0319516
R7815 dvss dvss.n234 0.0319516
R7816 dvss dvss.n4032 0.0319516
R7817 dvss.n1408 dvss.n1403 0.0311452
R7818 dvss.n1829 dvss.n1828 0.0311452
R7819 dvss.n3357 dvss.n3352 0.0311452
R7820 dvss dvss.n2692 0.0300608
R7821 dvss dvss.n2731 0.0300608
R7822 dvss dvss.n2770 0.0300608
R7823 dvss dvss.n2809 0.0300608
R7824 dvss dvss.n2848 0.0300608
R7825 dvss.n3163 dvss 0.0300608
R7826 dvss.n2011 dvss 0.0300608
R7827 dvss.n109 dvss 0.0300608
R7828 dvss dvss.n4336 0.0300608
R7829 dvss.n2244 dvss 0.0300608
R7830 dvss.n1346 dvss.n1345 0.0295323
R7831 dvss.n4272 dvss.n4271 0.029472
R7832 dvss.n4284 dvss.n4280 0.029472
R7833 dvss.n856 dvss 0.0287258
R7834 dvss.n1113 dvss 0.0282388
R7835 dvss.n1136 dvss 0.0282388
R7836 dvss.n1142 dvss 0.0282388
R7837 dvss dvss.n1173 0.0282388
R7838 dvss dvss.n1187 0.0282388
R7839 dvss.n1198 dvss 0.0282388
R7840 dvss.n632 dvss 0.0282388
R7841 dvss.n633 dvss 0.0282388
R7842 dvss.n1207 dvss 0.0282388
R7843 dvss.n1216 dvss 0.0282388
R7844 dvss dvss.n651 0.0282388
R7845 dvss.n1238 dvss 0.0282388
R7846 dvss dvss.n714 0.0282388
R7847 dvss.n701 dvss 0.0282388
R7848 dvss dvss.n569 0.0282388
R7849 dvss.n1486 dvss 0.0282388
R7850 dvss.n1483 dvss 0.0282388
R7851 dvss.n1496 dvss 0.0282388
R7852 dvss.n1522 dvss 0.0282388
R7853 dvss dvss.n1533 0.0282388
R7854 dvss dvss.n1560 0.0282388
R7855 dvss dvss.n1574 0.0282388
R7856 dvss.n1742 dvss 0.0282388
R7857 dvss dvss.n1741 0.0282388
R7858 dvss dvss.n1740 0.0282388
R7859 dvss dvss.n1736 0.0282388
R7860 dvss.n1668 dvss 0.0282388
R7861 dvss dvss.n1719 0.0282388
R7862 dvss dvss.n1708 0.0282388
R7863 dvss.n1695 dvss 0.0282388
R7864 dvss.n3438 dvss 0.0282388
R7865 dvss.n3435 dvss 0.0282388
R7866 dvss dvss.n3434 0.0282388
R7867 dvss.n3447 dvss 0.0282388
R7868 dvss.n3473 dvss 0.0282388
R7869 dvss dvss.n3484 0.0282388
R7870 dvss dvss.n3511 0.0282388
R7871 dvss dvss.n3526 0.0282388
R7872 dvss dvss.n393 0.0282388
R7873 dvss.n3558 dvss 0.0282388
R7874 dvss.n3555 dvss 0.0282388
R7875 dvss.n3566 dvss 0.0282388
R7876 dvss.n3598 dvss 0.0282388
R7877 dvss.n3610 dvss 0.0282388
R7878 dvss.n3632 dvss 0.0282388
R7879 dvss dvss.n3643 0.0282388
R7880 dvss.n3653 dvss 0.0282388
R7881 dvss dvss.n3656 0.0282388
R7882 dvss.n3671 dvss 0.0282388
R7883 dvss dvss.n3670 0.0282388
R7884 dvss.n3679 dvss 0.0282388
R7885 dvss.n3705 dvss 0.0282388
R7886 dvss dvss.n3713 0.0282388
R7887 dvss dvss.n3743 0.0282388
R7888 dvss dvss.n3757 0.0282388
R7889 dvss.n3767 dvss 0.0282388
R7890 dvss.n3873 dvss 0.0282388
R7891 dvss dvss.n3872 0.0282388
R7892 dvss dvss.n3871 0.0282388
R7893 dvss dvss.n3867 0.0282388
R7894 dvss.n3806 dvss 0.0282388
R7895 dvss dvss.n3850 0.0282388
R7896 dvss dvss.n4144 0.0282388
R7897 dvss.n211 dvss 0.0282388
R7898 dvss.n212 dvss 0.0282388
R7899 dvss.n4129 dvss 0.0282388
R7900 dvss dvss.n4128 0.0282388
R7901 dvss dvss.n4127 0.0282388
R7902 dvss dvss.n4123 0.0282388
R7903 dvss.n4084 dvss 0.0282388
R7904 dvss dvss.n4106 0.0282388
R7905 dvss.n4202 dvss 0.0282388
R7906 dvss.n4219 dvss 0.0282388
R7907 dvss dvss.n4218 0.0282388
R7908 dvss.n4233 dvss 0.0282388
R7909 dvss.n4234 dvss 0.0282388
R7910 dvss.n4241 dvss 0.0282388
R7911 dvss.n1021 dvss 0.0278876
R7912 dvss.n1023 dvss 0.0278876
R7913 dvss.n1024 dvss 0.0278876
R7914 dvss.n1025 dvss 0.0278876
R7915 dvss.n1026 dvss 0.0278876
R7916 dvss.n1027 dvss 0.0278876
R7917 dvss.n1033 dvss 0.0278876
R7918 dvss.n1034 dvss 0.0278876
R7919 dvss.n1056 dvss 0.0278876
R7920 dvss dvss.n1069 0.0278876
R7921 dvss.n787 dvss 0.0278876
R7922 dvss dvss.n753 0.0278876
R7923 dvss dvss.n1237 0.0278876
R7924 dvss.n1547 dvss 0.0278876
R7925 dvss dvss.n1718 0.0278876
R7926 dvss.n3498 dvss 0.0278876
R7927 dvss.n3614 dvss 0.0278876
R7928 dvss.n3730 dvss 0.0278876
R7929 dvss dvss.n3849 0.0278876
R7930 dvss dvss.n4105 0.0278876
R7931 dvss.n2119 dvss 0.027527
R7932 dvss dvss.n2552 0.027527
R7933 dvss.n1464 dvss.n578 0.0271854
R7934 dvss.n1584 dvss.n519 0.0271854
R7935 dvss.n3413 dvss.n458 0.0271854
R7936 dvss.n3536 dvss.n400 0.0271854
R7937 dvss dvss.n2565 0.0258378
R7938 dvss.n2553 dvss 0.0258378
R7939 dvss.n1121 dvss 0.0257809
R7940 dvss dvss.n643 0.0257809
R7941 dvss.n1502 dvss 0.0257809
R7942 dvss dvss.n1732 0.0257809
R7943 dvss.n3453 dvss 0.0257809
R7944 dvss.n3575 dvss 0.0257809
R7945 dvss.n3694 dvss 0.0257809
R7946 dvss dvss.n3863 0.0257809
R7947 dvss dvss.n4119 0.0257809
R7948 dvss.n1029 dvss 0.0247275
R7949 dvss.n2698 dvss 0.0233041
R7950 dvss.n2737 dvss 0.0233041
R7951 dvss.n2776 dvss 0.0233041
R7952 dvss.n2815 dvss 0.0233041
R7953 dvss.n2854 dvss 0.0233041
R7954 dvss.n3161 dvss 0.0233041
R7955 dvss dvss.n3233 0.0233041
R7956 dvss dvss.n4374 0.0233041
R7957 dvss.n4337 dvss 0.0233041
R7958 dvss.n2242 dvss 0.0233041
R7959 dvss dvss.n894 0.0230806
R7960 dvss dvss.n1296 0.0230806
R7961 dvss dvss.n1439 0.0230806
R7962 dvss dvss.n1779 0.0230806
R7963 dvss dvss.n3388 0.0230806
R7964 dvss dvss.n3333 0.0230806
R7965 dvss dvss.n3283 0.0230806
R7966 dvss dvss.n3910 0.0230806
R7967 dvss dvss.n4045 0.0230806
R7968 dvss.n870 dvss 0.0226774
R7969 dvss.n937 dvss 0.0226774
R7970 dvss.n594 dvss 0.0226774
R7971 dvss dvss.n1413 0.0226774
R7972 dvss.n474 dvss 0.0226774
R7973 dvss dvss.n3362 0.0226774
R7974 dvss dvss.n3307 0.0226774
R7975 dvss dvss.n3257 0.0226774
R7976 dvss.n228 dvss 0.0226774
R7977 dvss dvss.n4019 0.0226774
R7978 dvss.n2354 dvss 0.0226354
R7979 dvss.n2345 dvss 0.0226354
R7980 dvss.n2421 dvss 0.0226354
R7981 dvss dvss.n2431 0.0226354
R7982 dvss.n2502 dvss 0.0226354
R7983 dvss dvss.n2512 0.0226354
R7984 dvss.n2480 dvss 0.0226354
R7985 dvss.n4400 dvss 0.0226354
R7986 dvss.n4391 dvss 0.0226354
R7987 dvss.n914 dvss 0.0222742
R7988 dvss.n924 dvss 0.0222742
R7989 dvss dvss.n1301 0.0222742
R7990 dvss dvss.n1316 0.0222742
R7991 dvss dvss.n1435 0.0222742
R7992 dvss.n1423 dvss 0.0222742
R7993 dvss dvss.n1784 0.0222742
R7994 dvss dvss.n1799 0.0222742
R7995 dvss dvss.n3384 0.0222742
R7996 dvss.n3372 dvss 0.0222742
R7997 dvss dvss.n3329 0.0222742
R7998 dvss.n3317 dvss 0.0222742
R7999 dvss dvss.n3279 0.0222742
R8000 dvss.n3267 dvss 0.0222742
R8001 dvss dvss.n3915 0.0222742
R8002 dvss dvss.n3930 0.0222742
R8003 dvss dvss.n4041 0.0222742
R8004 dvss.n4029 dvss 0.0222742
R8005 dvss dvss.n928 0.0202581
R8006 dvss.n1332 dvss 0.0202581
R8007 dvss.n1371 dvss 0.0202581
R8008 dvss.n1815 dvss 0.0202581
R8009 dvss.n1854 dvss 0.0202581
R8010 dvss.n1885 dvss 0.0202581
R8011 dvss.n1916 dvss 0.0202581
R8012 dvss.n3946 dvss 0.0202581
R8013 dvss.n3996 dvss 0.0202581
R8014 dvss dvss.n1130 0.0201629
R8015 dvss dvss.n1225 0.0201629
R8016 dvss.n1515 dvss 0.0201629
R8017 dvss.n1667 dvss 0.0201629
R8018 dvss.n3466 dvss 0.0201629
R8019 dvss dvss.n3586 0.0201629
R8020 dvss.n3704 dvss 0.0201629
R8021 dvss.n3805 dvss 0.0201629
R8022 dvss.n4083 dvss 0.0201629
R8023 dvss.n1283 dvss 0.0198548
R8024 dvss dvss.n1449 0.0198548
R8025 dvss.n1766 dvss 0.0198548
R8026 dvss dvss.n3398 0.0198548
R8027 dvss.n3343 dvss 0.0198548
R8028 dvss.n3293 dvss 0.0198548
R8029 dvss.n3897 dvss 0.0198548
R8030 dvss dvss.n4055 0.0198548
R8031 dvss.n1195 dvss 0.0198118
R8032 dvss.n1467 dvss 0.0198118
R8033 dvss dvss.n512 0.0198118
R8034 dvss.n3416 dvss 0.0198118
R8035 dvss dvss.n392 0.0198118
R8036 dvss dvss.n330 0.0198118
R8037 dvss dvss.n267 0.0198118
R8038 dvss.n4133 dvss 0.0198118
R8039 dvss dvss.n73 0.0198118
R8040 dvss dvss.n1135 0.0194607
R8041 dvss.n1229 dvss 0.0194607
R8042 dvss.n1523 dvss 0.0194607
R8043 dvss.n1724 dvss 0.0194607
R8044 dvss.n3474 dvss 0.0194607
R8045 dvss dvss.n3597 0.0194607
R8046 dvss.n3706 dvss 0.0194607
R8047 dvss.n3855 dvss 0.0194607
R8048 dvss.n4111 dvss 0.0194607
R8049 dvss.n886 dvss 0.0194516
R8050 dvss.n858 dvss 0.0190484
R8051 dvss.n881 dvss 0.0186452
R8052 dvss dvss.n1157 0.0184073
R8053 dvss.n663 dvss 0.0184073
R8054 dvss dvss.n538 0.0184073
R8055 dvss.n1617 dvss 0.0184073
R8056 dvss dvss.n419 0.0184073
R8057 dvss dvss.n354 0.0184073
R8058 dvss dvss.n288 0.0184073
R8059 dvss.n3843 dvss 0.0184073
R8060 dvss.n4099 dvss 0.0184073
R8061 dvss.n2672 dvss 0.0182365
R8062 dvss dvss.n774 0.0173539
R8063 dvss.n1210 dvss 0.0173539
R8064 dvss dvss.n642 0.0173539
R8065 dvss dvss.n1482 0.0173539
R8066 dvss dvss.n558 0.0173539
R8067 dvss.n1737 dvss 0.0173539
R8068 dvss.n1597 dvss 0.0173539
R8069 dvss dvss.n3433 0.0173539
R8070 dvss dvss.n439 0.0173539
R8071 dvss dvss.n3554 0.0173539
R8072 dvss.n3572 dvss 0.0173539
R8073 dvss dvss.n3669 0.0173539
R8074 dvss.n3685 dvss 0.0173539
R8075 dvss.n3868 dvss 0.0173539
R8076 dvss.n3780 dvss 0.0173539
R8077 dvss.n4124 dvss 0.0173539
R8078 dvss.n154 dvss 0.0173539
R8079 dvss.n884 dvss 0.0170323
R8080 dvss.n1107 dvss 0.0170028
R8081 dvss dvss.n815 0.0166517
R8082 dvss.n1031 dvss 0.0163006
R8083 dvss.n1192 dvss 0.0163006
R8084 dvss dvss.n733 0.0163006
R8085 dvss.n707 dvss 0.0163006
R8086 dvss dvss.n709 0.0163006
R8087 dvss.n1579 dvss 0.0163006
R8088 dvss dvss.n522 0.0163006
R8089 dvss.n1701 dvss 0.0163006
R8090 dvss dvss.n1703 0.0163006
R8091 dvss.n3531 dvss 0.0163006
R8092 dvss dvss.n403 0.0163006
R8093 dvss.n3648 dvss 0.0163006
R8094 dvss dvss.n335 0.0163006
R8095 dvss.n3762 dvss 0.0163006
R8096 dvss dvss.n272 0.0163006
R8097 dvss.n4137 dvss 0.0163006
R8098 dvss dvss.n4139 0.0163006
R8099 dvss.n4213 dvss 0.0163006
R8100 dvss dvss.n87 0.0163006
R8101 dvss dvss.n1067 0.0159494
R8102 dvss dvss.n2647 0.0148581
R8103 dvss dvss.n2648 0.0148581
R8104 dvss dvss.n2649 0.0148581
R8105 dvss dvss.n2650 0.0148581
R8106 dvss dvss.n2651 0.0148581
R8107 dvss dvss.n2652 0.0148581
R8108 dvss dvss.n2653 0.0148581
R8109 dvss dvss.n2654 0.0148581
R8110 dvss dvss.n2655 0.0148581
R8111 dvss dvss.n2656 0.0148581
R8112 dvss.n2657 dvss 0.0148581
R8113 dvss dvss.n2664 0.0148581
R8114 dvss dvss.n2665 0.0148581
R8115 dvss.n2667 dvss 0.0148581
R8116 dvss dvss.n2666 0.0148581
R8117 dvss dvss.n2666 0.0148581
R8118 dvss dvss.n2672 0.0148581
R8119 dvss dvss.n2673 0.0148581
R8120 dvss dvss.n2674 0.0148581
R8121 dvss dvss.n2675 0.0148581
R8122 dvss dvss.n2676 0.0148581
R8123 dvss.n2678 dvss 0.0148581
R8124 dvss dvss.n2683 0.0148581
R8125 dvss dvss.n2684 0.0148581
R8126 dvss dvss.n2685 0.0148581
R8127 dvss dvss.n2686 0.0148581
R8128 dvss dvss.n2687 0.0148581
R8129 dvss dvss.n2688 0.0148581
R8130 dvss dvss.n2689 0.0148581
R8131 dvss dvss.n2690 0.0148581
R8132 dvss.n2700 dvss 0.0148581
R8133 dvss dvss.n2691 0.0148581
R8134 dvss.n2698 dvss 0.0148581
R8135 dvss dvss.n2692 0.0148581
R8136 dvss dvss.n2693 0.0148581
R8137 dvss.n2702 dvss 0.0148581
R8138 dvss dvss.n2695 0.0148581
R8139 dvss dvss.n2696 0.0148581
R8140 dvss dvss.n2697 0.0148581
R8141 dvss.n2707 dvss 0.0148581
R8142 dvss dvss.n2711 0.0148581
R8143 dvss dvss.n2712 0.0148581
R8144 dvss dvss.n2713 0.0148581
R8145 dvss dvss.n2714 0.0148581
R8146 dvss dvss.n2715 0.0148581
R8147 dvss.n2717 dvss 0.0148581
R8148 dvss dvss.n2722 0.0148581
R8149 dvss dvss.n2723 0.0148581
R8150 dvss dvss.n2724 0.0148581
R8151 dvss dvss.n2725 0.0148581
R8152 dvss dvss.n2726 0.0148581
R8153 dvss dvss.n2727 0.0148581
R8154 dvss dvss.n2728 0.0148581
R8155 dvss dvss.n2729 0.0148581
R8156 dvss.n2739 dvss 0.0148581
R8157 dvss dvss.n2730 0.0148581
R8158 dvss.n2737 dvss 0.0148581
R8159 dvss dvss.n2731 0.0148581
R8160 dvss dvss.n2732 0.0148581
R8161 dvss.n2741 dvss 0.0148581
R8162 dvss dvss.n2734 0.0148581
R8163 dvss dvss.n2735 0.0148581
R8164 dvss dvss.n2736 0.0148581
R8165 dvss.n2746 dvss 0.0148581
R8166 dvss dvss.n2750 0.0148581
R8167 dvss dvss.n2751 0.0148581
R8168 dvss dvss.n2752 0.0148581
R8169 dvss dvss.n2753 0.0148581
R8170 dvss dvss.n2754 0.0148581
R8171 dvss.n2756 dvss 0.0148581
R8172 dvss dvss.n2761 0.0148581
R8173 dvss dvss.n2762 0.0148581
R8174 dvss dvss.n2763 0.0148581
R8175 dvss dvss.n2764 0.0148581
R8176 dvss dvss.n2765 0.0148581
R8177 dvss dvss.n2766 0.0148581
R8178 dvss dvss.n2767 0.0148581
R8179 dvss dvss.n2768 0.0148581
R8180 dvss.n2778 dvss 0.0148581
R8181 dvss dvss.n2769 0.0148581
R8182 dvss.n2776 dvss 0.0148581
R8183 dvss dvss.n2770 0.0148581
R8184 dvss dvss.n2771 0.0148581
R8185 dvss.n2780 dvss 0.0148581
R8186 dvss dvss.n2773 0.0148581
R8187 dvss dvss.n2774 0.0148581
R8188 dvss dvss.n2775 0.0148581
R8189 dvss.n2785 dvss 0.0148581
R8190 dvss dvss.n2789 0.0148581
R8191 dvss dvss.n2790 0.0148581
R8192 dvss dvss.n2791 0.0148581
R8193 dvss dvss.n2792 0.0148581
R8194 dvss dvss.n2793 0.0148581
R8195 dvss.n2795 dvss 0.0148581
R8196 dvss dvss.n2800 0.0148581
R8197 dvss dvss.n2801 0.0148581
R8198 dvss dvss.n2802 0.0148581
R8199 dvss dvss.n2803 0.0148581
R8200 dvss dvss.n2804 0.0148581
R8201 dvss dvss.n2805 0.0148581
R8202 dvss dvss.n2806 0.0148581
R8203 dvss dvss.n2807 0.0148581
R8204 dvss.n2817 dvss 0.0148581
R8205 dvss dvss.n2808 0.0148581
R8206 dvss.n2815 dvss 0.0148581
R8207 dvss dvss.n2809 0.0148581
R8208 dvss dvss.n2810 0.0148581
R8209 dvss.n2819 dvss 0.0148581
R8210 dvss dvss.n2812 0.0148581
R8211 dvss dvss.n2813 0.0148581
R8212 dvss dvss.n2814 0.0148581
R8213 dvss.n2824 dvss 0.0148581
R8214 dvss dvss.n2828 0.0148581
R8215 dvss dvss.n2829 0.0148581
R8216 dvss dvss.n2830 0.0148581
R8217 dvss dvss.n2831 0.0148581
R8218 dvss dvss.n2832 0.0148581
R8219 dvss.n2834 dvss 0.0148581
R8220 dvss dvss.n2839 0.0148581
R8221 dvss dvss.n2840 0.0148581
R8222 dvss dvss.n2841 0.0148581
R8223 dvss dvss.n2842 0.0148581
R8224 dvss dvss.n2843 0.0148581
R8225 dvss dvss.n2844 0.0148581
R8226 dvss dvss.n2845 0.0148581
R8227 dvss dvss.n2846 0.0148581
R8228 dvss.n2856 dvss 0.0148581
R8229 dvss dvss.n2847 0.0148581
R8230 dvss.n2854 dvss 0.0148581
R8231 dvss dvss.n2848 0.0148581
R8232 dvss dvss.n2849 0.0148581
R8233 dvss.n2858 dvss 0.0148581
R8234 dvss dvss.n2851 0.0148581
R8235 dvss dvss.n2852 0.0148581
R8236 dvss dvss.n2853 0.0148581
R8237 dvss.n2863 dvss 0.0148581
R8238 dvss dvss.n2867 0.0148581
R8239 dvss dvss.n2868 0.0148581
R8240 dvss dvss.n2869 0.0148581
R8241 dvss dvss.n2870 0.0148581
R8242 dvss dvss.n2871 0.0148581
R8243 dvss.n2873 dvss 0.0148581
R8244 dvss dvss.n2878 0.0148581
R8245 dvss.n2880 dvss 0.0148581
R8246 dvss.n2879 dvss 0.0148581
R8247 dvss dvss.n3147 0.0148581
R8248 dvss dvss.n3148 0.0148581
R8249 dvss.n3150 dvss 0.0148581
R8250 dvss.n3149 dvss 0.0148581
R8251 dvss dvss.n3158 0.0148581
R8252 dvss dvss.n3159 0.0148581
R8253 dvss dvss.n3160 0.0148581
R8254 dvss dvss.n3161 0.0148581
R8255 dvss.n3163 dvss 0.0148581
R8256 dvss.n3162 dvss 0.0148581
R8257 dvss dvss.n2098 0.0148581
R8258 dvss.n2102 dvss 0.0148581
R8259 dvss.n2101 dvss 0.0148581
R8260 dvss.n3181 dvss 0.0148581
R8261 dvss.n3180 dvss 0.0148581
R8262 dvss dvss.n3190 0.0148581
R8263 dvss dvss.n3191 0.0148581
R8264 dvss.n3193 dvss 0.0148581
R8265 dvss.n3192 dvss 0.0148581
R8266 dvss dvss.n3202 0.0148581
R8267 dvss.n3203 dvss 0.0148581
R8268 dvss.n3209 dvss 0.0148581
R8269 dvss.n3208 dvss 0.0148581
R8270 dvss dvss.n3217 0.0148581
R8271 dvss dvss.n3218 0.0148581
R8272 dvss.n3220 dvss 0.0148581
R8273 dvss.n3219 dvss 0.0148581
R8274 dvss dvss.n3229 0.0148581
R8275 dvss dvss.n3230 0.0148581
R8276 dvss.n3231 dvss 0.0148581
R8277 dvss.n3234 dvss 0.0148581
R8278 dvss.n3233 dvss 0.0148581
R8279 dvss dvss.n2011 0.0148581
R8280 dvss dvss.n2016 0.0148581
R8281 dvss dvss.n2019 0.0148581
R8282 dvss.n2022 dvss 0.0148581
R8283 dvss.n2021 dvss 0.0148581
R8284 dvss.n2020 dvss 0.0148581
R8285 dvss dvss.n2004 0.0148581
R8286 dvss.n2069 dvss 0.0148581
R8287 dvss.n2068 dvss 0.0148581
R8288 dvss.n2067 dvss 0.0148581
R8289 dvss.n2064 dvss 0.0148581
R8290 dvss.n2063 dvss 0.0148581
R8291 dvss.n2062 dvss 0.0148581
R8292 dvss.n4388 dvss 0.0148581
R8293 dvss.n4385 dvss 0.0148581
R8294 dvss.n4384 dvss 0.0148581
R8295 dvss.n4383 dvss 0.0148581
R8296 dvss.n4380 dvss 0.0148581
R8297 dvss.n4379 dvss 0.0148581
R8298 dvss.n4378 dvss 0.0148581
R8299 dvss.n4372 dvss 0.0148581
R8300 dvss.n4375 dvss 0.0148581
R8301 dvss.n4374 dvss 0.0148581
R8302 dvss dvss.n109 0.0148581
R8303 dvss.n117 dvss 0.0148581
R8304 dvss.n114 dvss 0.0148581
R8305 dvss.n113 dvss 0.0148581
R8306 dvss.n111 dvss 0.0148581
R8307 dvss.n110 dvss 0.0148581
R8308 dvss dvss.n22 0.0148581
R8309 dvss.n4364 dvss 0.0148581
R8310 dvss.n4363 dvss 0.0148581
R8311 dvss.n4362 dvss 0.0148581
R8312 dvss.n4359 dvss 0.0148581
R8313 dvss.n4358 dvss 0.0148581
R8314 dvss.n4357 dvss 0.0148581
R8315 dvss.n4354 dvss 0.0148581
R8316 dvss.n4351 dvss 0.0148581
R8317 dvss.n4350 dvss 0.0148581
R8318 dvss.n4349 dvss 0.0148581
R8319 dvss.n4346 dvss 0.0148581
R8320 dvss.n4345 dvss 0.0148581
R8321 dvss.n4344 dvss 0.0148581
R8322 dvss.n4341 dvss 0.0148581
R8323 dvss.n4340 dvss 0.0148581
R8324 dvss dvss.n44 0.0148581
R8325 dvss.n4337 dvss 0.0148581
R8326 dvss.n4336 dvss 0.0148581
R8327 dvss.n4333 dvss 0.0148581
R8328 dvss.n4329 dvss 0.0148581
R8329 dvss.n4328 dvss 0.0148581
R8330 dvss.n4325 dvss 0.0148581
R8331 dvss.n4324 dvss 0.0148581
R8332 dvss.n4323 dvss 0.0148581
R8333 dvss.n4317 dvss 0.0148581
R8334 dvss.n4316 dvss 0.0148581
R8335 dvss.n4315 dvss 0.0148581
R8336 dvss dvss.n2184 0.0148581
R8337 dvss.n2185 dvss 0.0148581
R8338 dvss dvss.n2190 0.0148581
R8339 dvss.n2192 dvss 0.0148581
R8340 dvss.n2191 dvss 0.0148581
R8341 dvss dvss.n2200 0.0148581
R8342 dvss dvss.n2201 0.0148581
R8343 dvss.n2203 dvss 0.0148581
R8344 dvss.n2202 dvss 0.0148581
R8345 dvss dvss.n2239 0.0148581
R8346 dvss dvss.n2240 0.0148581
R8347 dvss dvss.n2241 0.0148581
R8348 dvss dvss.n2242 0.0148581
R8349 dvss.n2244 dvss 0.0148581
R8350 dvss.n2243 dvss 0.0148581
R8351 dvss dvss.n2154 0.0148581
R8352 dvss.n2158 dvss 0.0148581
R8353 dvss.n2157 dvss 0.0148581
R8354 dvss.n2262 dvss 0.0148581
R8355 dvss.n2261 dvss 0.0148581
R8356 dvss dvss.n2270 0.0148581
R8357 dvss dvss.n2271 0.0148581
R8358 dvss.n2515 dvss 0.0148581
R8359 dvss.n2570 dvss 0.0148581
R8360 dvss.n2569 dvss 0.0148581
R8361 dvss.n2566 dvss 0.0148581
R8362 dvss.n2565 dvss 0.0148581
R8363 dvss dvss.n2119 0.0148581
R8364 dvss.n2562 dvss 0.0148581
R8365 dvss.n2561 dvss 0.0148581
R8366 dvss.n2558 dvss 0.0148581
R8367 dvss.n2557 dvss 0.0148581
R8368 dvss dvss.n2125 0.0148581
R8369 dvss.n2553 dvss 0.0148581
R8370 dvss.n2552 dvss 0.0148581
R8371 dvss.n2549 dvss 0.0148581
R8372 dvss.n2545 dvss 0.0148581
R8373 dvss.n2544 dvss 0.0148581
R8374 dvss.n2541 dvss 0.0148581
R8375 dvss.n2540 dvss 0.0148581
R8376 dvss.n2539 dvss 0.0148581
R8377 dvss.n2535 dvss 0.0148581
R8378 dvss.n2534 dvss 0.0148581
R8379 dvss.n2531 dvss 0.0148581
R8380 dvss.n2530 dvss 0.0148581
R8381 dvss.n2529 dvss 0.0148581
R8382 dvss.n2526 dvss 0.0148581
R8383 dvss.n2525 dvss 0.0148581
R8384 dvss.n2524 dvss 0.0148581
R8385 dvss.n1098 dvss 0.0145449
R8386 dvss dvss.n2663 0.0140135
R8387 dvss dvss.n2129 0.0140135
R8388 dvss dvss.n893 0.0134032
R8389 dvss dvss.n900 0.0134032
R8390 dvss.n1295 dvss 0.0134032
R8391 dvss dvss.n1311 0.0134032
R8392 dvss.n1354 dvss 0.0134032
R8393 dvss dvss.n1430 0.0134032
R8394 dvss.n1778 dvss 0.0134032
R8395 dvss dvss.n1794 0.0134032
R8396 dvss.n1837 dvss 0.0134032
R8397 dvss dvss.n3379 0.0134032
R8398 dvss.n1869 dvss 0.0134032
R8399 dvss dvss.n3324 0.0134032
R8400 dvss.n1900 dvss 0.0134032
R8401 dvss dvss.n3274 0.0134032
R8402 dvss.n3909 dvss 0.0134032
R8403 dvss dvss.n3925 0.0134032
R8404 dvss.n3963 dvss 0.0134032
R8405 dvss dvss.n4036 0.0134032
R8406 dvss.n1174 dvss 0.0127893
R8407 dvss.n715 dvss 0.0127893
R8408 dvss.n1561 dvss 0.0127893
R8409 dvss.n1709 dvss 0.0127893
R8410 dvss.n3512 dvss 0.0127893
R8411 dvss.n3625 dvss 0.0127893
R8412 dvss.n3744 dvss 0.0127893
R8413 dvss.n4145 dvss 0.0127893
R8414 dvss.n4193 dvss 0.0127893
R8415 dvss.n907 dvss 0.0125968
R8416 dvss.n918 dvss 0.0125968
R8417 dvss dvss.n1285 0.0125968
R8418 dvss.n1312 dvss 0.0125968
R8419 dvss dvss.n1443 0.0125968
R8420 dvss.n1431 dvss 0.0125968
R8421 dvss dvss.n1768 0.0125968
R8422 dvss.n1795 dvss 0.0125968
R8423 dvss dvss.n3392 0.0125968
R8424 dvss.n3380 dvss 0.0125968
R8425 dvss dvss.n3337 0.0125968
R8426 dvss.n3325 dvss 0.0125968
R8427 dvss dvss.n3287 0.0125968
R8428 dvss.n3275 dvss 0.0125968
R8429 dvss dvss.n3899 0.0125968
R8430 dvss.n3926 dvss 0.0125968
R8431 dvss dvss.n4049 0.0125968
R8432 dvss.n4037 dvss 0.0125968
R8433 dvss.n2678 dvss 0.0123243
R8434 dvss.n2717 dvss 0.0123243
R8435 dvss.n2756 dvss 0.0123243
R8436 dvss.n2795 dvss 0.0123243
R8437 dvss.n2834 dvss 0.0123243
R8438 dvss.n2873 dvss 0.0123243
R8439 dvss.n3203 dvss 0.0123243
R8440 dvss dvss.n2062 0.0123243
R8441 dvss dvss.n4357 0.0123243
R8442 dvss.n2185 dvss 0.0123243
R8443 dvss.n1123 dvss 0.011736
R8444 dvss dvss.n1151 0.011736
R8445 dvss dvss.n644 0.011736
R8446 dvss dvss.n653 0.011736
R8447 dvss dvss.n1509 0.011736
R8448 dvss.n1534 dvss 0.011736
R8449 dvss.n1729 dvss 0.011736
R8450 dvss.n1720 dvss 0.011736
R8451 dvss dvss.n3460 0.011736
R8452 dvss.n3485 dvss 0.011736
R8453 dvss dvss.n375 0.011736
R8454 dvss dvss.n3592 0.011736
R8455 dvss.n3689 dvss 0.011736
R8456 dvss.n3714 dvss 0.011736
R8457 dvss.n3860 dvss 0.011736
R8458 dvss.n3851 dvss 0.011736
R8459 dvss.n4116 dvss 0.011736
R8460 dvss.n4107 dvss 0.011736
R8461 dvss dvss.n2694 0.0114797
R8462 dvss dvss.n2710 0.0114797
R8463 dvss dvss.n2733 0.0114797
R8464 dvss dvss.n2749 0.0114797
R8465 dvss dvss.n2772 0.0114797
R8466 dvss dvss.n2788 0.0114797
R8467 dvss dvss.n2811 0.0114797
R8468 dvss dvss.n2827 0.0114797
R8469 dvss dvss.n2850 0.0114797
R8470 dvss dvss.n2866 0.0114797
R8471 dvss.n3173 dvss 0.0114797
R8472 dvss.n3177 dvss 0.0114797
R8473 dvss dvss.n2018 0.0114797
R8474 dvss.n2072 dvss 0.0114797
R8475 dvss.n115 dvss 0.0114797
R8476 dvss.n4367 dvss 0.0114797
R8477 dvss dvss.n48 0.0114797
R8478 dvss.n4320 dvss 0.0114797
R8479 dvss.n2254 dvss 0.0114797
R8480 dvss.n2258 dvss 0.0114797
R8481 dvss dvss.n2539 0.0114797
R8482 dvss.n1122 dvss 0.0110337
R8483 dvss.n1152 dvss 0.0110337
R8484 dvss.n720 dvss 0.0110337
R8485 dvss.n1233 dvss 0.0110337
R8486 dvss.n1510 dvss 0.0110337
R8487 dvss dvss.n1529 0.0110337
R8488 dvss.n1604 dvss 0.0110337
R8489 dvss.n1714 dvss 0.0110337
R8490 dvss.n3461 dvss 0.0110337
R8491 dvss dvss.n3480 0.0110337
R8492 dvss dvss.n376 0.0110337
R8493 dvss.n3593 dvss 0.0110337
R8494 dvss dvss.n3693 0.0110337
R8495 dvss.n3712 dvss 0.0110337
R8496 dvss.n3787 dvss 0.0110337
R8497 dvss.n3845 dvss 0.0110337
R8498 dvss.n161 dvss 0.0110337
R8499 dvss.n4101 dvss 0.0110337
R8500 dvss dvss.n748 0.00998034
R8501 dvss.n670 dvss 0.00998034
R8502 dvss dvss.n1550 0.00998034
R8503 dvss.n1625 dvss 0.00998034
R8504 dvss dvss.n3501 0.00998034
R8505 dvss dvss.n3617 0.00998034
R8506 dvss dvss.n3733 0.00998034
R8507 dvss.n135 dvss 0.00998034
R8508 dvss.n4192 dvss 0.00998034
R8509 dvss dvss.n2691 0.00979054
R8510 dvss dvss.n2695 0.00979054
R8511 dvss dvss.n2730 0.00979054
R8512 dvss dvss.n2734 0.00979054
R8513 dvss dvss.n2769 0.00979054
R8514 dvss dvss.n2773 0.00979054
R8515 dvss dvss.n2808 0.00979054
R8516 dvss dvss.n2812 0.00979054
R8517 dvss dvss.n2847 0.00979054
R8518 dvss dvss.n2851 0.00979054
R8519 dvss.n3160 dvss 0.00979054
R8520 dvss.n2102 dvss 0.00979054
R8521 dvss.n3234 dvss 0.00979054
R8522 dvss.n2022 dvss 0.00979054
R8523 dvss.n4375 dvss 0.00979054
R8524 dvss dvss.n113 0.00979054
R8525 dvss.n44 dvss 0.00979054
R8526 dvss dvss.n4328 0.00979054
R8527 dvss.n2241 dvss 0.00979054
R8528 dvss.n2158 dvss 0.00979054
R8529 dvss.n2536 dvss 0.00979054
R8530 dvss.n883 dvss 0.00896774
R8531 dvss dvss.n2682 0.00894595
R8532 dvss dvss.n2721 0.00894595
R8533 dvss dvss.n2760 0.00894595
R8534 dvss dvss.n2799 0.00894595
R8535 dvss dvss.n2838 0.00894595
R8536 dvss dvss.n2877 0.00894595
R8537 dvss dvss.n3207 0.00894595
R8538 dvss.n2060 dvss 0.00894595
R8539 dvss.n4355 dvss 0.00894595
R8540 dvss dvss.n2189 0.00894595
R8541 dvss.n4389 dvss 0.00810135
R8542 dvss.n1065 dvss 0.00752247
R8543 dvss dvss.n841 0.00735484
R8544 dvss dvss.n842 0.00735484
R8545 dvss dvss.n847 0.00735484
R8546 dvss dvss.n848 0.00735484
R8547 dvss dvss.n849 0.00735484
R8548 dvss dvss.n850 0.00735484
R8549 dvss dvss.n858 0.00735484
R8550 dvss dvss.n859 0.00735484
R8551 dvss dvss.n860 0.00735484
R8552 dvss dvss.n872 0.00735484
R8553 dvss dvss.n873 0.00735484
R8554 dvss.n881 dvss 0.00735484
R8555 dvss dvss.n874 0.00735484
R8556 dvss dvss.n874 0.00735484
R8557 dvss dvss.n883 0.00735484
R8558 dvss dvss.n884 0.00735484
R8559 dvss dvss.n885 0.00735484
R8560 dvss dvss.n886 0.00735484
R8561 dvss dvss.n887 0.00735484
R8562 dvss dvss.n891 0.00735484
R8563 dvss dvss.n892 0.00735484
R8564 dvss.n907 dvss 0.00735484
R8565 dvss dvss.n893 0.00735484
R8566 dvss.n910 dvss 0.00735484
R8567 dvss dvss.n894 0.00735484
R8568 dvss dvss.n913 0.00735484
R8569 dvss.n914 dvss 0.00735484
R8570 dvss dvss.n899 0.00735484
R8571 dvss.n918 dvss 0.00735484
R8572 dvss dvss.n900 0.00735484
R8573 dvss dvss.n901 0.00735484
R8574 dvss dvss.n924 0.00735484
R8575 dvss dvss.n925 0.00735484
R8576 dvss dvss.n926 0.00735484
R8577 dvss dvss.n927 0.00735484
R8578 dvss.n931 dvss 0.00735484
R8579 dvss dvss.n937 0.00735484
R8580 dvss dvss.n938 0.00735484
R8581 dvss.n940 dvss 0.00735484
R8582 dvss.n939 dvss 0.00735484
R8583 dvss dvss.n1272 0.00735484
R8584 dvss dvss.n1273 0.00735484
R8585 dvss.n1275 dvss 0.00735484
R8586 dvss.n1274 dvss 0.00735484
R8587 dvss dvss.n1283 0.00735484
R8588 dvss dvss.n1284 0.00735484
R8589 dvss.n1287 dvss 0.00735484
R8590 dvss.n1286 dvss 0.00735484
R8591 dvss.n1285 dvss 0.00735484
R8592 dvss dvss.n1295 0.00735484
R8593 dvss.n1297 dvss 0.00735484
R8594 dvss.n1296 dvss 0.00735484
R8595 dvss.n1302 dvss 0.00735484
R8596 dvss.n1301 dvss 0.00735484
R8597 dvss.n610 dvss 0.00735484
R8598 dvss.n1312 dvss 0.00735484
R8599 dvss.n1311 dvss 0.00735484
R8600 dvss.n604 dvss 0.00735484
R8601 dvss.n1316 dvss 0.00735484
R8602 dvss.n601 dvss 0.00735484
R8603 dvss dvss.n1326 0.00735484
R8604 dvss dvss.n1327 0.00735484
R8605 dvss.n1328 dvss 0.00735484
R8606 dvss.n594 dvss 0.00735484
R8607 dvss.n593 dvss 0.00735484
R8608 dvss dvss.n1340 0.00735484
R8609 dvss dvss.n1346 0.00735484
R8610 dvss.n1455 dvss 0.00735484
R8611 dvss.n1454 dvss 0.00735484
R8612 dvss.n1453 dvss 0.00735484
R8613 dvss.n1450 dvss 0.00735484
R8614 dvss.n1449 dvss 0.00735484
R8615 dvss.n1448 dvss 0.00735484
R8616 dvss.n1445 dvss 0.00735484
R8617 dvss.n1444 dvss 0.00735484
R8618 dvss.n1443 dvss 0.00735484
R8619 dvss.n1354 dvss 0.00735484
R8620 dvss.n1440 dvss 0.00735484
R8621 dvss.n1439 dvss 0.00735484
R8622 dvss.n1436 dvss 0.00735484
R8623 dvss.n1435 dvss 0.00735484
R8624 dvss dvss.n1361 0.00735484
R8625 dvss.n1431 dvss 0.00735484
R8626 dvss.n1430 dvss 0.00735484
R8627 dvss.n1427 dvss 0.00735484
R8628 dvss.n1423 dvss 0.00735484
R8629 dvss.n1422 dvss 0.00735484
R8630 dvss.n1419 dvss 0.00735484
R8631 dvss.n1418 dvss 0.00735484
R8632 dvss.n1417 dvss 0.00735484
R8633 dvss.n1413 dvss 0.00735484
R8634 dvss.n1412 dvss 0.00735484
R8635 dvss.n1409 dvss 0.00735484
R8636 dvss.n1403 dvss 0.00735484
R8637 dvss dvss.n1755 0.00735484
R8638 dvss dvss.n1756 0.00735484
R8639 dvss.n1758 dvss 0.00735484
R8640 dvss.n1757 dvss 0.00735484
R8641 dvss dvss.n1766 0.00735484
R8642 dvss dvss.n1767 0.00735484
R8643 dvss.n1770 dvss 0.00735484
R8644 dvss.n1769 dvss 0.00735484
R8645 dvss.n1768 dvss 0.00735484
R8646 dvss dvss.n1778 0.00735484
R8647 dvss.n1780 dvss 0.00735484
R8648 dvss.n1779 dvss 0.00735484
R8649 dvss.n1785 dvss 0.00735484
R8650 dvss.n1784 dvss 0.00735484
R8651 dvss.n490 dvss 0.00735484
R8652 dvss.n1795 dvss 0.00735484
R8653 dvss.n1794 dvss 0.00735484
R8654 dvss.n484 dvss 0.00735484
R8655 dvss.n1799 dvss 0.00735484
R8656 dvss.n481 dvss 0.00735484
R8657 dvss dvss.n1809 0.00735484
R8658 dvss dvss.n1810 0.00735484
R8659 dvss.n1811 dvss 0.00735484
R8660 dvss.n474 dvss 0.00735484
R8661 dvss.n473 dvss 0.00735484
R8662 dvss dvss.n1823 0.00735484
R8663 dvss dvss.n1829 0.00735484
R8664 dvss.n3404 dvss 0.00735484
R8665 dvss.n3403 dvss 0.00735484
R8666 dvss.n3402 dvss 0.00735484
R8667 dvss.n3399 dvss 0.00735484
R8668 dvss.n3398 dvss 0.00735484
R8669 dvss.n3397 dvss 0.00735484
R8670 dvss.n3394 dvss 0.00735484
R8671 dvss.n3393 dvss 0.00735484
R8672 dvss.n3392 dvss 0.00735484
R8673 dvss.n1837 dvss 0.00735484
R8674 dvss.n3389 dvss 0.00735484
R8675 dvss.n3388 dvss 0.00735484
R8676 dvss.n3385 dvss 0.00735484
R8677 dvss.n3384 dvss 0.00735484
R8678 dvss dvss.n1844 0.00735484
R8679 dvss.n3380 dvss 0.00735484
R8680 dvss.n3379 dvss 0.00735484
R8681 dvss.n3376 dvss 0.00735484
R8682 dvss.n3372 dvss 0.00735484
R8683 dvss.n3371 dvss 0.00735484
R8684 dvss.n3368 dvss 0.00735484
R8685 dvss.n3367 dvss 0.00735484
R8686 dvss.n3366 dvss 0.00735484
R8687 dvss.n3362 dvss 0.00735484
R8688 dvss.n3361 dvss 0.00735484
R8689 dvss.n3358 dvss 0.00735484
R8690 dvss.n3352 dvss 0.00735484
R8691 dvss.n3351 dvss 0.00735484
R8692 dvss.n3348 dvss 0.00735484
R8693 dvss.n3347 dvss 0.00735484
R8694 dvss.n3346 dvss 0.00735484
R8695 dvss.n3343 dvss 0.00735484
R8696 dvss.n3342 dvss 0.00735484
R8697 dvss.n3341 dvss 0.00735484
R8698 dvss.n3338 dvss 0.00735484
R8699 dvss.n3337 dvss 0.00735484
R8700 dvss dvss.n1869 0.00735484
R8701 dvss.n3334 dvss 0.00735484
R8702 dvss.n3333 dvss 0.00735484
R8703 dvss.n3330 dvss 0.00735484
R8704 dvss.n3329 dvss 0.00735484
R8705 dvss dvss.n1875 0.00735484
R8706 dvss.n3325 dvss 0.00735484
R8707 dvss.n3324 dvss 0.00735484
R8708 dvss.n3321 dvss 0.00735484
R8709 dvss.n3317 dvss 0.00735484
R8710 dvss.n3316 dvss 0.00735484
R8711 dvss.n3313 dvss 0.00735484
R8712 dvss.n3312 dvss 0.00735484
R8713 dvss.n3311 dvss 0.00735484
R8714 dvss.n3307 dvss 0.00735484
R8715 dvss.n3306 dvss 0.00735484
R8716 dvss.n3303 dvss 0.00735484
R8717 dvss.n3302 dvss 0.00735484
R8718 dvss.n3301 dvss 0.00735484
R8719 dvss.n3298 dvss 0.00735484
R8720 dvss.n3297 dvss 0.00735484
R8721 dvss.n3296 dvss 0.00735484
R8722 dvss.n3293 dvss 0.00735484
R8723 dvss.n3292 dvss 0.00735484
R8724 dvss.n3291 dvss 0.00735484
R8725 dvss.n3288 dvss 0.00735484
R8726 dvss.n3287 dvss 0.00735484
R8727 dvss dvss.n1900 0.00735484
R8728 dvss.n3284 dvss 0.00735484
R8729 dvss.n3283 dvss 0.00735484
R8730 dvss.n3280 dvss 0.00735484
R8731 dvss.n3279 dvss 0.00735484
R8732 dvss dvss.n1906 0.00735484
R8733 dvss.n3275 dvss 0.00735484
R8734 dvss.n3274 dvss 0.00735484
R8735 dvss.n3271 dvss 0.00735484
R8736 dvss.n3267 dvss 0.00735484
R8737 dvss.n3266 dvss 0.00735484
R8738 dvss.n3263 dvss 0.00735484
R8739 dvss.n3262 dvss 0.00735484
R8740 dvss.n3261 dvss 0.00735484
R8741 dvss.n3257 dvss 0.00735484
R8742 dvss.n3256 dvss 0.00735484
R8743 dvss.n3253 dvss 0.00735484
R8744 dvss.n3252 dvss 0.00735484
R8745 dvss dvss.n3886 0.00735484
R8746 dvss dvss.n3887 0.00735484
R8747 dvss.n3889 dvss 0.00735484
R8748 dvss.n3888 dvss 0.00735484
R8749 dvss dvss.n3897 0.00735484
R8750 dvss dvss.n3898 0.00735484
R8751 dvss.n3901 dvss 0.00735484
R8752 dvss.n3900 dvss 0.00735484
R8753 dvss.n3899 dvss 0.00735484
R8754 dvss dvss.n3909 0.00735484
R8755 dvss.n3911 dvss 0.00735484
R8756 dvss.n3910 dvss 0.00735484
R8757 dvss.n3916 dvss 0.00735484
R8758 dvss.n3915 dvss 0.00735484
R8759 dvss.n244 dvss 0.00735484
R8760 dvss.n3926 dvss 0.00735484
R8761 dvss.n3925 dvss 0.00735484
R8762 dvss.n238 dvss 0.00735484
R8763 dvss.n3930 dvss 0.00735484
R8764 dvss.n235 dvss 0.00735484
R8765 dvss dvss.n3940 0.00735484
R8766 dvss dvss.n3941 0.00735484
R8767 dvss.n3942 dvss 0.00735484
R8768 dvss.n228 dvss 0.00735484
R8769 dvss.n227 dvss 0.00735484
R8770 dvss dvss.n3954 0.00735484
R8771 dvss dvss.n3955 0.00735484
R8772 dvss.n4061 dvss 0.00735484
R8773 dvss.n4060 dvss 0.00735484
R8774 dvss.n4059 dvss 0.00735484
R8775 dvss.n4056 dvss 0.00735484
R8776 dvss.n4055 dvss 0.00735484
R8777 dvss.n4054 dvss 0.00735484
R8778 dvss.n4051 dvss 0.00735484
R8779 dvss.n4050 dvss 0.00735484
R8780 dvss.n4049 dvss 0.00735484
R8781 dvss.n3963 dvss 0.00735484
R8782 dvss.n4046 dvss 0.00735484
R8783 dvss.n4045 dvss 0.00735484
R8784 dvss.n4042 dvss 0.00735484
R8785 dvss.n4041 dvss 0.00735484
R8786 dvss dvss.n3970 0.00735484
R8787 dvss.n4037 dvss 0.00735484
R8788 dvss.n4036 dvss 0.00735484
R8789 dvss.n4033 dvss 0.00735484
R8790 dvss.n4029 dvss 0.00735484
R8791 dvss.n4028 dvss 0.00735484
R8792 dvss.n4025 dvss 0.00735484
R8793 dvss.n4024 dvss 0.00735484
R8794 dvss.n4023 dvss 0.00735484
R8795 dvss.n4019 dvss 0.00735484
R8796 dvss.n4018 dvss 0.00735484
R8797 dvss.n4015 dvss 0.00735484
R8798 dvss.n4014 dvss 0.00735484
R8799 dvss.n4013 dvss 0.00735484
R8800 dvss.n4306 dvss 0.00735484
R8801 dvss.n4305 dvss 0.00735484
R8802 dvss.n4304 dvss 0.00735484
R8803 dvss.n4389 dvss.n9 0.00725676
R8804 dvss.n2125 dvss 0.00725676
R8805 dvss dvss.n2544 0.00725676
R8806 dvss.n859 dvss 0.00695161
R8807 dvss.n921 dvss 0.00695161
R8808 dvss.n1317 dvss 0.00695161
R8809 dvss dvss.n1365 0.00695161
R8810 dvss.n1800 dvss 0.00695161
R8811 dvss dvss.n1848 0.00695161
R8812 dvss dvss.n1879 0.00695161
R8813 dvss dvss.n1910 0.00695161
R8814 dvss.n3931 dvss 0.00695161
R8815 dvss dvss.n3990 0.00695161
R8816 dvss.n868 dvss.n861 0.00654839
R8817 dvss dvss.n1031 0.0064691
R8818 dvss dvss.n1107 0.0064691
R8819 dvss.n1113 dvss 0.0064691
R8820 dvss.n1112 dvss 0.0064691
R8821 dvss dvss.n1121 0.0064691
R8822 dvss dvss.n1122 0.0064691
R8823 dvss.n1123 dvss 0.0064691
R8824 dvss.n1131 dvss 0.0064691
R8825 dvss.n1130 dvss 0.0064691
R8826 dvss.n1136 dvss 0.0064691
R8827 dvss.n1135 dvss 0.0064691
R8828 dvss.n766 dvss 0.0064691
R8829 dvss.n1152 dvss 0.0064691
R8830 dvss.n1151 dvss 0.0064691
R8831 dvss.n1142 dvss 0.0064691
R8832 dvss.n749 dvss 0.0064691
R8833 dvss.n748 dvss 0.0064691
R8834 dvss.n1174 dvss 0.0064691
R8835 dvss.n1173 dvss 0.0064691
R8836 dvss.n1172 dvss 0.0064691
R8837 dvss.n1188 dvss 0.0064691
R8838 dvss.n1187 dvss 0.0064691
R8839 dvss.n1198 dvss 0.0064691
R8840 dvss.n1197 dvss 0.0064691
R8841 dvss dvss.n632 0.0064691
R8842 dvss dvss.n633 0.0064691
R8843 dvss dvss.n1207 0.0064691
R8844 dvss dvss.n1210 0.0064691
R8845 dvss.n1216 dvss 0.0064691
R8846 dvss.n1215 dvss 0.0064691
R8847 dvss dvss.n643 0.0064691
R8848 dvss.n720 dvss 0.0064691
R8849 dvss dvss.n644 0.0064691
R8850 dvss.n1226 dvss 0.0064691
R8851 dvss.n1225 dvss 0.0064691
R8852 dvss dvss.n651 0.0064691
R8853 dvss.n1229 dvss 0.0064691
R8854 dvss dvss.n652 0.0064691
R8855 dvss.n1233 dvss 0.0064691
R8856 dvss dvss.n653 0.0064691
R8857 dvss.n1238 dvss 0.0064691
R8858 dvss.n718 dvss 0.0064691
R8859 dvss dvss.n670 0.0064691
R8860 dvss.n715 dvss 0.0064691
R8861 dvss.n714 dvss 0.0064691
R8862 dvss.n713 dvss 0.0064691
R8863 dvss.n704 dvss 0.0064691
R8864 dvss.n701 dvss 0.0064691
R8865 dvss dvss.n1464 0.0064691
R8866 dvss.n1465 dvss 0.0064691
R8867 dvss dvss.n569 0.0064691
R8868 dvss.n1486 dvss 0.0064691
R8869 dvss.n1483 dvss 0.0064691
R8870 dvss.n1482 dvss 0.0064691
R8871 dvss dvss.n1496 0.0064691
R8872 dvss.n1497 dvss 0.0064691
R8873 dvss.n1502 dvss 0.0064691
R8874 dvss.n1510 dvss 0.0064691
R8875 dvss.n1509 dvss 0.0064691
R8876 dvss dvss.n1514 0.0064691
R8877 dvss.n1515 dvss 0.0064691
R8878 dvss dvss.n1522 0.0064691
R8879 dvss.n1523 dvss 0.0064691
R8880 dvss.n1530 dvss 0.0064691
R8881 dvss.n1529 dvss 0.0064691
R8882 dvss.n1534 dvss 0.0064691
R8883 dvss.n1533 dvss 0.0064691
R8884 dvss.n1551 dvss 0.0064691
R8885 dvss.n1550 dvss 0.0064691
R8886 dvss.n1561 dvss 0.0064691
R8887 dvss.n1560 dvss 0.0064691
R8888 dvss.n1559 dvss 0.0064691
R8889 dvss.n1575 dvss 0.0064691
R8890 dvss.n1574 dvss 0.0064691
R8891 dvss.n1584 dvss 0.0064691
R8892 dvss.n1583 dvss 0.0064691
R8893 dvss.n1742 dvss 0.0064691
R8894 dvss.n1741 dvss 0.0064691
R8895 dvss.n1740 dvss 0.0064691
R8896 dvss.n1737 dvss 0.0064691
R8897 dvss.n1736 dvss 0.0064691
R8898 dvss.n1735 dvss 0.0064691
R8899 dvss.n1732 dvss 0.0064691
R8900 dvss.n1604 dvss 0.0064691
R8901 dvss.n1729 dvss 0.0064691
R8902 dvss.n1728 dvss 0.0064691
R8903 dvss dvss.n1667 0.0064691
R8904 dvss.n1668 dvss 0.0064691
R8905 dvss.n1724 dvss 0.0064691
R8906 dvss.n1723 dvss 0.0064691
R8907 dvss.n1714 dvss 0.0064691
R8908 dvss.n1720 dvss 0.0064691
R8909 dvss.n1719 dvss 0.0064691
R8910 dvss.n1712 dvss 0.0064691
R8911 dvss dvss.n1625 0.0064691
R8912 dvss.n1709 dvss 0.0064691
R8913 dvss.n1708 dvss 0.0064691
R8914 dvss.n1707 dvss 0.0064691
R8915 dvss.n1698 dvss 0.0064691
R8916 dvss.n1695 dvss 0.0064691
R8917 dvss dvss.n3413 0.0064691
R8918 dvss.n3414 dvss 0.0064691
R8919 dvss.n3438 dvss 0.0064691
R8920 dvss.n3435 dvss 0.0064691
R8921 dvss.n3434 dvss 0.0064691
R8922 dvss.n3433 dvss 0.0064691
R8923 dvss dvss.n3447 0.0064691
R8924 dvss.n3448 dvss 0.0064691
R8925 dvss.n3453 dvss 0.0064691
R8926 dvss.n3461 dvss 0.0064691
R8927 dvss.n3460 dvss 0.0064691
R8928 dvss dvss.n3465 0.0064691
R8929 dvss.n3466 dvss 0.0064691
R8930 dvss dvss.n3473 0.0064691
R8931 dvss.n3474 dvss 0.0064691
R8932 dvss.n3481 dvss 0.0064691
R8933 dvss.n3480 dvss 0.0064691
R8934 dvss.n3485 dvss 0.0064691
R8935 dvss.n3484 dvss 0.0064691
R8936 dvss.n3502 dvss 0.0064691
R8937 dvss.n3501 dvss 0.0064691
R8938 dvss.n3512 dvss 0.0064691
R8939 dvss.n3511 dvss 0.0064691
R8940 dvss.n3510 dvss 0.0064691
R8941 dvss.n3527 dvss 0.0064691
R8942 dvss.n3526 dvss 0.0064691
R8943 dvss.n3536 dvss 0.0064691
R8944 dvss.n3535 dvss 0.0064691
R8945 dvss.n393 dvss 0.0064691
R8946 dvss.n3558 dvss 0.0064691
R8947 dvss.n3555 dvss 0.0064691
R8948 dvss.n3554 dvss 0.0064691
R8949 dvss dvss.n3566 0.0064691
R8950 dvss.n3567 dvss 0.0064691
R8951 dvss.n3575 dvss 0.0064691
R8952 dvss.n376 dvss 0.0064691
R8953 dvss.n375 dvss 0.0064691
R8954 dvss.n3587 dvss 0.0064691
R8955 dvss.n3586 dvss 0.0064691
R8956 dvss.n3598 dvss 0.0064691
R8957 dvss.n3597 dvss 0.0064691
R8958 dvss.n3601 dvss 0.0064691
R8959 dvss.n3593 dvss 0.0064691
R8960 dvss.n3592 dvss 0.0064691
R8961 dvss.n3610 dvss 0.0064691
R8962 dvss.n3618 dvss 0.0064691
R8963 dvss.n3617 dvss 0.0064691
R8964 dvss dvss.n3625 0.0064691
R8965 dvss.n3632 dvss 0.0064691
R8966 dvss.n3631 dvss 0.0064691
R8967 dvss.n3644 dvss 0.0064691
R8968 dvss.n3643 dvss 0.0064691
R8969 dvss.n3653 dvss 0.0064691
R8970 dvss.n3652 dvss 0.0064691
R8971 dvss.n3656 dvss 0.0064691
R8972 dvss.n3671 dvss 0.0064691
R8973 dvss.n3670 dvss 0.0064691
R8974 dvss.n3669 dvss 0.0064691
R8975 dvss dvss.n3679 0.0064691
R8976 dvss.n3680 dvss 0.0064691
R8977 dvss.n3694 dvss 0.0064691
R8978 dvss.n3693 dvss 0.0064691
R8979 dvss dvss.n3689 0.0064691
R8980 dvss.n3690 dvss 0.0064691
R8981 dvss dvss.n3704 0.0064691
R8982 dvss dvss.n3705 0.0064691
R8983 dvss.n3706 dvss 0.0064691
R8984 dvss.n3717 dvss 0.0064691
R8985 dvss dvss.n3712 0.0064691
R8986 dvss.n3714 dvss 0.0064691
R8987 dvss.n3713 dvss 0.0064691
R8988 dvss.n3734 dvss 0.0064691
R8989 dvss.n3733 dvss 0.0064691
R8990 dvss.n3744 dvss 0.0064691
R8991 dvss.n3743 dvss 0.0064691
R8992 dvss.n3742 dvss 0.0064691
R8993 dvss.n3758 dvss 0.0064691
R8994 dvss.n3757 dvss 0.0064691
R8995 dvss.n3767 dvss 0.0064691
R8996 dvss.n3766 dvss 0.0064691
R8997 dvss.n3873 dvss 0.0064691
R8998 dvss.n3872 dvss 0.0064691
R8999 dvss.n3871 dvss 0.0064691
R9000 dvss.n3868 dvss 0.0064691
R9001 dvss.n3867 dvss 0.0064691
R9002 dvss.n3866 dvss 0.0064691
R9003 dvss.n3863 dvss 0.0064691
R9004 dvss.n3787 dvss 0.0064691
R9005 dvss.n3860 dvss 0.0064691
R9006 dvss.n3859 dvss 0.0064691
R9007 dvss dvss.n3805 0.0064691
R9008 dvss.n3806 dvss 0.0064691
R9009 dvss.n3855 dvss 0.0064691
R9010 dvss.n3854 dvss 0.0064691
R9011 dvss.n3845 dvss 0.0064691
R9012 dvss.n3851 dvss 0.0064691
R9013 dvss.n3850 dvss 0.0064691
R9014 dvss.n4148 dvss 0.0064691
R9015 dvss.n135 dvss 0.0064691
R9016 dvss.n4145 dvss 0.0064691
R9017 dvss.n4144 dvss 0.0064691
R9018 dvss.n4143 dvss 0.0064691
R9019 dvss.n204 dvss 0.0064691
R9020 dvss dvss.n211 0.0064691
R9021 dvss.n212 dvss 0.0064691
R9022 dvss dvss.n138 0.0064691
R9023 dvss.n4129 dvss 0.0064691
R9024 dvss.n4128 dvss 0.0064691
R9025 dvss.n4127 dvss 0.0064691
R9026 dvss.n4124 dvss 0.0064691
R9027 dvss.n4123 dvss 0.0064691
R9028 dvss.n4122 dvss 0.0064691
R9029 dvss.n4119 dvss 0.0064691
R9030 dvss.n161 dvss 0.0064691
R9031 dvss.n4116 dvss 0.0064691
R9032 dvss.n4115 dvss 0.0064691
R9033 dvss dvss.n4083 0.0064691
R9034 dvss.n4084 dvss 0.0064691
R9035 dvss.n4111 dvss 0.0064691
R9036 dvss.n4110 dvss 0.0064691
R9037 dvss.n4101 dvss 0.0064691
R9038 dvss.n4107 dvss 0.0064691
R9039 dvss.n4106 dvss 0.0064691
R9040 dvss dvss.n4191 0.0064691
R9041 dvss dvss.n4192 0.0064691
R9042 dvss.n4193 dvss 0.0064691
R9043 dvss dvss.n4202 0.0064691
R9044 dvss.n4203 dvss 0.0064691
R9045 dvss.n4209 dvss 0.0064691
R9046 dvss.n4219 dvss 0.0064691
R9047 dvss.n4218 dvss 0.0064691
R9048 dvss.n4217 dvss 0.0064691
R9049 dvss dvss.n4233 0.0064691
R9050 dvss.n4234 dvss 0.0064691
R9051 dvss dvss.n4241 0.0064691
R9052 dvss.n2682 dvss.n2677 0.00641216
R9053 dvss.n2721 dvss.n2716 0.00641216
R9054 dvss.n2760 dvss.n2755 0.00641216
R9055 dvss.n2799 dvss.n2794 0.00641216
R9056 dvss.n2838 dvss.n2833 0.00641216
R9057 dvss.n2877 dvss.n2872 0.00641216
R9058 dvss.n3207 dvss.n2086 0.00641216
R9059 dvss.n2060 dvss.n2059 0.00641216
R9060 dvss.n4355 dvss.n32 0.00641216
R9061 dvss.n2189 dvss.n2174 0.00641216
R9062 dvss dvss.n1020 0.00611798
R9063 dvss dvss.n1022 0.00611798
R9064 dvss dvss.n805 0.00611798
R9065 dvss dvss.n806 0.00611798
R9066 dvss dvss.n807 0.00611798
R9067 dvss dvss.n808 0.00611798
R9068 dvss dvss.n809 0.00611798
R9069 dvss.n1032 dvss 0.00611798
R9070 dvss dvss.n811 0.00611798
R9071 dvss dvss.n812 0.00611798
R9072 dvss.n1070 dvss 0.00611798
R9073 dvss.n1068 dvss 0.00611798
R9074 dvss.n1057 dvss 0.00611798
R9075 dvss dvss.n785 0.00611798
R9076 dvss dvss.n1059 0.00611798
R9077 dvss.n1064 dvss 0.00611798
R9078 dvss.n1097 dvss 0.00611798
R9079 dvss.n788 dvss 0.00611798
R9080 dvss.n1158 dvss 0.00611798
R9081 dvss dvss.n662 0.00611798
R9082 dvss.n1546 dvss 0.00611798
R9083 dvss dvss.n1616 0.00611798
R9084 dvss.n3497 dvss 0.00611798
R9085 dvss.n3613 dvss 0.00611798
R9086 dvss.n3729 dvss 0.00611798
R9087 dvss dvss.n3842 0.00611798
R9088 dvss dvss.n4098 0.00611798
R9089 dvss.n931 dvss 0.00574194
R9090 dvss.n1328 dvss 0.00574194
R9091 dvss dvss.n1417 0.00574194
R9092 dvss.n1811 dvss 0.00574194
R9093 dvss dvss.n3366 0.00574194
R9094 dvss dvss.n3311 0.00574194
R9095 dvss dvss.n3261 0.00574194
R9096 dvss.n3942 dvss 0.00574194
R9097 dvss dvss.n4023 0.00574194
R9098 dvss.n2657 dvss 0.00556757
R9099 dvss.n2562 dvss 0.00556757
R9100 dvss.n2536 dvss.n2135 0.00556757
R9101 dvss.n819 dvss.n813 0.00541573
R9102 dvss dvss.n1112 0.00541573
R9103 dvss.n1156 dvss 0.00541573
R9104 dvss dvss.n1215 0.00541573
R9105 dvss.n719 dvss 0.00541573
R9106 dvss.n1497 dvss 0.00541573
R9107 dvss dvss.n1549 0.00541573
R9108 dvss dvss.n1735 0.00541573
R9109 dvss.n1713 dvss 0.00541573
R9110 dvss.n3448 dvss 0.00541573
R9111 dvss dvss.n3500 0.00541573
R9112 dvss.n3567 dvss 0.00541573
R9113 dvss dvss.n3616 0.00541573
R9114 dvss.n3680 dvss 0.00541573
R9115 dvss dvss.n3732 0.00541573
R9116 dvss dvss.n3866 0.00541573
R9117 dvss.n3844 dvss 0.00541573
R9118 dvss dvss.n4122 0.00541573
R9119 dvss.n4100 dvss 0.00541573
R9120 dvss dvss.n1172 0.00506461
R9121 dvss dvss.n631 0.00506461
R9122 dvss dvss.n713 0.00506461
R9123 dvss.n1468 dvss 0.00506461
R9124 dvss dvss.n1559 0.00506461
R9125 dvss.n1745 dvss 0.00506461
R9126 dvss dvss.n1707 0.00506461
R9127 dvss.n3417 dvss 0.00506461
R9128 dvss dvss.n3510 0.00506461
R9129 dvss.n3539 dvss 0.00506461
R9130 dvss dvss.n3631 0.00506461
R9131 dvss.n3657 dvss 0.00506461
R9132 dvss dvss.n3742 0.00506461
R9133 dvss.n3876 dvss 0.00506461
R9134 dvss dvss.n4143 0.00506461
R9135 dvss.n4132 dvss 0.00506461
R9136 dvss.n4203 dvss 0.00506461
R9137 dvss.n4230 dvss 0.00506461
R9138 dvss.n933 dvss 0.00493548
R9139 dvss.n1331 dvss 0.00493548
R9140 dvss.n1414 dvss 0.00493548
R9141 dvss.n1814 dvss 0.00493548
R9142 dvss.n3363 dvss 0.00493548
R9143 dvss.n3308 dvss 0.00493548
R9144 dvss.n3258 dvss 0.00493548
R9145 dvss.n3945 dvss 0.00493548
R9146 dvss.n4020 dvss 0.00493548
R9147 dvss.n856 dvss.n855 0.00412903
R9148 dvss.n871 dvss.n870 0.00412903
R9149 dvss.n1110 dvss 0.00401124
R9150 dvss.n1167 dvss.n733 0.00401124
R9151 dvss.n1213 dvss 0.00401124
R9152 dvss.n709 dvss.n705 0.00401124
R9153 dvss dvss.n1501 0.00401124
R9154 dvss.n1554 dvss.n522 0.00401124
R9155 dvss.n1733 dvss 0.00401124
R9156 dvss.n1703 dvss.n1699 0.00401124
R9157 dvss dvss.n3452 0.00401124
R9158 dvss.n3505 dvss.n403 0.00401124
R9159 dvss.n3571 dvss 0.00401124
R9160 dvss.n3626 dvss.n335 0.00401124
R9161 dvss.n3684 dvss 0.00401124
R9162 dvss.n3737 dvss.n272 0.00401124
R9163 dvss.n3864 dvss 0.00401124
R9164 dvss.n4139 dvss.n134 0.00401124
R9165 dvss.n4120 dvss 0.00401124
R9166 dvss.n4208 dvss.n87 0.00401124
R9167 dvss.n2704 dvss.n2694 0.00387838
R9168 dvss.n2710 dvss.n2709 0.00387838
R9169 dvss.n2743 dvss.n2733 0.00387838
R9170 dvss.n2749 dvss.n2748 0.00387838
R9171 dvss.n2782 dvss.n2772 0.00387838
R9172 dvss.n2788 dvss.n2787 0.00387838
R9173 dvss.n2821 dvss.n2811 0.00387838
R9174 dvss.n2827 dvss.n2826 0.00387838
R9175 dvss.n2860 dvss.n2850 0.00387838
R9176 dvss.n2866 dvss.n2865 0.00387838
R9177 dvss.n3174 dvss.n3173 0.00387838
R9178 dvss.n3178 dvss.n3177 0.00387838
R9179 dvss.n2018 dvss.n2017 0.00387838
R9180 dvss.n2073 dvss.n2072 0.00387838
R9181 dvss.n116 dvss.n115 0.00387838
R9182 dvss.n4368 dvss.n4367 0.00387838
R9183 dvss.n4332 dvss.n48 0.00387838
R9184 dvss.n4321 dvss.n4320 0.00387838
R9185 dvss.n2255 dvss.n2254 0.00387838
R9186 dvss.n2259 dvss.n2258 0.00387838
R9187 dvss.n855 dvss 0.00372581
R9188 dvss dvss.n871 0.00372581
R9189 dvss dvss.n899 0.00372581
R9190 dvss.n925 dvss 0.00372581
R9191 dvss dvss.n610 0.00372581
R9192 dvss dvss.n601 0.00372581
R9193 dvss.n1361 dvss 0.00372581
R9194 dvss dvss.n1422 0.00372581
R9195 dvss dvss.n490 0.00372581
R9196 dvss dvss.n481 0.00372581
R9197 dvss.n1844 dvss 0.00372581
R9198 dvss dvss.n3371 0.00372581
R9199 dvss.n1875 dvss 0.00372581
R9200 dvss dvss.n3316 0.00372581
R9201 dvss.n1906 dvss 0.00372581
R9202 dvss dvss.n3266 0.00372581
R9203 dvss dvss.n244 0.00372581
R9204 dvss dvss.n235 0.00372581
R9205 dvss.n3970 dvss 0.00372581
R9206 dvss dvss.n4028 0.00372581
R9207 dvss.n1029 dvss.n1028 0.00366011
R9208 dvss.n825 dvss.n815 0.00366011
R9209 dvss.n1345 dvss 0.00332258
R9210 dvss.n820 dvss 0.00330899
R9211 dvss dvss.n766 0.00330899
R9212 dvss dvss.n749 0.00330899
R9213 dvss dvss.n652 0.00330899
R9214 dvss dvss.n718 0.00330899
R9215 dvss.n1530 dvss 0.00330899
R9216 dvss.n1551 dvss 0.00330899
R9217 dvss dvss.n1723 0.00330899
R9218 dvss dvss.n1712 0.00330899
R9219 dvss.n3481 dvss 0.00330899
R9220 dvss.n3502 dvss 0.00330899
R9221 dvss.n3601 dvss 0.00330899
R9222 dvss.n3618 dvss 0.00330899
R9223 dvss.n3717 dvss 0.00330899
R9224 dvss.n3734 dvss 0.00330899
R9225 dvss dvss.n3854 0.00330899
R9226 dvss.n4148 dvss 0.00330899
R9227 dvss dvss.n4110 0.00330899
R9228 dvss.n4191 dvss 0.00330899
R9229 dvss.n2707 dvss 0.00303378
R9230 dvss.n2746 dvss 0.00303378
R9231 dvss.n2785 dvss 0.00303378
R9232 dvss.n2824 dvss 0.00303378
R9233 dvss.n2863 dvss 0.00303378
R9234 dvss dvss.n3180 0.00303378
R9235 dvss dvss.n2004 0.00303378
R9236 dvss dvss.n22 0.00303378
R9237 dvss dvss.n4323 0.00303378
R9238 dvss dvss.n2261 0.00303378
R9239 dvss dvss.n810 0.00295787
R9240 dvss dvss.n814 0.00295787
R9241 dvss.n1110 dvss.n774 0.00295787
R9242 dvss.n736 dvss 0.00295787
R9243 dvss.n1167 dvss 0.00295787
R9244 dvss.n1213 dvss.n642 0.00295787
R9245 dvss.n710 dvss 0.00295787
R9246 dvss.n705 dvss 0.00295787
R9247 dvss.n1501 dvss.n558 0.00295787
R9248 dvss.n525 dvss 0.00295787
R9249 dvss.n1554 dvss 0.00295787
R9250 dvss.n1733 dvss.n1597 0.00295787
R9251 dvss.n1704 dvss 0.00295787
R9252 dvss.n1699 dvss 0.00295787
R9253 dvss.n3452 dvss.n439 0.00295787
R9254 dvss.n406 dvss 0.00295787
R9255 dvss.n3505 dvss 0.00295787
R9256 dvss.n3572 dvss.n3571 0.00295787
R9257 dvss.n338 dvss 0.00295787
R9258 dvss.n3626 dvss 0.00295787
R9259 dvss.n3685 dvss.n3684 0.00295787
R9260 dvss.n275 dvss 0.00295787
R9261 dvss.n3737 dvss 0.00295787
R9262 dvss.n3864 dvss.n3780 0.00295787
R9263 dvss.n4140 dvss 0.00295787
R9264 dvss dvss.n134 0.00295787
R9265 dvss.n4120 dvss.n154 0.00295787
R9266 dvss.n90 dvss 0.00295787
R9267 dvss dvss.n4208 0.00295787
R9268 dvss.n910 dvss 0.00291935
R9269 dvss.n933 dvss.n928 0.00291935
R9270 dvss.n1297 dvss 0.00291935
R9271 dvss.n1332 dvss.n1331 0.00291935
R9272 dvss.n1440 dvss 0.00291935
R9273 dvss.n1414 dvss.n1371 0.00291935
R9274 dvss.n1780 dvss 0.00291935
R9275 dvss.n1815 dvss.n1814 0.00291935
R9276 dvss.n3389 dvss 0.00291935
R9277 dvss.n3363 dvss.n1854 0.00291935
R9278 dvss.n3334 dvss 0.00291935
R9279 dvss.n3308 dvss.n1885 0.00291935
R9280 dvss.n3284 dvss 0.00291935
R9281 dvss.n3258 dvss.n1916 0.00291935
R9282 dvss.n3911 dvss 0.00291935
R9283 dvss.n3946 dvss.n3945 0.00291935
R9284 dvss.n4046 dvss 0.00291935
R9285 dvss.n4020 dvss.n3996 0.00291935
R9286 dvss.n820 dvss 0.00260674
R9287 dvss.n1131 dvss 0.00260674
R9288 dvss.n1191 dvss.n736 0.00260674
R9289 dvss.n1226 dvss 0.00260674
R9290 dvss.n710 dvss.n675 0.00260674
R9291 dvss.n1514 dvss 0.00260674
R9292 dvss.n1578 dvss.n525 0.00260674
R9293 dvss dvss.n1728 0.00260674
R9294 dvss.n1704 dvss.n1630 0.00260674
R9295 dvss.n3465 dvss 0.00260674
R9296 dvss.n3530 dvss.n406 0.00260674
R9297 dvss.n3587 dvss 0.00260674
R9298 dvss.n3647 dvss.n338 0.00260674
R9299 dvss.n3690 dvss 0.00260674
R9300 dvss.n3761 dvss.n275 0.00260674
R9301 dvss dvss.n3859 0.00260674
R9302 dvss.n4140 dvss.n133 0.00260674
R9303 dvss dvss.n4115 0.00260674
R9304 dvss.n4212 dvss.n90 0.00260674
R9305 dvss.n1192 dvss.n1191 0.00190449
R9306 dvss.n1195 dvss.n631 0.00190449
R9307 dvss.n707 dvss.n675 0.00190449
R9308 dvss.n1468 dvss.n1467 0.00190449
R9309 dvss.n1579 dvss.n1578 0.00190449
R9310 dvss.n1745 dvss.n512 0.00190449
R9311 dvss.n1701 dvss.n1630 0.00190449
R9312 dvss.n3417 dvss.n3416 0.00190449
R9313 dvss.n3531 dvss.n3530 0.00190449
R9314 dvss.n3539 dvss.n392 0.00190449
R9315 dvss.n3648 dvss.n3647 0.00190449
R9316 dvss.n3657 dvss.n330 0.00190449
R9317 dvss.n3762 dvss.n3761 0.00190449
R9318 dvss.n3876 dvss.n267 0.00190449
R9319 dvss.n4137 dvss.n133 0.00190449
R9320 dvss.n4133 dvss.n4132 0.00190449
R9321 dvss.n4213 dvss.n4212 0.00190449
R9322 dvss.n4230 dvss.n73 0.00190449
R9323 dvss dvss.n1408 0.00170968
R9324 dvss.n1828 dvss 0.00170968
R9325 dvss dvss.n3357 0.00170968
R9326 dvss.n1157 dvss.n1156 0.00155337
R9327 dvss dvss.n1197 0.00155337
R9328 dvss.n719 dvss.n663 0.00155337
R9329 dvss dvss.n578 0.00155337
R9330 dvss.n1465 dvss 0.00155337
R9331 dvss.n1549 dvss.n538 0.00155337
R9332 dvss dvss.n519 0.00155337
R9333 dvss dvss.n1583 0.00155337
R9334 dvss.n1713 dvss.n1617 0.00155337
R9335 dvss dvss.n458 0.00155337
R9336 dvss.n3414 dvss 0.00155337
R9337 dvss.n3500 dvss.n419 0.00155337
R9338 dvss dvss.n400 0.00155337
R9339 dvss dvss.n3535 0.00155337
R9340 dvss.n3616 dvss.n354 0.00155337
R9341 dvss dvss.n3652 0.00155337
R9342 dvss.n3732 dvss.n288 0.00155337
R9343 dvss dvss.n3766 0.00155337
R9344 dvss.n3844 dvss.n3843 0.00155337
R9345 dvss dvss.n138 0.00155337
R9346 dvss.n4100 dvss.n4099 0.00155337
R9347 dvss dvss.n4217 0.00155337
R9348 dvss.n2663 dvss.n2662 0.00134459
R9349 dvss.n2548 dvss.n2129 0.00134459
R9350 dvss dvss.n2534 0.00134459
R9351 dvss.n868 dvss 0.00130645
R9352 dvss dvss.n819 0.00120225
R9353 dvss.n922 dvss.n921 0.000903226
R9354 dvss.n938 dvss 0.000903226
R9355 dvss.n1317 dvss.n600 0.000903226
R9356 dvss dvss.n593 0.000903226
R9357 dvss.n1426 dvss.n1365 0.000903226
R9358 dvss dvss.n1412 0.000903226
R9359 dvss.n1800 dvss.n480 0.000903226
R9360 dvss dvss.n473 0.000903226
R9361 dvss.n3375 dvss.n1848 0.000903226
R9362 dvss dvss.n3361 0.000903226
R9363 dvss.n3320 dvss.n1879 0.000903226
R9364 dvss dvss.n3306 0.000903226
R9365 dvss.n3270 dvss.n1910 0.000903226
R9366 dvss dvss.n3256 0.000903226
R9367 dvss.n3931 dvss.n234 0.000903226
R9368 dvss dvss.n227 0.000903226
R9369 dvss.n4032 dvss.n3990 0.000903226
R9370 dvss dvss.n4018 0.000903226
R9371 dvss.n1022 dvss.n1021 0.000851124
R9372 dvss.n1023 dvss.n805 0.000851124
R9373 dvss.n1024 dvss.n806 0.000851124
R9374 dvss.n1025 dvss.n807 0.000851124
R9375 dvss.n1026 dvss.n808 0.000851124
R9376 dvss.n1027 dvss.n809 0.000851124
R9377 dvss.n1028 dvss.n810 0.000851124
R9378 dvss.n1032 dvss.n811 0.000851124
R9379 dvss.n1033 dvss.n812 0.000851124
R9380 dvss.n1034 dvss.n813 0.000851124
R9381 dvss.n825 dvss.n814 0.000851124
R9382 dvss.n1070 dvss.n1056 0.000851124
R9383 dvss.n1069 dvss.n1068 0.000851124
R9384 dvss.n1067 dvss.n1057 0.000851124
R9385 dvss.n1059 dvss.n785 0.000851124
R9386 dvss.n1065 dvss.n1064 0.000851124
R9387 dvss.n1098 dvss.n1097 0.000851124
R9388 dvss.n788 dvss.n787 0.000851124
R9389 dvss.n1158 dvss.n753 0.000851124
R9390 dvss.n1188 dvss 0.000851124
R9391 dvss.n1237 dvss.n662 0.000851124
R9392 dvss dvss.n704 0.000851124
R9393 dvss.n1547 dvss.n1546 0.000851124
R9394 dvss.n1575 dvss 0.000851124
R9395 dvss.n1718 dvss.n1616 0.000851124
R9396 dvss dvss.n1698 0.000851124
R9397 dvss.n3498 dvss.n3497 0.000851124
R9398 dvss.n3527 dvss 0.000851124
R9399 dvss.n3614 dvss.n3613 0.000851124
R9400 dvss.n3644 dvss 0.000851124
R9401 dvss.n3730 dvss.n3729 0.000851124
R9402 dvss.n3758 dvss 0.000851124
R9403 dvss.n3849 dvss.n3842 0.000851124
R9404 dvss.n204 dvss 0.000851124
R9405 dvss.n4105 dvss.n4098 0.000851124
R9406 dvss.n4209 dvss 0.000851124
R9407 avss.n68 avss.n67 2.18688e+07
R9408 avss.n370 avss.n369 188352
R9409 avss.n882 avss.n846 160432
R9410 avss.n845 avss.n844 110146
R9411 avss.n66 avss.n50 100279
R9412 avss.n1013 avss.n50 100279
R9413 avss.n66 avss.n51 100279
R9414 avss.n1013 avss.n51 100279
R9415 avss.n369 avss.n368 92956.3
R9416 avss.n308 avss.n69 68021.9
R9417 avss.n997 avss.n363 64733.3
R9418 avss.n369 avss.t273 48414.6
R9419 avss.n871 avss.n360 45524.4
R9420 avss.n871 avss.n361 45524.4
R9421 avss.n999 avss.n360 45524.4
R9422 avss.n999 avss.n361 45524.4
R9423 avss.n577 avss.n573 45524.4
R9424 avss.n777 avss.n573 45524.4
R9425 avss.n776 avss.n577 45524.4
R9426 avss.n777 avss.n776 45524.4
R9427 avss.n308 avss.n307 45183
R9428 avss.n1096 avss.n8 37415.6
R9429 avss.n997 avss.n996 29160.7
R9430 avss.n846 avss.t384 29031.2
R9431 avss.n1016 avss.n47 21059.4
R9432 avss.n1016 avss.n48 21059.4
R9433 avss.n1018 avss.n47 21059.4
R9434 avss.n1018 avss.n48 21059.4
R9435 avss.n982 avss.n372 18174.6
R9436 avss.n989 avss.n372 18174.6
R9437 avss.n989 avss.n371 18174.6
R9438 avss.n982 avss.n371 18174.6
R9439 avss.n828 avss.n553 18174.6
R9440 avss.n800 avss.n553 18174.6
R9441 avss.n828 avss.n827 18174.6
R9442 avss.n827 avss.n800 18174.6
R9443 avss.n843 avss.n564 17601.7
R9444 avss.n344 avss.n63 16300.9
R9445 avss.n340 avss.n63 16300.9
R9446 avss.n344 avss.n65 16300.9
R9447 avss.n340 avss.n65 16300.9
R9448 avss.n883 avss.n882 13864
R9449 avss.n117 avss.n69 12588.9
R9450 avss.n880 avss.n848 12517.1
R9451 avss.n874 avss.n848 12517.1
R9452 avss.n874 avss.n847 12517.1
R9453 avss.n880 avss.n847 12517.1
R9454 avss.n443 avss.n439 7742.83
R9455 avss.n445 avss.n439 7742.83
R9456 avss.n444 avss.n443 7742.83
R9457 avss.n445 avss.n444 7742.83
R9458 avss.n861 avss.n19 7610.36
R9459 avss.n861 avss.n20 7610.36
R9460 avss.n1073 avss.n20 7610.36
R9461 avss.n1073 avss.n19 7610.36
R9462 avss.n846 avss.n845 7383.98
R9463 avss.n54 avss.n52 6515.58
R9464 avss.n1012 avss.n52 6515.58
R9465 avss.n1011 avss.n54 6515.58
R9466 avss.n1012 avss.n1011 6515.58
R9467 avss.n1076 avss.n12 5644.38
R9468 avss.n1076 avss.n13 5644.38
R9469 avss.n1087 avss.n13 5644.38
R9470 avss.n1087 avss.n12 5644.38
R9471 avss.n69 avss.n68 4523.98
R9472 avss.n442 avss.n437 4175.68
R9473 avss.n446 avss.n437 4175.68
R9474 avss.n442 avss.n438 4175.68
R9475 avss.n446 avss.n438 4175.68
R9476 avss.n976 avss.n379 4139.43
R9477 avss.n972 avss.n379 4139.43
R9478 avss.n976 avss.n380 4139.43
R9479 avss.n972 avss.n380 4139.43
R9480 avss.n832 avss.n793 4139.43
R9481 avss.n798 avss.n793 4139.43
R9482 avss.n798 avss.n794 4139.43
R9483 avss.n832 avss.n794 4139.43
R9484 avss.n561 avss.n557 3978.07
R9485 avss.n561 avss.n558 3978.07
R9486 avss.n886 avss.n558 3978.07
R9487 avss.n886 avss.n557 3978.07
R9488 avss.n995 avss.n365 3978.07
R9489 avss.n991 avss.n365 3978.07
R9490 avss.n991 avss.n364 3978.07
R9491 avss.n995 avss.n364 3978.07
R9492 avss.t282 avss.t171 3966.94
R9493 avss.t280 avss.t282 3966.94
R9494 avss.t278 avss.t284 3966.94
R9495 avss.t284 avss.t193 3966.94
R9496 avss.n845 avss.n843 3945.98
R9497 avss.n1090 avss.n9 3902.33
R9498 avss.n1090 avss.n10 3902.33
R9499 avss.n1094 avss.n10 3902.33
R9500 avss.n1094 avss.n9 3902.33
R9501 avss.n882 avss.n881 3318.88
R9502 avss.n322 avss.n321 2998.14
R9503 avss.n1000 avss.n359 2957.93
R9504 avss.n778 avss.n571 2957.93
R9505 avss.n576 avss.n572 2957.93
R9506 avss.n778 avss.n572 2957.93
R9507 avss.n576 avss.n574 2940.24
R9508 avss.n870 avss.n359 2935.34
R9509 avss.n129 avss.n128 2905.02
R9510 avss.n141 avss.n140 2905.02
R9511 avss.n153 avss.n152 2905.02
R9512 avss.n165 avss.n164 2905.02
R9513 avss.n177 avss.n176 2905.02
R9514 avss.n189 avss.n188 2905.02
R9515 avss.n201 avss.n200 2905.02
R9516 avss.n213 avss.n212 2905.02
R9517 avss.n225 avss.n224 2905.02
R9518 avss.n237 avss.n236 2905.02
R9519 avss.n249 avss.n248 2905.02
R9520 avss.n261 avss.n260 2905.02
R9521 avss.n273 avss.n272 2905.02
R9522 avss.n285 avss.n284 2905.02
R9523 avss.n297 avss.n296 2905.02
R9524 avss.n1098 avss.n1097 2538.7
R9525 avss.t39 avss.n793 2436.62
R9526 avss.n794 avss.t384 2436.62
R9527 avss.n379 avss.t52 2436.62
R9528 avss.n1019 avss.n45 2366.87
R9529 avss.n1019 avss.n44 2366.87
R9530 avss.n1015 avss.n44 2344.28
R9531 avss.n1015 avss.n45 2344.28
R9532 avss.n829 avss.t171 2304.08
R9533 avss.t193 avss.n562 2304.08
R9534 avss.n489 avss.n473 2087.09
R9535 avss.n514 avss.n463 2084.98
R9536 avss.n825 avss.n552 2054.02
R9537 avss.n890 avss.n552 2054.02
R9538 avss.n988 avss.n373 2054.02
R9539 avss.n983 avss.n373 2054.02
R9540 avss.n507 avss.n505 2039.85
R9541 avss.n531 avss.n530 2039.84
R9542 avss.n826 avss.t280 1983.47
R9543 avss.n826 avss.t278 1983.47
R9544 avss.n890 avss.n889 1894.78
R9545 avss.n825 avss.n801 1894.78
R9546 avss.n985 avss.n983 1894.78
R9547 avss.n988 avss.n987 1894.78
R9548 avss.n339 avss.n338 1813.84
R9549 avss.n1100 avss.n6 1735.47
R9550 avss.n1101 avss.n6 1735.47
R9551 avss.n1101 avss.n5 1735.47
R9552 avss.n1100 avss.n5 1735.47
R9553 avss.t46 avss.n49 1637.21
R9554 avss.n346 avss.n62 1602.64
R9555 avss.n864 avss.n863 1487.81
R9556 avss.n863 avss.n357 1487.81
R9557 avss.n870 avss.n864 1439.24
R9558 avss.n1000 avss.n357 1439.24
R9559 avss.n875 avss.n860 1435.48
R9560 avss.n875 avss.n859 1435.48
R9561 avss.n321 avss.n320 1414.29
R9562 avss.t174 avss.t231 1389.88
R9563 avss.n879 avss.n850 1385.79
R9564 avss.n879 avss.n849 1385.79
R9565 avss.n831 avss.t27 1301
R9566 avss.n831 avss.t31 1301
R9567 avss.n977 avss.t48 1301
R9568 avss.t58 avss.n977 1301
R9569 avss.n996 avss.t231 1143.92
R9570 avss.t31 avss.t37 1081.77
R9571 avss.t52 avss.t44 1081.77
R9572 avss.t29 avss.t39 1081.77
R9573 avss.t33 avss.t29 1081.77
R9574 avss.t35 avss.t33 1081.77
R9575 avss.t27 avss.t35 1081.77
R9576 avss.t37 avss.t25 1081.77
R9577 avss.t25 avss.t382 1081.77
R9578 avss.t44 avss.t56 1081.77
R9579 avss.t56 avss.t54 1081.77
R9580 avss.n441 avss.n434 976.942
R9581 avss.n441 avss.n440 976.942
R9582 avss.n448 avss.n447 976.188
R9583 avss.n447 avss.n436 974.683
R9584 avss.t271 avss.n49 964.784
R9585 avss.n321 avss.n308 939.895
R9586 avss.n799 avss.t27 925.769
R9587 avss.t31 avss.n799 925.769
R9588 avss.n830 avss.t384 887.293
R9589 avss.n1072 avss.n21 874.542
R9590 avss.n22 avss.n21 874.542
R9591 avss.n128 avss.n115 815.444
R9592 avss.n140 avss.n112 815.444
R9593 avss.n152 avss.n109 815.444
R9594 avss.n164 avss.n106 815.444
R9595 avss.n176 avss.n103 815.444
R9596 avss.n188 avss.n100 815.444
R9597 avss.n200 avss.n97 815.444
R9598 avss.n212 avss.n94 815.444
R9599 avss.n224 avss.n91 815.444
R9600 avss.n236 avss.n88 815.444
R9601 avss.n248 avss.n85 815.444
R9602 avss.n260 avss.n82 815.444
R9603 avss.n272 avss.n79 815.444
R9604 avss.n284 avss.n76 815.444
R9605 avss.n296 avss.n73 815.444
R9606 avss.n307 avss.n70 815.444
R9607 avss.n59 avss.n58 796.612
R9608 avss.n64 avss.n58 782.683
R9609 avss.n312 avss.n309 769.572
R9610 avss.n1070 avss.n1069 765.741
R9611 avss.n1071 avss.n1070 765.741
R9612 avss.n56 avss.n55 759.718
R9613 avss.n117 avss.t267 755.986
R9614 avss.n129 avss.t95 755.986
R9615 avss.n141 avss.t245 755.986
R9616 avss.n153 avss.t22 755.986
R9617 avss.n165 avss.t73 755.986
R9618 avss.n177 avss.t378 755.986
R9619 avss.n189 avss.t17 755.986
R9620 avss.n201 avss.t376 755.986
R9621 avss.n213 avss.t100 755.986
R9622 avss.n225 avss.t306 755.986
R9623 avss.n237 avss.t396 755.986
R9624 avss.n249 avss.t78 755.986
R9625 avss.n261 avss.t253 755.986
R9626 avss.n273 avss.t340 755.986
R9627 avss.n285 avss.t300 755.986
R9628 avss.n297 avss.t311 755.986
R9629 avss.t327 avss.t325 731.963
R9630 avss.t286 avss.t290 731.963
R9631 avss.t290 avss.n884 684.673
R9632 avss.n885 avss.t325 668.225
R9633 avss.n1086 avss.n14 649.788
R9634 avss.n1077 avss.n14 649.788
R9635 avss.n998 avss.n997 627.813
R9636 avss.n506 avss.t169 625.516
R9637 avss.n513 avss.t169 625.516
R9638 avss.t169 avss.n457 614.321
R9639 avss.n524 avss.t169 614.321
R9640 avss.n844 avss.t327 602.431
R9641 avss.n57 avss.n56 598.966
R9642 avss.t169 avss.n496 598.606
R9643 avss.n497 avss.t169 598.606
R9644 avss.n482 avss.t169 588.343
R9645 avss.n480 avss.t169 588.343
R9646 avss.n319 avss.n318 585
R9647 avss.n320 avss.n319 585
R9648 avss.n311 avss.n310 585
R9649 avss.n503 avss.n502 585
R9650 avss.n501 avss.n470 585
R9651 avss.n470 avss.n469 585
R9652 avss.n500 avss.n499 585
R9653 avss.n499 avss.n498 585
R9654 avss.n472 avss.n471 585
R9655 avss.n497 avss.n472 585
R9656 avss.n495 avss.n494 585
R9657 avss.n496 avss.n495 585
R9658 avss.n493 avss.n474 585
R9659 avss.n474 avss.n473 585
R9660 avss.n492 avss.n491 585
R9661 avss.n476 avss.n475 585
R9662 avss.n518 avss.n517 585
R9663 avss.n515 avss.n465 585
R9664 avss.n515 avss.n514 585
R9665 avss.n512 avss.n511 585
R9666 avss.n513 avss.n512 585
R9667 avss.n510 avss.n466 585
R9668 avss.n506 avss.n466 585
R9669 avss.n509 avss.n508 585
R9670 avss.n508 avss.n507 585
R9671 avss.n468 avss.n467 585
R9672 avss.n519 avss.n464 585
R9673 avss.n521 avss.n520 585
R9674 avss.n522 avss.n521 585
R9675 avss.n462 avss.n461 585
R9676 avss.n523 avss.n462 585
R9677 avss.n526 avss.n525 585
R9678 avss.n525 avss.n524 585
R9679 avss.n527 avss.n459 585
R9680 avss.n459 avss.n457 585
R9681 avss.n529 avss.n528 585
R9682 avss.n530 avss.n529 585
R9683 avss.n460 avss.n458 585
R9684 avss.n454 avss.n452 585
R9685 avss.n487 avss.n486 585
R9686 avss.n488 avss.n487 585
R9687 avss.n485 avss.n478 585
R9688 avss.n478 avss.n477 585
R9689 avss.n484 avss.n483 585
R9690 avss.n483 avss.n482 585
R9691 avss.n481 avss.n479 585
R9692 avss.n481 avss.n480 585
R9693 avss.n453 avss.n451 585
R9694 avss.n455 avss.n453 585
R9695 avss.n534 avss.n533 585
R9696 avss.n533 avss.n532 585
R9697 avss.n635 avss.n634 585
R9698 avss.n634 avss.n633 585
R9699 avss.n641 avss.n640 585
R9700 avss.n642 avss.n641 585
R9701 avss.n632 avss.n631 585
R9702 avss.n643 avss.n632 585
R9703 avss.n647 avss.n646 585
R9704 avss.n646 avss.n645 585
R9705 avss.n627 avss.n626 585
R9706 avss.n644 avss.n626 585
R9707 avss.n655 avss.n654 585
R9708 avss.n656 avss.n655 585
R9709 avss.n624 avss.n622 585
R9710 avss.n657 avss.n624 585
R9711 avss.n662 avss.n661 585
R9712 avss.n661 avss.n660 585
R9713 avss.n625 avss.n623 585
R9714 avss.n659 avss.n625 585
R9715 avss.n618 avss.n617 585
R9716 avss.n658 avss.n617 585
R9717 avss.n675 avss.n674 585
R9718 avss.n676 avss.n675 585
R9719 avss.n616 avss.n615 585
R9720 avss.n677 avss.n616 585
R9721 avss.n681 avss.n680 585
R9722 avss.n680 avss.n679 585
R9723 avss.n611 avss.n610 585
R9724 avss.n678 avss.n610 585
R9725 avss.n696 avss.n695 585
R9726 avss.n697 avss.n696 585
R9727 avss.n694 avss.n608 585
R9728 avss.n698 avss.n608 585
R9729 avss.n700 avss.n609 585
R9730 avss.n700 avss.n699 585
R9731 avss.n701 avss.n607 585
R9732 avss.n702 avss.n701 585
R9733 avss.n706 avss.n705 585
R9734 avss.n705 avss.n704 585
R9735 avss.n605 avss.n604 585
R9736 avss.n703 avss.n604 585
R9737 avss.n716 avss.n715 585
R9738 avss.n717 avss.n716 585
R9739 avss.n603 avss.n602 585
R9740 avss.n718 avss.n603 585
R9741 avss.n722 avss.n721 585
R9742 avss.n721 avss.n720 585
R9743 avss.n598 avss.n597 585
R9744 avss.n719 avss.n597 585
R9745 avss.n730 avss.n729 585
R9746 avss.n731 avss.n730 585
R9747 avss.n596 avss.n595 585
R9748 avss.n732 avss.n596 585
R9749 avss.n736 avss.n735 585
R9750 avss.n735 avss.n734 585
R9751 avss.n592 avss.n591 585
R9752 avss.n733 avss.n591 585
R9753 avss.n744 avss.n743 585
R9754 avss.n745 avss.n744 585
R9755 avss.n590 avss.n589 585
R9756 avss.n746 avss.n590 585
R9757 avss.n750 avss.n749 585
R9758 avss.n749 avss.n748 585
R9759 avss.n586 avss.n585 585
R9760 avss.n747 avss.n585 585
R9761 avss.n760 avss.n759 585
R9762 avss.n761 avss.n760 585
R9763 avss.n584 avss.n583 585
R9764 avss.n762 avss.n584 585
R9765 avss.n765 avss.n764 585
R9766 avss.n764 avss.n763 585
R9767 avss.n580 avss.n579 585
R9768 avss.n579 avss.n578 585
R9769 avss.n773 avss.n772 585
R9770 avss.n774 avss.n773 585
R9771 avss.n567 avss.n566 585
R9772 avss.n566 avss.n565 585
R9773 avss.n841 avss.n840 585
R9774 avss.n842 avss.n841 585
R9775 avss.n119 avss.n118 585
R9776 avss.n118 avss.n117 585
R9777 avss.n120 avss.n116 585
R9778 avss.n116 avss.n115 585
R9779 avss.n127 avss.n126 585
R9780 avss.n128 avss.n127 585
R9781 avss.n131 avss.n130 585
R9782 avss.n130 avss.n129 585
R9783 avss.n114 avss.n113 585
R9784 avss.n113 avss.n112 585
R9785 avss.n139 avss.n138 585
R9786 avss.n140 avss.n139 585
R9787 avss.n143 avss.n142 585
R9788 avss.n142 avss.n141 585
R9789 avss.n111 avss.n110 585
R9790 avss.n110 avss.n109 585
R9791 avss.n151 avss.n150 585
R9792 avss.n152 avss.n151 585
R9793 avss.n155 avss.n154 585
R9794 avss.n154 avss.n153 585
R9795 avss.n108 avss.n107 585
R9796 avss.n107 avss.n106 585
R9797 avss.n163 avss.n162 585
R9798 avss.n164 avss.n163 585
R9799 avss.n167 avss.n166 585
R9800 avss.n166 avss.n165 585
R9801 avss.n105 avss.n104 585
R9802 avss.n104 avss.n103 585
R9803 avss.n175 avss.n174 585
R9804 avss.n176 avss.n175 585
R9805 avss.n179 avss.n178 585
R9806 avss.n178 avss.n177 585
R9807 avss.n102 avss.n101 585
R9808 avss.n101 avss.n100 585
R9809 avss.n187 avss.n186 585
R9810 avss.n188 avss.n187 585
R9811 avss.n191 avss.n190 585
R9812 avss.n190 avss.n189 585
R9813 avss.n99 avss.n98 585
R9814 avss.n98 avss.n97 585
R9815 avss.n199 avss.n198 585
R9816 avss.n200 avss.n199 585
R9817 avss.n203 avss.n202 585
R9818 avss.n202 avss.n201 585
R9819 avss.n96 avss.n95 585
R9820 avss.n95 avss.n94 585
R9821 avss.n211 avss.n210 585
R9822 avss.n212 avss.n211 585
R9823 avss.n215 avss.n214 585
R9824 avss.n214 avss.n213 585
R9825 avss.n93 avss.n92 585
R9826 avss.n92 avss.n91 585
R9827 avss.n223 avss.n222 585
R9828 avss.n224 avss.n223 585
R9829 avss.n227 avss.n226 585
R9830 avss.n226 avss.n225 585
R9831 avss.n90 avss.n89 585
R9832 avss.n89 avss.n88 585
R9833 avss.n235 avss.n234 585
R9834 avss.n236 avss.n235 585
R9835 avss.n239 avss.n238 585
R9836 avss.n238 avss.n237 585
R9837 avss.n87 avss.n86 585
R9838 avss.n86 avss.n85 585
R9839 avss.n247 avss.n246 585
R9840 avss.n248 avss.n247 585
R9841 avss.n251 avss.n250 585
R9842 avss.n250 avss.n249 585
R9843 avss.n84 avss.n83 585
R9844 avss.n83 avss.n82 585
R9845 avss.n259 avss.n258 585
R9846 avss.n260 avss.n259 585
R9847 avss.n263 avss.n262 585
R9848 avss.n262 avss.n261 585
R9849 avss.n81 avss.n80 585
R9850 avss.n80 avss.n79 585
R9851 avss.n271 avss.n270 585
R9852 avss.n272 avss.n271 585
R9853 avss.n275 avss.n274 585
R9854 avss.n274 avss.n273 585
R9855 avss.n78 avss.n77 585
R9856 avss.n77 avss.n76 585
R9857 avss.n283 avss.n282 585
R9858 avss.n284 avss.n283 585
R9859 avss.n287 avss.n286 585
R9860 avss.n286 avss.n285 585
R9861 avss.n75 avss.n74 585
R9862 avss.n74 avss.n73 585
R9863 avss.n295 avss.n294 585
R9864 avss.n296 avss.n295 585
R9865 avss.n299 avss.n298 585
R9866 avss.n298 avss.n297 585
R9867 avss.n72 avss.n71 585
R9868 avss.n71 avss.n70 585
R9869 avss.n306 avss.n305 585
R9870 avss.n307 avss.n306 585
R9871 avss.n1078 avss.n15 540.989
R9872 avss.n1085 avss.n15 540.989
R9873 avss.n319 avss.n310 539.294
R9874 avss.n641 avss.n634 539.294
R9875 avss.n641 avss.n632 539.294
R9876 avss.n646 avss.n632 539.294
R9877 avss.n646 avss.n626 539.294
R9878 avss.n655 avss.n626 539.294
R9879 avss.n655 avss.n624 539.294
R9880 avss.n661 avss.n624 539.294
R9881 avss.n661 avss.n625 539.294
R9882 avss.n625 avss.n617 539.294
R9883 avss.n675 avss.n617 539.294
R9884 avss.n675 avss.n616 539.294
R9885 avss.n680 avss.n616 539.294
R9886 avss.n680 avss.n610 539.294
R9887 avss.n696 avss.n610 539.294
R9888 avss.n696 avss.n608 539.294
R9889 avss.n700 avss.n608 539.294
R9890 avss.n701 avss.n700 539.294
R9891 avss.n705 avss.n701 539.294
R9892 avss.n705 avss.n604 539.294
R9893 avss.n716 avss.n604 539.294
R9894 avss.n716 avss.n603 539.294
R9895 avss.n721 avss.n603 539.294
R9896 avss.n721 avss.n597 539.294
R9897 avss.n730 avss.n597 539.294
R9898 avss.n730 avss.n596 539.294
R9899 avss.n735 avss.n596 539.294
R9900 avss.n735 avss.n591 539.294
R9901 avss.n744 avss.n591 539.294
R9902 avss.n744 avss.n590 539.294
R9903 avss.n749 avss.n590 539.294
R9904 avss.n749 avss.n585 539.294
R9905 avss.n760 avss.n585 539.294
R9906 avss.n760 avss.n584 539.294
R9907 avss.n764 avss.n584 539.294
R9908 avss.n764 avss.n579 539.294
R9909 avss.n773 avss.n579 539.294
R9910 avss.n773 avss.n566 539.294
R9911 avss.n841 avss.n566 539.294
R9912 avss.n298 avss.n71 539.294
R9913 avss.n306 avss.n71 539.294
R9914 avss.n286 avss.n74 539.294
R9915 avss.n295 avss.n74 539.294
R9916 avss.n274 avss.n77 539.294
R9917 avss.n283 avss.n77 539.294
R9918 avss.n262 avss.n80 539.294
R9919 avss.n271 avss.n80 539.294
R9920 avss.n250 avss.n83 539.294
R9921 avss.n259 avss.n83 539.294
R9922 avss.n238 avss.n86 539.294
R9923 avss.n247 avss.n86 539.294
R9924 avss.n226 avss.n89 539.294
R9925 avss.n235 avss.n89 539.294
R9926 avss.n214 avss.n92 539.294
R9927 avss.n223 avss.n92 539.294
R9928 avss.n202 avss.n95 539.294
R9929 avss.n211 avss.n95 539.294
R9930 avss.n190 avss.n98 539.294
R9931 avss.n199 avss.n98 539.294
R9932 avss.n178 avss.n101 539.294
R9933 avss.n187 avss.n101 539.294
R9934 avss.n166 avss.n104 539.294
R9935 avss.n175 avss.n104 539.294
R9936 avss.n154 avss.n107 539.294
R9937 avss.n163 avss.n107 539.294
R9938 avss.n142 avss.n110 539.294
R9939 avss.n151 avss.n110 539.294
R9940 avss.n130 avss.n113 539.294
R9941 avss.n139 avss.n113 539.294
R9942 avss.n118 avss.n116 539.294
R9943 avss.n127 avss.n116 539.294
R9944 avss.n321 avss.t330 492.382
R9945 avss.n378 avss.t174 488.039
R9946 avss.n797 avss.n792 477.741
R9947 avss.n833 avss.n792 477.741
R9948 avss.n974 avss.n973 477.741
R9949 avss.n975 avss.n974 477.741
R9950 avss.t288 avss.n883 474.954
R9951 avss.n887 avss.n556 459.295
R9952 avss.n560 avss.n556 459.295
R9953 avss.n560 avss.n559 459.295
R9954 avss.n994 avss.n366 459.295
R9955 avss.n994 avss.n993 459.295
R9956 avss.n993 avss.n992 459.295
R9957 avss.n483 avss.n481 456.416
R9958 avss.n525 avss.n459 456.416
R9959 avss.n512 avss.n466 456.416
R9960 avss.n495 avss.n472 456.416
R9961 avss.n1093 avss.n11 425.264
R9962 avss.n1091 avss.n11 420.43
R9963 avss.n1092 avss.n1091 420.43
R9964 avss.n1093 avss.n1092 420.43
R9965 avss.n834 avss.n791 401.812
R9966 avss.n796 avss.n791 401.812
R9967 avss.n382 avss.n381 401.812
R9968 avss.n971 avss.n382 401.812
R9969 avss.n25 avss.t140 392.769
R9970 avss.n24 avss.t213 392.692
R9971 avss.n23 avss.t185 392.664
R9972 avss.n61 avss.t149 384.515
R9973 avss.n323 avss.t209 384.515
R9974 avss.n325 avss.t205 384.515
R9975 avss.n326 avss.t211 384.515
R9976 avss.n327 avss.t207 384.515
R9977 avss.n328 avss.t183 384.515
R9978 avss.n329 avss.t158 384.515
R9979 avss.n336 avss.t138 384.515
R9980 avss.n334 avss.t160 384.515
R9981 avss.n333 avss.t142 384.515
R9982 avss.n332 avss.t196 384.515
R9983 avss.n331 avss.t156 384.515
R9984 avss.n330 avss.t187 384.515
R9985 avss.n324 avss.t215 384.454
R9986 avss.n335 avss.t151 384.454
R9987 avss.n872 avss.t128 382.757
R9988 avss.n507 avss.n506 363.548
R9989 avss.n514 avss.n513 363.548
R9990 avss.n530 avss.n457 357.041
R9991 avss.n524 avss.n523 357.041
R9992 avss.n523 avss.n522 357.041
R9993 avss.n522 avss.n463 357.041
R9994 avss.n496 avss.n473 347.908
R9995 avss.n498 avss.n497 347.908
R9996 avss.n498 avss.n469 347.908
R9997 avss.n505 avss.n469 347.908
R9998 avss.n489 avss.n488 341.943
R9999 avss.n488 avss.n477 341.943
R10000 avss.n482 avss.n477 341.943
R10001 avss.n480 avss.n455 341.943
R10002 avss.n532 avss.n455 341.943
R10003 avss.n532 avss.n531 341.943
R10004 avss.n830 avss.n829 340.805
R10005 avss.n363 avss.t0 338.375
R10006 avss.n419 avss.n406 333.334
R10007 avss.n414 avss.n413 333.334
R10008 avss.n429 avss.n404 333.334
R10009 avss.t296 avss.n7 323.332
R10010 avss.t296 avss.n1098 323.332
R10011 avss.n888 avss.n555 318.495
R10012 avss.n984 avss.n367 318.495
R10013 avss.n321 avss.n7 301.202
R10014 avss.n516 avss.n463 283.521
R10015 avss.n505 avss.n504 283.521
R10016 avss.n339 avss.n55 274.072
R10017 avss.n345 avss.n59 270.683
R10018 avss.n881 avss.t67 262.885
R10019 avss.n873 avss.t67 262.885
R10020 avss.n490 avss.n489 262.719
R10021 avss.n531 avss.n456 262.719
R10022 avss.n998 avss.t146 239.365
R10023 avss.n346 avss.n345 238.306
R10024 avss.n884 avss.n562 227.298
R10025 avss.t220 avss.n11 209.756
R10026 avss.n1092 avss.t220 209.756
R10027 avss.n64 avss.n57 208.189
R10028 avss.n1099 avss.n4 202.918
R10029 avss.n1102 avss.n4 202.918
R10030 avss.n320 avss.n309 200.215
R10031 avss.t382 avss.n830 194.476
R10032 avss.n1099 avss.n3 193.918
R10033 avss.n862 avss.t146 188.975
R10034 avss.n1103 avss.n1102 186.73
R10035 avss.t115 avss.t5 185.605
R10036 avss.t5 avss.t320 185.605
R10037 avss.t320 avss.t105 185.605
R10038 avss.t105 avss.t240 185.605
R10039 avss.t240 avss.t11 185.605
R10040 avss.t11 avss.t249 185.605
R10041 avss.t249 avss.t20 185.605
R10042 avss.t20 avss.t235 185.605
R10043 avss.n755 avss.n754 185
R10044 avss.n424 avss.n423 185
R10045 avss.n425 avss.n411 185
R10046 avss.n417 avss.n416 185
R10047 avss.n418 avss.n406 185
R10048 avss.t168 avss.n406 185
R10049 avss.n420 avss.n419 185
R10050 avss.n422 avss.n421 185
R10051 avss.n413 avss.n412 185
R10052 avss.n415 avss.n414 185
R10053 avss.n405 avss.n403 185
R10054 avss.n430 avss.n429 185
R10055 avss.n429 avss.t168 185
R10056 avss.n404 avss.n402 185
R10057 avss.n427 avss.n426 185
R10058 avss.n310 avss.n309 184.572
R10059 avss.n741 avss.t81 163.472
R10060 avss.t104 avss.t302 160.929
R10061 avss.t409 avss.t104 160.929
R10062 avss.t401 avss.t409 160.929
R10063 avss.t60 avss.t401 160.929
R10064 avss.t6 avss.t60 160.929
R10065 avss.t69 avss.t256 160.929
R10066 avss.t256 avss.t103 160.929
R10067 avss.t103 avss.t65 160.929
R10068 avss.t106 avss.t402 160.339
R10069 avss.t270 avss.t106 160.339
R10070 avss.t9 avss.t270 160.339
R10071 avss.t132 avss.t9 160.339
R10072 avss.t407 avss.t62 160.339
R10073 avss.t62 avss.t387 160.339
R10074 avss.t387 avss.t322 160.339
R10075 avss.t322 avss.t241 160.339
R10076 avss.t241 avss.t404 160.339
R10077 avss.t404 avss.t41 160.339
R10078 avss.t41 avss.t260 160.339
R10079 avss.t260 avss.t257 160.339
R10080 avss.t257 avss.t237 160.339
R10081 avss.t237 avss.t261 160.339
R10082 avss.n889 avss.n554 159.248
R10083 avss.n801 avss.n554 159.248
R10084 avss.n986 avss.n985 159.248
R10085 avss.n987 avss.n986 159.248
R10086 avss.n846 avss.n563 157.524
R10087 avss.n68 avss.t132 157.37
R10088 avss.n316 avss.t331 149.067
R10089 avss.n837 avss.t389 149.067
R10090 avss.n768 avss.t87 149.067
R10091 avss.n302 avss.t312 149.067
R10092 avss.n291 avss.t301 149.067
R10093 avss.n279 avss.t341 149.067
R10094 avss.n267 avss.t254 149.067
R10095 avss.n255 avss.t79 149.067
R10096 avss.n243 avss.t397 149.067
R10097 avss.n231 avss.t307 149.067
R10098 avss.n219 avss.t101 149.067
R10099 avss.n207 avss.t377 149.067
R10100 avss.n195 avss.t18 149.067
R10101 avss.n183 avss.t379 149.067
R10102 avss.n171 avss.t74 149.067
R10103 avss.n159 avss.t23 149.067
R10104 avss.n147 avss.t246 149.067
R10105 avss.n135 avss.t96 149.067
R10106 avss.n123 avss.t268 149.067
R10107 avss.n341 avss.t116 142.101
R10108 avss.n322 avss.t115 132.919
R10109 avss.n487 avss.n478 132.635
R10110 avss.n483 avss.n478 132.635
R10111 avss.n481 avss.n453 132.635
R10112 avss.n533 avss.n453 132.635
R10113 avss.n529 avss.n458 132.635
R10114 avss.n529 avss.n459 132.635
R10115 avss.n525 avss.n462 132.635
R10116 avss.n521 avss.n462 132.635
R10117 avss.n521 avss.n464 132.635
R10118 avss.n508 avss.n468 132.635
R10119 avss.n508 avss.n466 132.635
R10120 avss.n515 avss.n512 132.635
R10121 avss.n517 avss.n515 132.635
R10122 avss.n491 avss.n474 132.635
R10123 avss.n495 avss.n474 132.635
R10124 avss.n499 avss.n472 132.635
R10125 avss.n499 avss.n470 132.635
R10126 avss.n503 avss.n470 132.635
R10127 avss.n739 avss.t355 126.32
R10128 avss.n916 avss.t429 125.388
R10129 avss.n637 avss.t357 124.695
R10130 avss.n917 avss.t418 124.674
R10131 avss.n916 avss.t416 124.674
R10132 avss.n918 avss.t230 123.24
R10133 avss.n918 avss.t173 122.623
R10134 avss.t117 avss.n49 118.332
R10135 avss.t263 avss.t239 118.26
R10136 avss.t239 avss.t232 118.26
R10137 avss.t232 avss.t107 118.26
R10138 avss.t107 avss.t12 118.26
R10139 avss.t12 avss.t64 118.26
R10140 avss.n793 avss.n791 117.001
R10141 avss.n794 avss.n792 117.001
R10142 avss.n557 avss.n556 117.001
R10143 avss.n844 avss.n557 117.001
R10144 avss.n559 avss.n558 117.001
R10145 avss.n883 avss.n558 117.001
R10146 avss.n995 avss.n994 117.001
R10147 avss.n996 avss.n995 117.001
R10148 avss.n974 avss.n380 117.001
R10149 avss.n380 avss.n370 117.001
R10150 avss.n992 avss.n991 117.001
R10151 avss.n991 avss.n990 117.001
R10152 avss.n382 avss.n379 117.001
R10153 avss.n1100 avss.n1099 117.001
R10154 avss.t296 avss.n1100 117.001
R10155 avss.n1102 avss.n1101 117.001
R10156 avss.n1101 avss.t296 117.001
R10157 avss.n416 avss.n406 113.334
R10158 avss.n429 avss.n405 113.334
R10159 avss.n873 avss.n872 111.906
R10160 avss.t64 avss.t394 110.1
R10161 avss.t71 avss.n564 108.138
R10162 avss.t65 avss.n563 108.138
R10163 avss.t402 avss.n67 107.742
R10164 avss.n843 avss.t69 102.603
R10165 avss.n726 avss.n600 100.05
R10166 avss.n712 avss.n711 100.05
R10167 avss.n690 avss.n689 100.05
R10168 avss.n686 avss.n613 100.05
R10169 avss.n671 avss.n670 100.05
R10170 avss.n665 avss.n620 100.05
R10171 avss.n650 avss.n629 100.05
R10172 avss.n559 avss.n555 99.0123
R10173 avss.n992 avss.n367 99.0123
R10174 avss.n5 avss.n3 97.5005
R10175 avss.n7 avss.n5 97.5005
R10176 avss.n6 avss.n4 97.5005
R10177 avss.n1098 avss.n6 97.5005
R10178 avss.t68 avss.t14 96.6926
R10179 avss.n343 avss.t265 94.5922
R10180 avss.t318 avss.t259 91.065
R10181 avss.n782 avss.t40 88.2028
R10182 avss.n786 avss.t385 88.2028
R10183 avss.n930 avss.t110 88.2028
R10184 avss.n384 avss.t53 88.2028
R10185 avss.n388 avss.t274 88.2028
R10186 avss.n894 avss.t289 88.2028
R10187 avss.n932 avss.t175 87.8727
R10188 avss.n896 avss.t326 87.8727
R10189 avss.n411 avss.n409 87.6787
R10190 avss.n423 avss.n409 87.6787
R10191 avss.n931 avss.t112 87.5075
R10192 avss.n930 avss.t108 87.5075
R10193 avss.n895 avss.t287 87.5075
R10194 avss.n894 avss.t291 87.5075
R10195 avss.n1072 avss.n1071 86.2123
R10196 avss.n1069 avss.n22 86.2123
R10197 avss.n1086 avss.n1085 86.2123
R10198 avss.n1078 avss.n1077 86.2123
R10199 avss.n1104 avss.t297 85.1191
R10200 avss.t394 avss.n1096 84.4142
R10201 avss.n899 avss.t204 82.9912
R10202 avss.n540 avss.t195 82.9912
R10203 avss.n807 avss.t179 82.9912
R10204 avss.t172 avss.n818 82.9912
R10205 avss.t134 avss.n963 82.9912
R10206 avss.t177 avss.n960 82.9912
R10207 avss.n935 avss.t219 82.9912
R10208 avss.n922 avss.t155 82.9912
R10209 avss.n889 avss.n888 82.824
R10210 avss.n801 avss.n555 82.824
R10211 avss.n985 avss.n984 82.824
R10212 avss.n987 avss.n367 82.824
R10213 avss.t321 avss.t316 81.8562
R10214 avss.t168 avss.n407 77.7851
R10215 avss.t168 avss.n408 77.7851
R10216 avss.t313 avss.t238 76.3526
R10217 avss.t266 avss.t150 75.5042
R10218 avss.t94 avss.t93 75.5042
R10219 avss.t210 avss.t248 75.5042
R10220 avss.t247 avss.t216 75.5042
R10221 avss.t21 avss.t24 75.5042
R10222 avss.t206 avss.t75 75.5042
R10223 avss.t75 avss.t72 75.5042
R10224 avss.t212 avss.t380 75.5042
R10225 avss.t381 avss.t208 75.5042
R10226 avss.t16 avss.t19 75.5042
R10227 avss.t184 avss.t374 75.5042
R10228 avss.t375 avss.t159 75.5042
R10229 avss.t99 avss.t102 75.5042
R10230 avss.t139 avss.t309 75.5042
R10231 avss.t308 avss.t152 75.5042
R10232 avss.t152 avss.t395 75.5042
R10233 avss.t398 avss.t161 75.5042
R10234 avss.t77 avss.t76 75.5042
R10235 avss.t143 avss.t252 75.5042
R10236 avss.t255 avss.t197 75.5042
R10237 avss.t157 avss.t299 75.5042
R10238 avss.t298 avss.t188 75.5042
R10239 avss.t314 avss.t313 75.5042
R10240 avss.t113 avss.t398 73.8075
R10241 avss.n1097 avss.t235 73.162
R10242 avss.t63 avss.t212 72.9591
R10243 avss.n1097 avss.t263 71.6444
R10244 avss.n784 avss.n783 70.9775
R10245 avss.n782 avss.n781 70.9775
R10246 avss.n788 avss.n787 70.9775
R10247 avss.n786 avss.n785 70.9775
R10248 avss.n386 avss.n385 70.9775
R10249 avss.n384 avss.n383 70.9775
R10250 avss.n390 avss.n389 70.9775
R10251 avss.n388 avss.n387 70.9775
R10252 avss.n546 avss.n545 70.9612
R10253 avss.n544 avss.n543 70.9612
R10254 avss.n550 avss.n549 70.9612
R10255 avss.n823 avss.n822 70.9612
R10256 avss.n806 avss.n803 70.9612
R10257 avss.n820 avss.n819 70.9612
R10258 avss.n928 avss.n927 70.9612
R10259 avss.n926 avss.n925 70.9612
R10260 avss.n396 avss.n395 70.9612
R10261 avss.n394 avss.n393 70.9612
R10262 avss.n965 avss.n964 70.9612
R10263 avss.n962 avss.n961 70.9612
R10264 avss.t168 avss.n410 70.8113
R10265 avss.t168 avss.n428 70.8113
R10266 avss.t334 avss.t114 70.601
R10267 avss.n423 avss.n422 70.0005
R10268 avss.n427 avss.n411 70.0005
R10269 avss.t24 avss.t7 68.7174
R10270 avss.t130 avss.t131 67.9453
R10271 avss.t129 avss.t130 67.9453
R10272 avss.t128 avss.t129 67.9453
R10273 avss.t309 avss.t405 67.869
R10274 avss.t188 avss.t250 67.0206
R10275 avss.t2 avss.t77 64.4756
R10276 avss.t58 avss.t50 63.8987
R10277 avss.n885 avss.t286 63.7388
R10278 avss.t262 avss.t381 63.6272
R10279 avss.n378 avss.t48 63.1818
R10280 avss.n363 avss.n362 61.8334
R10281 avss.t8 avss.t303 61.3923
R10282 avss.n1089 avss.t136 61.1365
R10283 avss.n1095 avss.t4 60.3691
R10284 avss.n458 avss.n456 59.5655
R10285 avss.n491 avss.n490 59.5655
R10286 avss.n490 avss.n476 59.5655
R10287 avss.n456 avss.n454 59.5655
R10288 avss.t267 avss.n115 59.46
R10289 avss.t95 avss.n112 59.46
R10290 avss.t245 avss.n109 59.46
R10291 avss.t22 avss.n106 59.46
R10292 avss.t73 avss.n103 59.46
R10293 avss.t378 avss.n100 59.46
R10294 avss.t17 avss.n97 59.46
R10295 avss.t376 avss.n94 59.46
R10296 avss.t100 avss.n91 59.46
R10297 avss.t306 avss.n88 59.46
R10298 avss.t396 avss.n85 59.46
R10299 avss.t78 avss.n82 59.46
R10300 avss.t253 avss.n79 59.46
R10301 avss.t340 avss.n76 59.46
R10302 avss.t300 avss.n73 59.46
R10303 avss.t311 avss.n70 59.46
R10304 avss.t216 avss.t61 59.3854
R10305 avss.t102 avss.t1 58.5371
R10306 avss.n843 avss.t6 58.3266
R10307 avss.t299 avss.t251 57.6887
R10308 avss.n855 avss.t144 57.0602
R10309 avss.n979 avss.t271 56.675
R10310 avss.t243 avss.t143 55.1437
R10311 avss.t328 avss.t242 54.4857
R10312 avss.t386 avss.t16 54.2953
R10313 avss.t233 avss.t266 53.4469
R10314 avss.n800 avss.n554 53.1823
R10315 avss.n800 avss.n562 53.1823
R10316 avss.n828 avss.n552 53.1823
R10317 avss.n829 avss.n828 53.1823
R10318 avss.n373 avss.n371 53.1823
R10319 avss.n979 avss.n371 53.1823
R10320 avss.n986 avss.n372 53.1823
R10321 avss.n979 avss.n372 53.1823
R10322 avss.n18 avss.t70 52.9509
R10323 avss.n46 avss.t221 51.9277
R10324 avss.t248 avss.t66 50.0535
R10325 avss.n834 avss.n833 49.8123
R10326 avss.n797 avss.n796 49.8123
R10327 avss.n973 avss.n971 49.8123
R10328 avss.n975 avss.n381 49.8123
R10329 avss.t159 avss.t269 49.2052
R10330 avss.t168 avss.n409 48.6621
R10331 avss.t338 avss.t275 48.3568
R10332 avss.n884 avss.t288 47.2902
R10333 avss.t42 avss.t255 45.8117
R10334 avss.t324 avss.t336 45.5327
R10335 avss.t186 avss.t337 45.5327
R10336 avss.t141 avss.t305 45.5327
R10337 avss.n11 avss.n9 45.0005
R10338 avss.t221 avss.n9 45.0005
R10339 avss.n1092 avss.n10 45.0005
R10340 avss.t221 avss.n10 45.0005
R10341 avss.t13 avss.t184 44.9634
R10342 avss.n980 avss.t46 44.1554
R10343 avss.n978 avss.t273 44.1554
R10344 avss.t244 avss.t94 44.115
R10345 avss.t264 avss.n18 43.7421
R10346 avss.n343 avss.t261 43.6909
R10347 avss.t339 avss.n342 43.6909
R10348 avss.n419 avss.n410 43.3803
R10349 avss.n428 avss.n404 43.3803
R10350 avss.n422 avss.n410 43.3803
R10351 avss.n428 avss.n427 43.3803
R10352 avss.t131 avss.n49 42.7523
R10353 avss.n1075 avss.n1074 42.7189
R10354 avss.n990 avss.n370 42.3223
R10355 avss.t276 avss.t328 42.2073
R10356 avss.n642 avss.n633 40.8713
R10357 avss.n645 avss.n643 40.8713
R10358 avss.n657 avss.n656 40.8713
R10359 avss.n677 avss.n676 40.8713
R10360 avss.n679 avss.n678 40.8713
R10361 avss.n704 avss.n703 40.8713
R10362 avss.n718 avss.n717 40.8713
R10363 avss.n734 avss.n732 40.8713
R10364 avss.n748 avss.n746 40.8713
R10365 avss.n774 avss.n578 40.8713
R10366 avss.n842 avss.n565 40.8713
R10367 avss.t93 avss.t258 40.7216
R10368 avss.t374 avss.t97 39.8732
R10369 avss.n990 avss.t273 39.7462
R10370 avss.n644 avss.t364 39.5941
R10371 avss.t358 avss.n702 39.5941
R10372 avss.n761 avss.t15 39.5941
R10373 avss.n763 avss.t234 39.5941
R10374 avss.t197 avss.t236 39.0249
R10375 avss.n1010 avss.n1009 38.6099
R10376 avss.n1010 avss.n53 38.6076
R10377 avss.n1009 avss.n1008 38.5956
R10378 avss.t80 avss.n745 37.8912
R10379 avss.t388 avss.n774 37.8912
R10380 avss.n697 avss.t342 37.0397
R10381 avss.t354 avss.n733 37.0397
R10382 avss.n745 avss.t3 37.0397
R10383 avss.t302 avss.n842 37.0397
R10384 avss.t236 avss.t339 36.4798
R10385 avss.t14 avss.n1095 36.324
R10386 avss.n318 avss.n311 36.1417
R10387 avss.n312 avss.n311 36.1417
R10388 avss.n640 avss.n635 36.1417
R10389 avss.n640 avss.n631 36.1417
R10390 avss.n647 avss.n631 36.1417
R10391 avss.n647 avss.n627 36.1417
R10392 avss.n654 avss.n627 36.1417
R10393 avss.n654 avss.n622 36.1417
R10394 avss.n662 avss.n622 36.1417
R10395 avss.n662 avss.n623 36.1417
R10396 avss.n623 avss.n618 36.1417
R10397 avss.n674 avss.n618 36.1417
R10398 avss.n674 avss.n615 36.1417
R10399 avss.n681 avss.n615 36.1417
R10400 avss.n681 avss.n611 36.1417
R10401 avss.n695 avss.n611 36.1417
R10402 avss.n695 avss.n694 36.1417
R10403 avss.n694 avss.n609 36.1417
R10404 avss.n609 avss.n607 36.1417
R10405 avss.n706 avss.n607 36.1417
R10406 avss.n706 avss.n605 36.1417
R10407 avss.n715 avss.n605 36.1417
R10408 avss.n715 avss.n602 36.1417
R10409 avss.n722 avss.n602 36.1417
R10410 avss.n722 avss.n598 36.1417
R10411 avss.n729 avss.n598 36.1417
R10412 avss.n729 avss.n595 36.1417
R10413 avss.n736 avss.n595 36.1417
R10414 avss.n736 avss.n592 36.1417
R10415 avss.n743 avss.n592 36.1417
R10416 avss.n743 avss.n589 36.1417
R10417 avss.n750 avss.n589 36.1417
R10418 avss.n750 avss.n586 36.1417
R10419 avss.n759 avss.n586 36.1417
R10420 avss.n759 avss.n583 36.1417
R10421 avss.n765 avss.n583 36.1417
R10422 avss.n765 avss.n580 36.1417
R10423 avss.n772 avss.n580 36.1417
R10424 avss.n772 avss.n567 36.1417
R10425 avss.n840 avss.n567 36.1417
R10426 avss.n299 avss.n72 36.1417
R10427 avss.n305 avss.n72 36.1417
R10428 avss.n287 avss.n75 36.1417
R10429 avss.n294 avss.n75 36.1417
R10430 avss.n275 avss.n78 36.1417
R10431 avss.n282 avss.n78 36.1417
R10432 avss.n263 avss.n81 36.1417
R10433 avss.n270 avss.n81 36.1417
R10434 avss.n251 avss.n84 36.1417
R10435 avss.n258 avss.n84 36.1417
R10436 avss.n239 avss.n87 36.1417
R10437 avss.n246 avss.n87 36.1417
R10438 avss.n227 avss.n90 36.1417
R10439 avss.n234 avss.n90 36.1417
R10440 avss.n215 avss.n93 36.1417
R10441 avss.n222 avss.n93 36.1417
R10442 avss.n203 avss.n96 36.1417
R10443 avss.n210 avss.n96 36.1417
R10444 avss.n191 avss.n99 36.1417
R10445 avss.n198 avss.n99 36.1417
R10446 avss.n179 avss.n102 36.1417
R10447 avss.n186 avss.n102 36.1417
R10448 avss.n167 avss.n105 36.1417
R10449 avss.n174 avss.n105 36.1417
R10450 avss.n155 avss.n108 36.1417
R10451 avss.n162 avss.n108 36.1417
R10452 avss.n143 avss.n111 36.1417
R10453 avss.n150 avss.n111 36.1417
R10454 avss.n131 avss.n114 36.1417
R10455 avss.n138 avss.n114 36.1417
R10456 avss.n120 avss.n119 36.1417
R10457 avss.n126 avss.n120 36.1417
R10458 avss.n338 avss.n62 36.1417
R10459 avss.n1007 avss.n53 35.7393
R10460 avss.t97 avss.t375 35.6315
R10461 avss.n420 avss.n418 35.5561
R10462 avss.n415 avss.n412 35.5561
R10463 avss.n487 avss.n476 35.1094
R10464 avss.n533 avss.n454 35.1094
R10465 avss.t258 avss.t210 34.7831
R10466 avss.n658 avss.t370 34.4853
R10467 avss.n720 avss.t362 34.4853
R10468 avss.n731 avss.t98 34.4853
R10469 avss.n340 avss.n339 34.4123
R10470 avss.n341 avss.n340 34.4123
R10471 avss.n345 avss.n344 34.4123
R10472 avss.n344 avss.n343 34.4123
R10473 avss.n762 avss.t84 33.6338
R10474 avss.n1017 avss.t277 33.2544
R10475 avss.t86 avss.n762 32.7823
R10476 avss.n861 avss.n22 32.5005
R10477 avss.t128 avss.n861 32.5005
R10478 avss.n859 avss.n847 32.5005
R10479 avss.n847 avss.t67 32.5005
R10480 avss.n860 avss.n848 32.5005
R10481 avss.n848 avss.t67 32.5005
R10482 avss.n1094 avss.n1093 32.5005
R10483 avss.n1095 avss.n1094 32.5005
R10484 avss.n1091 avss.n1090 32.5005
R10485 avss.n1090 avss.n1089 32.5005
R10486 avss.n1087 avss.n1086 32.5005
R10487 avss.n1088 avss.n1087 32.5005
R10488 avss.n1077 avss.n1076 32.5005
R10489 avss.n1076 avss.n1075 32.5005
R10490 avss.n1073 avss.n1072 32.5005
R10491 avss.n1074 avss.n1073 32.5005
R10492 avss.t368 avss.n658 31.9308
R10493 avss.n720 avss.t350 31.9308
R10494 avss.n342 avss.t338 31.8139
R10495 avss.n1075 avss.t8 31.4638
R10496 avss.t150 avss.t244 31.3897
R10497 avss.t19 avss.t13 30.5413
R10498 avss.t252 avss.t42 29.693
R10499 avss.n494 avss.n471 29.6559
R10500 avss.n511 avss.n510 29.6559
R10501 avss.n527 avss.n526 29.6559
R10502 avss.n416 avss.n407 29.4328
R10503 avss.n413 avss.n408 29.4328
R10504 avss.n414 avss.n407 29.4328
R10505 avss.n408 avss.n405 29.4328
R10506 avss.t356 avss.n642 29.3764
R10507 avss.t352 avss.n697 29.3764
R10508 avss.n699 avss.t10 29.3764
R10509 avss.n888 avss.n887 28.9887
R10510 avss.n984 avss.n366 28.9887
R10511 avss.t43 avss.t186 28.9058
R10512 avss.t214 avss.t117 28.65
R10513 avss.t275 avss.t157 27.1479
R10514 avss.n860 avss.n850 27.1064
R10515 avss.n859 avss.n849 27.1064
R10516 avss.n538 avss.n537 26.8634
R10517 avss.t0 avss.t146 26.5545
R10518 avss.n1035 avss.t189 26.4633
R10519 avss.n1030 avss.t162 26.4633
R10520 avss.n41 avss.t180 26.4633
R10521 avss.n1025 avss.t198 26.4633
R10522 avss.n1044 avss.t225 26.4633
R10523 avss.n1050 avss.t135 26.4633
R10524 avss.n1060 avss.t222 26.4633
R10525 avss.n1055 avss.t228 26.4633
R10526 avss.n28 avss.t145 26.4633
R10527 avss.n36 avss.t166 26.4633
R10528 avss.t269 avss.t99 26.2995
R10529 avss.t259 avss.t334 26.092
R10530 avss.t66 avss.t247 25.4512
R10531 avss.n856 avss.t164 25.2191
R10532 avss.n853 avss.t200 25.2191
R10533 avss.t366 avss.n657 24.2676
R10534 avss.t310 avss.n659 24.2676
R10535 avss.t221 avss.t276 23.7898
R10536 avss.n16 avss.t333 23.7186
R10537 avss.n1080 avss.t304 23.4728
R10538 avss.n1083 avss.t335 23.4728
R10539 avss.n16 avss.t329 23.4728
R10540 avss.t323 avss.t214 23.2782
R10541 avss.n748 avss.t82 22.5646
R10542 avss.n1074 avss.t277 22.5108
R10543 avss.n887 avss.n886 22.5005
R10544 avss.n886 avss.n885 22.5005
R10545 avss.n561 avss.n560 22.5005
R10546 avss.n885 avss.n561 22.5005
R10547 avss.n366 avss.n364 22.5005
R10548 avss.n377 avss.n364 22.5005
R10549 avss.n993 avss.n365 22.5005
R10550 avss.n377 avss.n365 22.5005
R10551 avss.n1088 avss.t114 22.255
R10552 avss.t337 avss.t323 22.255
R10553 avss.n981 avss.t58 22.0815
R10554 avss.t265 avss.t233 22.0578
R10555 avss.t406 avss.n644 21.7131
R10556 avss.n679 avss.t348 21.7131
R10557 avss.n732 avss.t344 21.7131
R10558 avss.n779 avss.n570 21.3347
R10559 avss.n754 avss.t83 21.2805
R10560 avss.n754 avss.t85 21.2805
R10561 avss.n600 avss.t363 21.2805
R10562 avss.n600 avss.t345 21.2805
R10563 avss.n711 avss.t361 21.2805
R10564 avss.n711 avss.t351 21.2805
R10565 avss.n689 avss.t347 21.2805
R10566 avss.n689 avss.t359 21.2805
R10567 avss.n613 avss.t343 21.2805
R10568 avss.n613 avss.t353 21.2805
R10569 avss.n670 avss.t371 21.2805
R10570 avss.n670 avss.t349 21.2805
R10571 avss.n620 avss.t367 21.2805
R10572 avss.n620 avss.t369 21.2805
R10573 avss.n629 avss.t373 21.2805
R10574 avss.n629 avss.t365 21.2805
R10575 avss.t208 avss.t386 21.2094
R10576 avss.n575 avss.n570 21.1018
R10577 avss.n575 avss.n569 20.9741
R10578 avss.n833 avss.n832 20.8934
R10579 avss.n832 avss.n831 20.8934
R10580 avss.n798 avss.n797 20.8934
R10581 avss.n799 avss.n798 20.8934
R10582 avss.n973 avss.n972 20.8934
R10583 avss.n972 avss.n376 20.8934
R10584 avss.n976 avss.n975 20.8934
R10585 avss.n977 avss.n976 20.8934
R10586 avss.t303 avss.t120 20.7202
R10587 avss.t346 avss.n8 20.4359
R10588 avss.n1034 avss.n1033 20.3733
R10589 avss.n1032 avss.n1031 20.3733
R10590 avss.n1022 avss.n1021 20.3733
R10591 avss.n1024 avss.n1023 20.3733
R10592 avss.n1047 avss.n1046 20.3733
R10593 avss.n1049 avss.n1048 20.3733
R10594 avss.n1059 avss.n1058 20.3733
R10595 avss.n1057 avss.n1056 20.3733
R10596 avss.n33 avss.n32 20.3733
R10597 avss.n35 avss.n34 20.3733
R10598 avss.t76 avss.t243 20.361
R10599 avss avss.n424 20.2672
R10600 avss.n14 avss.n12 20.1729
R10601 avss.n18 avss.n12 20.1729
R10602 avss.n15 avss.n13 20.1729
R10603 avss.n18 avss.n13 20.1729
R10604 avss.n1082 avss.n1081 20.1668
R10605 avss.t50 avss.n980 19.7448
R10606 avss.t271 avss.n978 19.7448
R10607 avss.n349 avss.t403 19.4214
R10608 avss.n633 avss.t71 19.1587
R10609 avss.t344 avss.n731 19.1587
R10610 avss.t82 avss.n747 18.3072
R10611 avss.t238 avss.n341 18.2402
R10612 avss.n1035 avss.t191 18.0193
R10613 avss.t163 avss.n1030 18.0193
R10614 avss.n41 avss.t182 18.0193
R10615 avss.n1025 avss.t199 18.0193
R10616 avss.n1044 avss.t227 18.0193
R10617 avss.n1050 avss.t137 18.0193
R10618 avss.n1060 avss.t224 18.0193
R10619 avss.t229 avss.n1055 18.0193
R10620 avss.n28 avss.t148 18.0193
R10621 avss.n36 avss.t167 18.0193
R10622 avss.n517 avss.n516 17.9618
R10623 avss.n504 avss.n468 17.9618
R10624 avss.n504 avss.n503 17.9618
R10625 avss.n516 avss.n464 17.9618
R10626 avss.n431 avss.n430 17.9561
R10627 avss.t251 avss.t298 17.816
R10628 avss.n574 avss.n571 17.6946
R10629 avss.n431 avss.n402 17.6005
R10630 avss.n856 avss.t165 17.2863
R10631 avss.n853 avss.t201 17.2863
R10632 avss.t1 avss.t139 16.9676
R10633 avss.n484 avss 16.7292
R10634 avss.t336 avss.t43 16.6274
R10635 avss.n660 avss.t366 16.6043
R10636 avss.n660 avss.t310 16.6043
R10637 avss.n717 avss.t360 16.6043
R10638 avss.n783 avss.t36 16.5305
R10639 avss.n783 avss.t28 16.5305
R10640 avss.n781 avss.t30 16.5305
R10641 avss.n781 avss.t34 16.5305
R10642 avss.n787 avss.t32 16.5305
R10643 avss.n787 avss.t38 16.5305
R10644 avss.n785 avss.t26 16.5305
R10645 avss.n785 avss.t383 16.5305
R10646 avss.n545 avss.t285 16.5305
R10647 avss.n545 avss.t203 16.5305
R10648 avss.n543 avss.t294 16.5305
R10649 avss.n543 avss.t194 16.5305
R10650 avss.n549 avss.t281 16.5305
R10651 avss.n549 avss.t279 16.5305
R10652 avss.n822 avss.t292 16.5305
R10653 avss.n822 avss.t295 16.5305
R10654 avss.t179 avss.n806 16.5305
R10655 avss.n806 avss.t283 16.5305
R10656 avss.n819 avss.t172 16.5305
R10657 avss.n819 avss.t293 16.5305
R10658 avss.n385 avss.t55 16.5305
R10659 avss.n385 avss.t49 16.5305
R10660 avss.n383 avss.t45 16.5305
R10661 avss.n383 avss.t57 16.5305
R10662 avss.n389 avss.t59 16.5305
R10663 avss.n389 avss.t51 16.5305
R10664 avss.n387 avss.t47 16.5305
R10665 avss.n387 avss.t272 16.5305
R10666 avss.n927 avss.t90 16.5305
R10667 avss.n927 avss.t218 16.5305
R10668 avss.n925 avss.t392 16.5305
R10669 avss.n925 avss.t154 16.5305
R10670 avss.n395 avss.t89 16.5305
R10671 avss.n395 avss.t92 16.5305
R10672 avss.n393 avss.t391 16.5305
R10673 avss.n393 avss.t390 16.5305
R10674 avss.n964 avss.t134 16.5305
R10675 avss.n964 avss.t91 16.5305
R10676 avss.n961 avss.t177 16.5305
R10677 avss.n961 avss.t393 16.5305
R10678 avss.t61 avss.t21 16.1193
R10679 avss.n757 avss.n756 16.0275
R10680 avss.n780 avss.n569 15.8429
R10681 avss.t408 avss.t360 15.3271
R10682 avss.n425 avss 15.2894
R10683 avss.n755 avss.n753 15.2801
R10684 avss.n1071 avss.n17 14.9605
R10685 avss.n1085 avss.n1084 14.9605
R10686 avss.n1079 avss.n1078 14.9605
R10687 avss.n1069 avss.n1068 14.9605
R10688 avss.t316 avss.t264 14.8368
R10689 avss.t120 avss.t321 14.581
R10690 avss.n899 avss.t202 14.0925
R10691 avss.n540 avss.t192 14.0925
R10692 avss.n807 avss.t178 14.0925
R10693 avss.n818 avss.t170 14.0925
R10694 avss.n963 avss.t133 14.0925
R10695 avss.n960 avss.t176 14.0925
R10696 avss.n935 avss.t217 14.0925
R10697 avss.n922 avss.t153 14.0925
R10698 avss.n46 avss.t332 14.0694
R10699 avss.n645 avss.t372 14.0498
R10700 avss.t315 avss.n677 14.0498
R10701 avss.n699 avss.t346 14.0498
R10702 avss.t117 avss.n1014 13.0463
R10703 avss.n479 avss 12.9272
R10704 avss.n1089 avss.t242 12.7905
R10705 avss.n21 avss.n19 12.7179
R10706 avss.t130 avss.n19 12.7179
R10707 avss.n1070 avss.n20 12.7179
R10708 avss.t130 avss.n20 12.7179
R10709 avss.t111 avss.n376 12.513
R10710 avss.n1096 avss.t68 12.2789
R10711 avss.n358 avss.n355 12.189
R10712 avss.n421 avss.n420 12.0894
R10713 avss.n418 avss.n417 12.0894
R10714 avss.n426 avss.n402 12.0894
R10715 avss.n430 avss.n403 12.0894
R10716 avss.n867 avss.t400 11.9874
R10717 avss.t380 avss.t262 11.8775
R10718 avss.n1104 avss.n1103 11.8447
R10719 avss.n362 avss.t146 11.7601
R10720 avss.n643 avss.t356 11.4954
R10721 avss.n698 avss.t352 11.4954
R10722 avss.t10 avss.n698 11.4954
R10723 avss.n377 avss.t111 11.409
R10724 avss.t161 avss.t2 11.0291
R10725 avss.n368 avss.n49 10.9999
R10726 avss.n981 avss.n376 10.673
R10727 avss.n392 avss.n381 10.3632
R10728 avss.n971 avss.n970 10.3105
R10729 avss.n835 avss.n834 10.3105
R10730 avss.n796 avss.n795 10.3105
R10731 avss.n1038 avss.n1020 9.42076
R10732 avss.n1028 avss.n1020 9.42076
R10733 avss.n636 avss.n635 9.36464
R10734 avss.n352 avss.n57 9.35869
R10735 avss.n351 avss.n58 9.35222
R10736 avss.n350 avss.n59 9.34791
R10737 avss.n353 avss.n56 9.33929
R10738 avss.n354 avss.n55 9.33929
R10739 avss.n317 avss.n316 9.30641
R10740 avss.n316 avss.n315 9.3005
R10741 avss.n318 avss.n317 9.3005
R10742 avss.n314 avss.n311 9.3005
R10743 avss.n313 avss.n312 9.3005
R10744 avss.n638 avss.n637 9.3005
R10745 avss.n637 avss.n636 9.3005
R10746 avss.n650 avss.n649 9.3005
R10747 avss.n666 avss.n665 9.3005
R10748 avss.n665 avss.n664 9.3005
R10749 avss.n665 avss.n621 9.3005
R10750 avss.n671 avss.n614 9.3005
R10751 avss.n672 avss.n671 9.3005
R10752 avss.n671 avss.n668 9.3005
R10753 avss.n687 avss.n686 9.3005
R10754 avss.n686 avss.n685 9.3005
R10755 avss.n686 avss.n684 9.3005
R10756 avss.n691 avss.n690 9.3005
R10757 avss.n712 avss.n601 9.3005
R10758 avss.n713 avss.n712 9.3005
R10759 avss.n712 avss.n709 9.3005
R10760 avss.n727 avss.n726 9.3005
R10761 avss.n726 avss.n599 9.3005
R10762 avss.n726 avss.n725 9.3005
R10763 avss.n756 avss.n587 9.3005
R10764 avss.n769 avss.n768 9.3005
R10765 avss.n768 avss.n767 9.3005
R10766 avss.n838 avss.n837 9.3005
R10767 avss.n837 avss.n568 9.3005
R10768 avss.n740 avss.n739 9.3005
R10769 avss.n739 avss.n738 9.3005
R10770 avss.n640 avss.n639 9.3005
R10771 avss.n631 avss.n630 9.3005
R10772 avss.n648 avss.n647 9.3005
R10773 avss.n628 avss.n627 9.3005
R10774 avss.n654 avss.n653 9.3005
R10775 avss.n652 avss.n622 9.3005
R10776 avss.n663 avss.n662 9.3005
R10777 avss.n623 avss.n619 9.3005
R10778 avss.n667 avss.n618 9.3005
R10779 avss.n674 avss.n673 9.3005
R10780 avss.n669 avss.n615 9.3005
R10781 avss.n682 avss.n681 9.3005
R10782 avss.n683 avss.n611 9.3005
R10783 avss.n695 avss.n612 9.3005
R10784 avss.n694 avss.n693 9.3005
R10785 avss.n692 avss.n609 9.3005
R10786 avss.n688 avss.n607 9.3005
R10787 avss.n707 avss.n706 9.3005
R10788 avss.n708 avss.n605 9.3005
R10789 avss.n715 avss.n714 9.3005
R10790 avss.n710 avss.n602 9.3005
R10791 avss.n723 avss.n722 9.3005
R10792 avss.n724 avss.n598 9.3005
R10793 avss.n729 avss.n728 9.3005
R10794 avss.n595 avss.n594 9.3005
R10795 avss.n737 avss.n736 9.3005
R10796 avss.n593 avss.n592 9.3005
R10797 avss.n743 avss.n742 9.3005
R10798 avss.n589 avss.n588 9.3005
R10799 avss.n751 avss.n750 9.3005
R10800 avss.n752 avss.n586 9.3005
R10801 avss.n759 avss.n758 9.3005
R10802 avss.n583 avss.n582 9.3005
R10803 avss.n766 avss.n765 9.3005
R10804 avss.n581 avss.n580 9.3005
R10805 avss.n772 avss.n771 9.3005
R10806 avss.n770 avss.n567 9.3005
R10807 avss.n840 avss.n839 9.3005
R10808 avss.n877 avss.n850 9.3005
R10809 avss.n851 avss.n849 9.3005
R10810 avss.n865 avss.n864 9.3005
R10811 avss.n1002 avss.n357 9.3005
R10812 avss.n124 avss.n123 9.3005
R10813 avss.n123 avss.n122 9.3005
R10814 avss.n136 avss.n135 9.3005
R10815 avss.n135 avss.n134 9.3005
R10816 avss.n148 avss.n147 9.3005
R10817 avss.n147 avss.n146 9.3005
R10818 avss.n160 avss.n159 9.3005
R10819 avss.n159 avss.n158 9.3005
R10820 avss.n172 avss.n171 9.3005
R10821 avss.n171 avss.n170 9.3005
R10822 avss.n184 avss.n183 9.3005
R10823 avss.n183 avss.n182 9.3005
R10824 avss.n196 avss.n195 9.3005
R10825 avss.n195 avss.n194 9.3005
R10826 avss.n208 avss.n207 9.3005
R10827 avss.n207 avss.n206 9.3005
R10828 avss.n220 avss.n219 9.3005
R10829 avss.n219 avss.n218 9.3005
R10830 avss.n232 avss.n231 9.3005
R10831 avss.n231 avss.n230 9.3005
R10832 avss.n244 avss.n243 9.3005
R10833 avss.n243 avss.n242 9.3005
R10834 avss.n256 avss.n255 9.3005
R10835 avss.n255 avss.n254 9.3005
R10836 avss.n268 avss.n267 9.3005
R10837 avss.n267 avss.n266 9.3005
R10838 avss.n280 avss.n279 9.3005
R10839 avss.n279 avss.n278 9.3005
R10840 avss.n292 avss.n291 9.3005
R10841 avss.n291 avss.n290 9.3005
R10842 avss.n302 avss.n0 9.3005
R10843 avss.n303 avss.n302 9.3005
R10844 avss.n132 avss.n131 9.3005
R10845 avss.n133 avss.n114 9.3005
R10846 avss.n138 avss.n137 9.3005
R10847 avss.n144 avss.n143 9.3005
R10848 avss.n145 avss.n111 9.3005
R10849 avss.n150 avss.n149 9.3005
R10850 avss.n156 avss.n155 9.3005
R10851 avss.n157 avss.n108 9.3005
R10852 avss.n162 avss.n161 9.3005
R10853 avss.n168 avss.n167 9.3005
R10854 avss.n169 avss.n105 9.3005
R10855 avss.n174 avss.n173 9.3005
R10856 avss.n180 avss.n179 9.3005
R10857 avss.n181 avss.n102 9.3005
R10858 avss.n186 avss.n185 9.3005
R10859 avss.n192 avss.n191 9.3005
R10860 avss.n193 avss.n99 9.3005
R10861 avss.n198 avss.n197 9.3005
R10862 avss.n204 avss.n203 9.3005
R10863 avss.n205 avss.n96 9.3005
R10864 avss.n210 avss.n209 9.3005
R10865 avss.n216 avss.n215 9.3005
R10866 avss.n217 avss.n93 9.3005
R10867 avss.n222 avss.n221 9.3005
R10868 avss.n228 avss.n227 9.3005
R10869 avss.n229 avss.n90 9.3005
R10870 avss.n234 avss.n233 9.3005
R10871 avss.n240 avss.n239 9.3005
R10872 avss.n241 avss.n87 9.3005
R10873 avss.n246 avss.n245 9.3005
R10874 avss.n252 avss.n251 9.3005
R10875 avss.n253 avss.n84 9.3005
R10876 avss.n258 avss.n257 9.3005
R10877 avss.n264 avss.n263 9.3005
R10878 avss.n265 avss.n81 9.3005
R10879 avss.n270 avss.n269 9.3005
R10880 avss.n276 avss.n275 9.3005
R10881 avss.n277 avss.n78 9.3005
R10882 avss.n282 avss.n281 9.3005
R10883 avss.n288 avss.n287 9.3005
R10884 avss.n289 avss.n75 9.3005
R10885 avss.n294 avss.n293 9.3005
R10886 avss.n300 avss.n299 9.3005
R10887 avss.n301 avss.n72 9.3005
R10888 avss.n305 avss.n304 9.3005
R10889 avss.n119 avss.n60 9.3005
R10890 avss.n121 avss.n120 9.3005
R10891 avss.n126 avss.n125 9.3005
R10892 avss.n347 avss.n346 9.3005
R10893 avss.n1005 avss.n1004 9.20927
R10894 avss.n659 avss.t368 8.94099
R10895 avss.n703 avss.t408 8.94099
R10896 avss.t350 avss.n718 8.94099
R10897 avss.t48 avss.n377 8.83289
R10898 avss.t46 avss.n979 8.83289
R10899 avss.n868 avss.n866 8.81442
R10900 avss.n815 avss.t440 8.80038
R10901 avss.n814 avss.t428 8.80038
R10902 avss.n813 avss.t421 8.80038
R10903 avss.n812 avss.t444 8.80038
R10904 avss.n811 avss.t423 8.80038
R10905 avss.n810 avss.t410 8.80038
R10906 avss.n809 avss.t434 8.80038
R10907 avss.n539 avss.t426 8.80038
R10908 avss.n957 avss.t422 8.80038
R10909 avss.n956 avss.t425 8.80038
R10910 avss.n955 avss.t433 8.80038
R10911 avss.n954 avss.t413 8.80038
R10912 avss.n953 avss.t431 8.80038
R10913 avss.n952 avss.t443 8.80038
R10914 avss.n951 avss.t420 8.80038
R10915 avss.n950 avss.t427 8.80038
R10916 avss.n905 avss.t430 8.73382
R10917 avss.n906 avss.t417 8.73382
R10918 avss.n907 avss.t411 8.73382
R10919 avss.n908 avss.t436 8.73382
R10920 avss.n909 avss.t412 8.73382
R10921 avss.n910 avss.t437 8.73382
R10922 avss.n911 avss.t419 8.73382
R10923 avss.n912 avss.t415 8.73382
R10924 avss.n941 avss.t435 8.73382
R10925 avss.n942 avss.t438 8.73382
R10926 avss.n943 avss.t442 8.73382
R10927 avss.n944 avss.t424 8.73382
R10928 avss.n945 avss.t441 8.73382
R10929 avss.n946 avss.t414 8.73382
R10930 avss.n947 avss.t432 8.73382
R10931 avss.n948 avss.t439 8.73382
R10932 avss.n492 avss.n475 8.61832
R10933 avss.n493 avss.n492 8.61832
R10934 avss.n494 avss.n493 8.61832
R10935 avss.n500 avss.n471 8.61832
R10936 avss.n501 avss.n500 8.61832
R10937 avss.n502 avss.n501 8.61832
R10938 avss.n509 avss.n467 8.61832
R10939 avss.n510 avss.n509 8.61832
R10940 avss.n511 avss.n465 8.61832
R10941 avss.n518 avss.n465 8.61832
R10942 avss.n460 avss.n452 8.61832
R10943 avss.n528 avss.n460 8.61832
R10944 avss.n528 avss.n527 8.61832
R10945 avss.n526 avss.n461 8.61832
R10946 avss.n520 avss.n461 8.61832
R10947 avss.n520 avss.n519 8.61832
R10948 avss.n486 avss.n485 8.61832
R10949 avss.n485 avss.n484 8.61832
R10950 avss.n479 avss.n451 8.61832
R10951 avss.t250 avss.t314 8.48406
R10952 avss.n866 avss.n358 8.4666
R10953 avss.n877 avss.n876 8.37766
R10954 avss.n876 avss.n851 8.37766
R10955 avss.n38 avss.n30 8.11041
R10956 avss.n1064 avss.n30 8.11041
R10957 avss.n763 avss.t86 8.08952
R10958 avss.n1002 avss.n1001 8.02619
R10959 avss.n1001 avss.n358 8.00675
R10960 avss.n878 avss.n851 7.938
R10961 avss.n878 avss.n877 7.938
R10962 avss avss.n836 7.87749
R10963 avss.t405 avss.t308 7.63571
R10964 avss.n913 avss.n539 7.62598
R10965 avss.n950 avss.n949 7.62598
R10966 avss.n869 avss.n865 7.48375
R10967 avss.n424 avss.n421 7.46717
R10968 avss.n426 avss.n425 7.46717
R10969 avss.n417 avss.n415 7.46717
R10970 avss.n412 avss.n403 7.46717
R10971 avss.t84 avss.n761 7.23804
R10972 avss.n869 avss.n868 7.16066
R10973 avss.n920 avss.n919 7.079
R10974 avss.t332 avss.t4 6.90708
R10975 avss.n865 avss.n356 6.89147
R10976 avss.n1002 avss.n356 6.89083
R10977 avss.n48 avss.n45 6.88285
R10978 avss.n362 avss.n48 6.88285
R10979 avss.n47 avss.n44 6.88285
R10980 avss.n47 avss.n46 6.88285
R10981 avss.t7 avss.t206 6.78735
R10982 avss.n880 avss.n879 6.5005
R10983 avss.n881 avss.n880 6.5005
R10984 avss.n875 avss.n874 6.5005
R10985 avss.n874 avss.n873 6.5005
R10986 avss.n891 avss.n551 6.47706
R10987 avss.n891 avss.n547 6.47706
R10988 avss.n824 avss.n821 6.47706
R10989 avss.n824 avss.n542 6.47706
R10990 avss.n966 avss.n375 6.47706
R10991 avss.n929 avss.n375 6.47706
R10992 avss.n401 avss.n374 6.47706
R10993 avss.n924 avss.n374 6.47706
R10994 avss.n535 avss.n451 6.46387
R10995 avss.n676 avss.t370 6.38657
R10996 avss.n702 avss.n8 6.38657
R10997 avss.t362 avss.n719 6.38657
R10998 avss.n719 avss.t98 6.38657
R10999 avss.n1106 avss.n1105 6.05765
R11000 avss.n1016 avss.n1015 5.90959
R11001 avss.n1017 avss.n1016 5.90959
R11002 avss.n1019 avss.n1018 5.90959
R11003 avss.n1018 avss.n1017 5.90959
R11004 avss.n368 avss.t141 5.88388
R11005 avss.n1105 avss.n2 5.78505
R11006 avss.n867 avss.n858 5.7846
R11007 avss.n857 avss.n856 5.76099
R11008 avss.n854 avss.n853 5.76099
R11009 avss.n836 avss.n780 5.71512
R11010 avss.n1029 avss.n1028 5.70305
R11011 avss.n1027 avss.n1026 5.70305
R11012 avss.n1052 avss.n1051 5.70305
R11013 avss.n1054 avss.n1053 5.70305
R11014 avss.n38 avss.n37 5.70305
R11015 avss.n852 avss.n851 5.6605
R11016 avss.n1036 avss.n1035 5.6605
R11017 avss.n1030 avss.n1029 5.6605
R11018 avss.n1038 avss.n1037 5.6605
R11019 avss.n42 avss.n41 5.6605
R11020 avss.n1026 avss.n1025 5.6605
R11021 avss.n1040 avss.n1039 5.6605
R11022 avss.n1045 avss.n1044 5.6605
R11023 avss.n1051 avss.n1050 5.6605
R11024 avss.n1043 avss.n31 5.6605
R11025 avss.n1061 avss.n1060 5.6605
R11026 avss.n1055 avss.n1054 5.6605
R11027 avss.n1063 avss.n1062 5.6605
R11028 avss.n29 avss.n28 5.6605
R11029 avss.n37 avss.n36 5.6605
R11030 avss.n1065 avss.n1064 5.6605
R11031 avss.n877 avss.n858 5.6605
R11032 avss.t70 avss.t318 5.62808
R11033 avss.n780 avss.n779 5.46789
R11034 avss.n776 avss.n572 5.27077
R11035 avss.n776 avss.n775 5.27077
R11036 avss.n573 avss.n571 5.27077
R11037 avss.n775 avss.n573 5.27077
R11038 avss.n1000 avss.n999 5.27077
R11039 avss.n999 avss.n998 5.27077
R11040 avss.n871 avss.n870 5.27077
R11041 avss.n872 avss.n871 5.27077
R11042 avss.t372 avss.t406 5.10935
R11043 avss.t348 avss.t315 5.10935
R11044 avss.n544 avss.n542 5.07277
R11045 avss.n824 avss.n823 5.07277
R11046 avss.n821 avss.n820 5.07277
R11047 avss.n926 avss.n924 5.07277
R11048 avss.n394 avss.n374 5.07277
R11049 avss.n962 avss.n401 5.07277
R11050 avss.n778 avss.n777 5.0436
R11051 avss.n777 avss.n563 5.0436
R11052 avss.n577 avss.n576 5.0436
R11053 avss.n577 avss.n564 5.0436
R11054 avss.n361 avss.n359 5.0436
R11055 avss.t0 avss.n361 5.0436
R11056 avss.n863 avss.n360 5.0436
R11057 avss.t0 avss.n360 5.0436
R11058 avss.n1013 avss.n1012 5.0436
R11059 avss.n1014 avss.n1013 5.0436
R11060 avss.n66 avss.n54 5.0436
R11061 avss.n67 avss.n66 5.0436
R11062 avss.n447 avss.n446 5.0005
R11063 avss.n446 avss.n445 5.0005
R11064 avss.n438 avss.n434 5.0005
R11065 avss.n444 avss.n438 5.0005
R11066 avss.n442 avss.n441 5.0005
R11067 avss.n443 avss.n442 5.0005
R11068 avss.n440 avss.n437 5.0005
R11069 avss.n439 avss.n437 5.0005
R11070 avss.n547 avss.n546 4.95167
R11071 avss.n803 avss.n551 4.95167
R11072 avss.n929 avss.n928 4.95167
R11073 avss.n966 avss.n965 4.95167
R11074 avss.n1007 avss.n1006 4.86769
R11075 avss.n63 avss.n62 4.6805
R11076 avss.t159 avss.n63 4.6805
R11077 avss.n65 avss.n64 4.6805
R11078 avss.t159 avss.n65 4.6805
R11079 avss.n651 avss.n650 4.63624
R11080 avss.n690 avss.n606 4.63624
R11081 avss.n949 avss.n948 4.60905
R11082 avss.n913 avss.n912 4.60905
R11083 avss.n541 avss.n540 4.5005
R11084 avss.n900 avss.n899 4.5005
R11085 avss.n892 avss.n891 4.5005
R11086 avss.n902 avss.n901 4.5005
R11087 avss.n904 avss.n903 4.5005
R11088 avss.n818 avss.n817 4.5005
R11089 avss.n808 avss.n807 4.5005
R11090 avss.n816 avss.n802 4.5005
R11091 avss.n805 avss.n804 4.5005
R11092 avss.n397 avss.n375 4.5005
R11093 avss.n923 avss.n922 4.5005
R11094 avss.n936 avss.n935 4.5005
R11095 avss.n940 avss.n939 4.5005
R11096 avss.n938 avss.n937 4.5005
R11097 avss.n960 avss.n959 4.5005
R11098 avss.n963 avss.n399 4.5005
R11099 avss.n958 avss.n400 4.5005
R11100 avss.n968 avss.n967 4.5005
R11101 avss.n435 avss.n432 4.3603
R11102 avss.n449 avss.n433 4.34678
R11103 avss.n435 avss.n433 4.34003
R11104 avss.n852 avss.n26 4.00655
R11105 avss.n827 avss.n825 3.9532
R11106 avss.n827 avss.n826 3.9532
R11107 avss.n890 avss.n553 3.9532
R11108 avss.n826 avss.n553 3.9532
R11109 avss.n983 avss.n982 3.9532
R11110 avss.n982 avss.n981 3.9532
R11111 avss.n989 avss.n988 3.9532
R11112 avss.n990 avss.n989 3.9532
R11113 avss.n1105 avss.n1104 3.94537
R11114 avss.n915 avss.n914 3.9105
R11115 avss.n1014 avss.t305 3.83749
R11116 avss.n678 avss.t342 3.83214
R11117 avss.n734 avss.t354 3.83214
R11118 avss.n733 avss.t3 3.83214
R11119 avss.n450 avss.n449 3.78259
R11120 avss.n805 avss.n548 3.77378
R11121 avss.n969 avss.n968 3.77378
R11122 avss.n893 avss.n892 3.77209
R11123 avss.n398 avss.n397 3.77209
R11124 avss.n901 avss.n898 3.77014
R11125 avss.n937 avss.n934 3.77014
R11126 avss.n1068 avss.n1067 3.68964
R11127 avss.n1037 avss.n40 3.57087
R11128 avss.n1041 avss.n1040 3.57087
R11129 avss.n1043 avss.n1042 3.57087
R11130 avss.n1062 avss.n27 3.57087
R11131 avss.n1066 avss.n1065 3.57087
R11132 avss.n392 avss.n391 3.4105
R11133 avss.n933 avss.n932 3.4105
R11134 avss.n897 avss.n896 3.4105
R11135 avss.n790 avss.n789 3.4105
R11136 avss.n1033 avss.t122 3.3065
R11137 avss.n1033 avss.t190 3.3065
R11138 avss.n1031 avss.t163 3.3065
R11139 avss.n1031 avss.t121 3.3065
R11140 avss.n1021 avss.t126 3.3065
R11141 avss.n1021 avss.t181 3.3065
R11142 avss.t199 avss.n1024 3.3065
R11143 avss.n1024 avss.t123 3.3065
R11144 avss.n1046 avss.t118 3.3065
R11145 avss.n1046 avss.t226 3.3065
R11146 avss.t137 avss.n1049 3.3065
R11147 avss.n1049 avss.t399 3.3065
R11148 avss.n1058 avss.t124 3.3065
R11149 avss.n1058 avss.t223 3.3065
R11150 avss.n1056 avss.t229 3.3065
R11151 avss.n1056 avss.t127 3.3065
R11152 avss.n32 avss.t119 3.3065
R11153 avss.n32 avss.t147 3.3065
R11154 avss.t167 avss.n35 3.3065
R11155 avss.n35 avss.t125 3.3065
R11156 avss.n1081 avss.t319 3.3065
R11157 avss.n1081 avss.t317 3.3065
R11158 avss.t128 avss.n862 3.2875
R11159 avss.n804 avss.n551 3.23878
R11160 avss.n902 avss.n547 3.23878
R11161 avss.n821 avss.n802 3.23878
R11162 avss.n903 avss.n542 3.23878
R11163 avss.n967 avss.n966 3.23878
R11164 avss.n938 avss.n929 3.23878
R11165 avss.n401 avss.n400 3.23878
R11166 avss.n939 avss.n924 3.23878
R11167 avss.n949 avss.n921 3.22196
R11168 avss.n905 avss.n904 3.21858
R11169 avss.n941 avss.n940 3.21858
R11170 avss.n816 avss.n815 3.12292
R11171 avss.n958 avss.n957 3.12292
R11172 avss.n536 avss.n535 3.1005
R11173 avss.n746 avss.t80 2.98066
R11174 avss.n68 avss.t407 2.96975
R11175 avss.n1008 avss.n1007 2.83532
R11176 avss.n1103 avss.n3 2.6005
R11177 avss.n775 avss.n565 2.55493
R11178 avss.t72 avss.t63 2.54557
R11179 avss.n1064 avss.n1063 2.42291
R11180 avss.n1063 avss.n31 2.42291
R11181 avss.n1039 avss.n1038 2.42291
R11182 avss.n1028 avss.n1027 2.42291
R11183 avss.n1053 avss.n1052 2.42291
R11184 avss.n1053 avss.n38 2.42291
R11185 avss.n502 avss.n467 2.40842
R11186 avss.n519 avss.n518 2.40842
R11187 avss.n537 avss.n431 2.32925
R11188 avss.n1003 avss.n1002 2.31886
R11189 avss.n865 avss.n26 2.31886
R11190 avss.n486 avss.n475 2.28169
R11191 avss.n534 avss.n452 2.28169
R11192 avss.n440 avss.n436 2.25932
R11193 avss.n868 avss.n867 2.2505
R11194 avss.n915 avss.n355 2.221
R11195 avss.n536 avss.n450 2.17339
R11196 avss.n535 avss.n534 2.15496
R11197 avss avss.n918 2.13136
R11198 avss.n914 avss.n913 2.12151
R11199 avss.n804 avss.n802 2.11769
R11200 avss.n903 avss.n902 2.11769
R11201 avss.n967 avss.n400 2.11769
R11202 avss.n939 avss.n938 2.11769
R11203 avss.n1004 avss.n355 2.058
R11204 avss.n914 avss.n538 1.90581
R11205 avss.n897 avss.n538 1.80585
R11206 avss.n1039 avss.n43 1.80222
R11207 avss.n1027 avss.n39 1.80222
R11208 avss.t395 avss.t113 1.69721
R11209 avss.n352 avss.n351 1.6605
R11210 avss.n920 avss.n915 1.65831
R11211 avss.n969 avss.n398 1.58008
R11212 avss.n934 avss.n398 1.58008
R11213 avss.n898 avss.n893 1.58008
R11214 avss.n893 avss.n548 1.58008
R11215 avss.n1011 avss.n51 1.50436
R11216 avss.n342 avss.n51 1.50436
R11217 avss.n52 avss.n50 1.50436
R11218 avss.n342 avss.n50 1.50436
R11219 avss.n348 avss.n60 1.48467
R11220 avss.n919 avss 1.41066
R11221 avss.n330 avss.n1 1.34141
R11222 avss.n351 avss.n350 1.338
R11223 avss.n347 avss.n61 1.32209
R11224 avss.n1017 avss.t324 1.2795
R11225 avss.n656 avss.t364 1.27771
R11226 avss.n704 avss.t358 1.27771
R11227 avss.n747 avss.t15 1.27771
R11228 avss.t234 avss.n578 1.27771
R11229 avss.n354 avss.n353 1.27675
R11230 avss.t116 avss.n322 1.27303
R11231 avss.n862 avss.n363 1.27293
R11232 avss.n325 avss.n324 1.14936
R11233 avss.n335 avss.n334 1.14936
R11234 avss.n336 avss.n335 1.14839
R11235 avss.n324 avss.n323 1.14811
R11236 avss.n323 avss.n61 1.08686
R11237 avss.n326 avss.n325 1.08686
R11238 avss.n327 avss.n326 1.08686
R11239 avss.n329 avss.n328 1.08686
R11240 avss.n334 avss.n333 1.08686
R11241 avss.n333 avss.n332 1.08686
R11242 avss.n332 avss.n331 1.08686
R11243 avss.n331 avss.n330 1.08686
R11244 avss.n328 avss.n327 1.08005
R11245 avss.n1034 avss.n1032 1.05355
R11246 avss.n1023 avss.n1022 1.05355
R11247 avss.n1048 avss.n1047 1.05355
R11248 avss.n1059 avss.n1057 1.05355
R11249 avss.n34 avss.n33 1.05355
R11250 avss.n353 avss.n352 1.00987
R11251 avss.n337 avss.n336 1.00505
R11252 avss.n933 avss.n921 1.00226
R11253 avss.n857 avss.n855 0.955426
R11254 avss.n855 avss.n854 0.953203
R11255 avss.n1005 avss.n1 0.902375
R11256 avss.n349 avss.n348 0.839875
R11257 avss.n815 avss.n814 0.807835
R11258 avss.n814 avss.n813 0.807835
R11259 avss.n813 avss.n812 0.807835
R11260 avss.n812 avss.n811 0.807835
R11261 avss.n811 avss.n810 0.807835
R11262 avss.n810 avss.n809 0.807835
R11263 avss.n809 avss.n539 0.807835
R11264 avss.n957 avss.n956 0.807835
R11265 avss.n956 avss.n955 0.807835
R11266 avss.n955 avss.n954 0.807835
R11267 avss.n954 avss.n953 0.807835
R11268 avss.n953 avss.n952 0.807835
R11269 avss.n952 avss.n951 0.807835
R11270 avss.n951 avss.n950 0.807835
R11271 avss.n906 avss.n905 0.80776
R11272 avss.n907 avss.n906 0.80776
R11273 avss.n908 avss.n907 0.80776
R11274 avss.n909 avss.n908 0.80776
R11275 avss.n910 avss.n909 0.80776
R11276 avss.n911 avss.n910 0.80776
R11277 avss.n912 avss.n911 0.80776
R11278 avss.n942 avss.n941 0.80776
R11279 avss.n943 avss.n942 0.80776
R11280 avss.n944 avss.n943 0.80776
R11281 avss.n945 avss.n944 0.80776
R11282 avss.n946 avss.n945 0.80776
R11283 avss.n947 avss.n946 0.80776
R11284 avss.n948 avss.n947 0.80776
R11285 avss.n1107 avss.n1106 0.79175
R11286 avss.n448 avss.n434 0.753441
R11287 avss.n756 avss.n755 0.747945
R11288 avss.n788 avss.n786 0.695812
R11289 avss.n900 avss.n541 0.695812
R11290 avss.n546 avss.n544 0.695812
R11291 avss.n820 avss.n803 0.695812
R11292 avss.n817 avss.n808 0.695812
R11293 avss.n931 avss.n930 0.695812
R11294 avss.n390 avss.n388 0.695812
R11295 avss.n928 avss.n926 0.695812
R11296 avss.n396 avss.n394 0.695812
R11297 avss.n965 avss.n962 0.695812
R11298 avss.n936 avss.n923 0.695812
R11299 avss.n959 avss.n399 0.695812
R11300 avss.n895 avss.n894 0.695812
R11301 avss.t54 avss.n378 0.69443
R11302 avss.n917 avss.n916 0.693859
R11303 avss.n784 avss.n782 0.679185
R11304 avss.n386 avss.n384 0.679185
R11305 avss.n823 avss.n550 0.676856
R11306 avss.n789 avss.n788 0.654797
R11307 avss.n391 avss.n390 0.654797
R11308 avss.n1068 avss.n25 0.635318
R11309 avss.n921 avss.n920 0.622375
R11310 avss.n43 avss.n31 0.62119
R11311 avss.n1052 avss.n39 0.62119
R11312 avss.n904 avss.n541 0.572766
R11313 avss.n817 avss.n816 0.572766
R11314 avss.n940 avss.n923 0.572766
R11315 avss.n959 avss.n958 0.572766
R11316 avss.n450 avss.n432 0.571446
R11317 avss.n1032 avss.n1029 0.527027
R11318 avss.n1036 avss.n1034 0.527027
R11319 avss.n1026 avss.n1023 0.527027
R11320 avss.n1022 avss.n42 0.527027
R11321 avss.n1051 avss.n1048 0.527027
R11322 avss.n1047 avss.n1045 0.527027
R11323 avss.n1057 avss.n1054 0.527027
R11324 avss.n1061 avss.n1059 0.527027
R11325 avss.n37 avss.n34 0.527027
R11326 avss.n33 avss.n29 0.527027
R11327 avss.t136 avss.n1088 0.512098
R11328 avss.n1067 avss.n26 0.505881
R11329 avss.n1067 avss.n1066 0.497189
R11330 avss.n1066 avss.n27 0.478977
R11331 avss.n1042 avss.n27 0.478977
R11332 avss.n1042 avss.n1041 0.478977
R11333 avss.n1041 avss.n40 0.478977
R11334 avss.n901 avss.n900 0.451672
R11335 avss.n892 avss.n550 0.451672
R11336 avss.n808 avss.n805 0.451672
R11337 avss.n397 avss.n396 0.451672
R11338 avss.n937 avss.n936 0.451672
R11339 avss.n968 avss.n399 0.451672
R11340 avss.n775 avss.t388 0.426238
R11341 avss.n919 avss.n917 0.416516
R11342 avss.n1004 avss.n1003 0.387296
R11343 avss.n1003 avss.n40 0.380881
R11344 avss.n1106 avss.n1 0.364875
R11345 avss.n980 avss.t88 0.344476
R11346 avss.n932 avss.n931 0.311047
R11347 avss.n896 avss.n895 0.311047
R11348 avss.n1083 avss.n1082 0.291392
R11349 avss.n1082 avss.n1080 0.291392
R11350 avss.n436 avss.n435 0.274029
R11351 avss.n447 avss.n433 0.266214
R11352 avss.n449 avss.n448 0.266214
R11353 avss.n441 avss.n432 0.266214
R11354 avss.n132 avss 0.248811
R11355 avss.n144 avss 0.248811
R11356 avss.n156 avss 0.248811
R11357 avss.n168 avss 0.248811
R11358 avss.n180 avss 0.248811
R11359 avss.n192 avss 0.248811
R11360 avss.n204 avss 0.248811
R11361 avss.n216 avss 0.248811
R11362 avss.n228 avss 0.248811
R11363 avss.n240 avss 0.248811
R11364 avss.n252 avss 0.248811
R11365 avss.n264 avss 0.248811
R11366 avss.n276 avss 0.248811
R11367 avss.n288 avss 0.248811
R11368 avss.n300 avss 0.248811
R11369 avss.n934 avss.n933 0.237405
R11370 avss.n898 avss.n897 0.237405
R11371 avss.n23 avss.n17 0.182466
R11372 avss.n978 avss.t109 0.176117
R11373 avss.n350 avss.n349 0.153
R11374 avss.n348 avss.n347 0.128909
R11375 avss.n1084 avss.n16 0.119588
R11376 avss.n970 avss.n969 0.118318
R11377 avss.n795 avss.n548 0.118318
R11378 avss.n45 avss.n43 0.11675
R11379 avss.n44 avss.n39 0.11675
R11380 avss.n24 avss.n23 0.11673
R11381 avss.n970 avss.n392 0.114189
R11382 avss.n795 avss.n790 0.114189
R11383 avss.n25 avss.n24 0.113554
R11384 avss.n879 avss.n878 0.109912
R11385 avss.n876 avss.n875 0.109912
R11386 avss avss.n1107 0.107764
R11387 avss.n1006 avss.n1005 0.10175
R11388 avss.n1015 avss.n30 0.0994362
R11389 avss.n1020 avss.n1019 0.0994362
R11390 avss.n574 avss.n569 0.0907913
R11391 avss.n870 avss.n869 0.0890714
R11392 avss.n1001 avss.n1000 0.0890714
R11393 avss.n572 avss.n570 0.0890714
R11394 avss.n863 avss.n356 0.0866111
R11395 avss.n1009 avss.n54 0.0850455
R11396 avss.n1012 avss.n53 0.0850455
R11397 avss.n866 avss.n359 0.0850455
R11398 avss.n576 avss.n575 0.0850455
R11399 avss.n779 avss.n778 0.0850455
R11400 avss.n337 avss.n329 0.0823182
R11401 avss.n314 avss.n313 0.0815811
R11402 avss.n121 avss.n60 0.0815811
R11403 avss.n133 avss.n132 0.0815811
R11404 avss.n145 avss.n144 0.0815811
R11405 avss.n157 avss.n156 0.0815811
R11406 avss.n169 avss.n168 0.0815811
R11407 avss.n181 avss.n180 0.0815811
R11408 avss.n193 avss.n192 0.0815811
R11409 avss.n205 avss.n204 0.0815811
R11410 avss.n217 avss.n216 0.0815811
R11411 avss.n229 avss.n228 0.0815811
R11412 avss.n241 avss.n240 0.0815811
R11413 avss.n253 avss.n252 0.0815811
R11414 avss.n265 avss.n264 0.0815811
R11415 avss.n277 avss.n276 0.0815811
R11416 avss.n289 avss.n288 0.0815811
R11417 avss.n301 avss.n300 0.0815811
R11418 avss.n836 avss.n835 0.0798919
R11419 avss.n648 avss.n630 0.0794474
R11420 avss.n653 avss.n652 0.0794474
R11421 avss.n683 avss.n682 0.0794474
R11422 avss.n693 avss.n692 0.0794474
R11423 avss.n708 avss.n707 0.0794474
R11424 avss.n737 avss.n594 0.0794474
R11425 avss.n751 avss.n588 0.0794474
R11426 avss.n766 avss.n582 0.0794474
R11427 avss.n771 avss.n770 0.0794474
R11428 avss.n338 avss.n337 0.0793136
R11429 avss.n537 avss.n536 0.0784703
R11430 avss.n668 avss.n667 0.072046
R11431 avss.n725 avss.n723 0.072046
R11432 avss.n891 avss.n890 0.0674065
R11433 avss.n825 avss.n824 0.0674065
R11434 avss.n988 avss.n374 0.0674065
R11435 avss.n983 avss.n375 0.0674065
R11436 avss.n667 avss.n666 0.0671118
R11437 avss.n723 avss.n601 0.0671118
R11438 avss.n757 avss.n582 0.0638224
R11439 avss.n741 avss.n588 0.0621776
R11440 avss.n753 avss.n751 0.0555987
R11441 avss.n125 avss.n122 0.0553986
R11442 avss.n137 avss.n134 0.0553986
R11443 avss.n149 avss.n146 0.0553986
R11444 avss.n161 avss.n158 0.0553986
R11445 avss.n173 avss.n170 0.0553986
R11446 avss.n185 avss.n182 0.0553986
R11447 avss.n197 avss.n194 0.0553986
R11448 avss.n209 avss.n206 0.0553986
R11449 avss.n221 avss.n218 0.0553986
R11450 avss.n233 avss.n230 0.0553986
R11451 avss.n245 avss.n242 0.0553986
R11452 avss.n257 avss.n254 0.0553986
R11453 avss.n269 avss.n266 0.0553986
R11454 avss.n281 avss.n278 0.0553986
R11455 avss.n293 avss.n290 0.0553986
R11456 avss.n304 avss.n303 0.0553986
R11457 avss.n767 avss.n581 0.0539539
R11458 avss.n839 avss.n568 0.0539539
R11459 avss.n1079 avss.n17 0.0538514
R11460 avss.n835 avss.n790 0.0532162
R11461 avss.n652 avss.n621 0.0523092
R11462 avss.n673 avss.n672 0.0523092
R11463 avss.n687 avss.n612 0.0523092
R11464 avss.n709 avss.n708 0.0523092
R11465 avss.n724 avss.n599 0.0523092
R11466 avss.n738 avss.n593 0.0498421
R11467 avss.n649 avss.n628 0.047375
R11468 avss.n664 avss.n619 0.047375
R11469 avss.n682 avss.n614 0.047375
R11470 avss.n691 avss.n688 0.047375
R11471 avss.n713 avss.n710 0.047375
R11472 avss.n727 avss.n594 0.047375
R11473 avss.n1107 avss 0.04675
R11474 avss.n639 avss.n638 0.0449079
R11475 avss.n758 avss.n587 0.0440855
R11476 avss.n858 avss.n857 0.0436892
R11477 avss.n1037 avss.n1036 0.0430541
R11478 avss.n1040 avss.n42 0.0430541
R11479 avss.n1045 avss.n1043 0.0430541
R11480 avss.n1062 avss.n1061 0.0430541
R11481 avss.n1065 avss.n29 0.0430541
R11482 avss.n1084 avss.n1083 0.0430541
R11483 avss.n854 avss.n852 0.0430541
R11484 avss.n651 avss.n628 0.0428468
R11485 avss.n688 avss.n606 0.0428468
R11486 avss.n1080 avss.n1079 0.0427365
R11487 avss.n313 avss 0.0410405
R11488 avss.n742 avss 0.0399737
R11489 avss.n771 avss 0.0399737
R11490 avss.n653 avss.n651 0.0379126
R11491 avss.n707 avss.n606 0.0379126
R11492 avss.n752 avss.n587 0.0358618
R11493 avss.n124 avss 0.0351284
R11494 avss.n136 avss 0.0351284
R11495 avss.n148 avss 0.0351284
R11496 avss.n160 avss 0.0351284
R11497 avss.n172 avss 0.0351284
R11498 avss.n184 avss 0.0351284
R11499 avss.n196 avss 0.0351284
R11500 avss.n208 avss 0.0351284
R11501 avss.n220 avss 0.0351284
R11502 avss.n232 avss 0.0351284
R11503 avss.n244 avss 0.0351284
R11504 avss.n256 avss 0.0351284
R11505 avss.n268 avss 0.0351284
R11506 avss.n280 avss 0.0351284
R11507 avss.n292 avss 0.0351284
R11508 avss avss.n0 0.0351284
R11509 avss.n638 avss.n630 0.0350395
R11510 avss avss.n769 0.0342171
R11511 avss.n838 avss 0.0342171
R11512 avss.n315 avss.n2 0.0334392
R11513 avss.n649 avss.n648 0.0325724
R11514 avss.n664 avss.n663 0.0325724
R11515 avss.n669 avss.n614 0.0325724
R11516 avss.n685 avss 0.0325724
R11517 avss.n692 avss.n691 0.0325724
R11518 avss.n714 avss.n713 0.0325724
R11519 avss.n728 avss.n727 0.0325724
R11520 avss.n738 avss.n737 0.0301053
R11521 avss avss.n740 0.0301053
R11522 avss.n663 avss.n621 0.0276382
R11523 avss.n672 avss.n669 0.0276382
R11524 avss avss.n684 0.0276382
R11525 avss.n693 avss.n687 0.0276382
R11526 avss.n714 avss.n709 0.0276382
R11527 avss.n728 avss.n599 0.0276382
R11528 avss.n315 avss.n314 0.0266824
R11529 avss.n122 avss.n121 0.0266824
R11530 avss.n134 avss.n133 0.0266824
R11531 avss.n146 avss.n145 0.0266824
R11532 avss.n158 avss.n157 0.0266824
R11533 avss.n170 avss.n169 0.0266824
R11534 avss.n182 avss.n181 0.0266824
R11535 avss.n194 avss.n193 0.0266824
R11536 avss.n206 avss.n205 0.0266824
R11537 avss.n218 avss.n217 0.0266824
R11538 avss.n230 avss.n229 0.0266824
R11539 avss.n242 avss.n241 0.0266824
R11540 avss.n254 avss.n253 0.0266824
R11541 avss.n266 avss.n265 0.0266824
R11542 avss.n278 avss.n277 0.0266824
R11543 avss.n290 avss.n289 0.0266824
R11544 avss.n303 avss.n301 0.0266824
R11545 avss.n767 avss.n766 0.0259934
R11546 avss.n770 avss.n568 0.0259934
R11547 avss.n1008 avss.n52 0.0258406
R11548 avss.n1011 avss.n1010 0.0258406
R11549 avss.n753 avss.n752 0.0243487
R11550 avss.n317 avss.n2 0.0224595
R11551 avss.n789 avss.n784 0.0190811
R11552 avss.n391 avss.n386 0.0190811
R11553 avss.n742 avss.n741 0.0177697
R11554 avss.n758 avss.n757 0.016125
R11555 avss.n639 avss.n636 0.0153026
R11556 avss.n666 avss.n619 0.0128355
R11557 avss.n684 avss.n683 0.0128355
R11558 avss.n710 avss.n601 0.0128355
R11559 avss.n740 avss.n593 0.0103684
R11560 avss.n673 avss.n668 0.00790132
R11561 avss.n685 avss.n612 0.00790132
R11562 avss.n725 avss.n724 0.00790132
R11563 avss.n125 avss.n124 0.00641216
R11564 avss.n137 avss.n136 0.00641216
R11565 avss.n149 avss.n148 0.00641216
R11566 avss.n161 avss.n160 0.00641216
R11567 avss.n173 avss.n172 0.00641216
R11568 avss.n185 avss.n184 0.00641216
R11569 avss.n197 avss.n196 0.00641216
R11570 avss.n209 avss.n208 0.00641216
R11571 avss.n221 avss.n220 0.00641216
R11572 avss.n233 avss.n232 0.00641216
R11573 avss.n245 avss.n244 0.00641216
R11574 avss.n257 avss.n256 0.00641216
R11575 avss.n269 avss.n268 0.00641216
R11576 avss.n281 avss.n280 0.00641216
R11577 avss.n293 avss.n292 0.00641216
R11578 avss.n304 avss.n0 0.00641216
R11579 avss.n769 avss.n581 0.00625658
R11580 avss.n839 avss.n838 0.00625658
R11581 avss.n1006 avss.n354 0.004875
R11582 comparator_0.vinn.n7 comparator_0.vinn.t27 51.0275
R11583 comparator_0.vinn.n0 comparator_0.vinn.n29 48.371
R11584 comparator_0.vinn.n1 comparator_0.vinn.n32 48.371
R11585 comparator_0.vinn.n35 comparator_0.vinn.n2 48.371
R11586 comparator_0.vinn.n3 comparator_0.vinn.n10 48.371
R11587 comparator_0.vinn.n4 comparator_0.vinn.n12 48.371
R11588 comparator_0.vinn.n22 comparator_0.vinn.n6 48.371
R11589 comparator_0.vinn.n20 comparator_0.vinn.n7 48.371
R11590 comparator_0.vinn.n8 comparator_0.vinn.n26 48.371
R11591 comparator_0.vinn.n11 comparator_0.vinn.n8 45.4885
R11592 comparator_0.vinn.n25 comparator_0.vinn.n0 45.4885
R11593 comparator_0.vinn.n28 comparator_0.vinn.n1 45.4885
R11594 comparator_0.vinn.n31 comparator_0.vinn.n2 45.4885
R11595 comparator_0.vinn.n3 comparator_0.vinn.n36 45.4885
R11596 comparator_0.vinn.n4 comparator_0.vinn.n23 45.4885
R11597 comparator_0.vinn.n6 comparator_0.vinn.n21 45.4885
R11598 comparator_0.vinn.n53 comparator_0.vinn.n52 45.3881
R11599 comparator_0.vinn.n19 comparator_0.vinn.t24 20.2802
R11600 comparator_0.vinn.n66 comparator_0.vinn.n65 17.7666
R11601 comparator_0.vinn.n63 comparator_0.vinn.n62 17.7666
R11602 comparator_0.vinn.n60 comparator_0.vinn.n59 17.7666
R11603 comparator_0.vinn.n57 comparator_0.vinn.n56 17.7666
R11604 comparator_0.vinn.n13 comparator_0.vinn.n9 17.7666
R11605 comparator_0.vinn.n16 comparator_0.vinn.n15 17.7666
R11606 comparator_0.vinn.n19 comparator_0.vinn.n18 17.7666
R11607 comparator_0.vinn.n53 comparator_0.vinn.n37 17.6963
R11608 comparator_0.vinn.n64 comparator_0.vinn.n63 16.9742
R11609 comparator_0.vinn.n61 comparator_0.vinn.n60 16.9742
R11610 comparator_0.vinn.n58 comparator_0.vinn.n57 16.9742
R11611 comparator_0.vinn.n55 comparator_0.vinn.n54 16.9742
R11612 comparator_0.vinn.n14 comparator_0.vinn.n13 16.9742
R11613 comparator_0.vinn.n17 comparator_0.vinn.n16 16.9742
R11614 comparator_0.vinn.n67 comparator_0.vinn.n66 16.9742
R11615 comparator_0.vinn.n45 comparator_0.vinn.t50 9.72783
R11616 comparator_0.vinn.n38 comparator_0.vinn.t56 9.65028
R11617 comparator_0.vinn.n52 comparator_0.vinn.n44 8.96563
R11618 comparator_0.vinn.n51 comparator_0.vinn.t63 8.73727
R11619 comparator_0.vinn.n50 comparator_0.vinn.t48 8.73727
R11620 comparator_0.vinn.n49 comparator_0.vinn.t52 8.73727
R11621 comparator_0.vinn.n48 comparator_0.vinn.t60 8.73727
R11622 comparator_0.vinn.n47 comparator_0.vinn.t51 8.73727
R11623 comparator_0.vinn.n46 comparator_0.vinn.t57 8.73727
R11624 comparator_0.vinn.n45 comparator_0.vinn.t62 8.73727
R11625 comparator_0.vinn.n44 comparator_0.vinn.t54 8.65985
R11626 comparator_0.vinn.n43 comparator_0.vinn.t55 8.65985
R11627 comparator_0.vinn.n42 comparator_0.vinn.t59 8.65985
R11628 comparator_0.vinn.n41 comparator_0.vinn.t49 8.65985
R11629 comparator_0.vinn.n40 comparator_0.vinn.t58 8.65985
R11630 comparator_0.vinn.n39 comparator_0.vinn.t61 8.65985
R11631 comparator_0.vinn.n38 comparator_0.vinn.t53 8.65985
R11632 comparator_0.vinn.n52 comparator_0.vinn.n51 5.98511
R11633 comparator_0.vinn.t32 comparator_0.vinn.n11 5.5395
R11634 comparator_0.vinn.n11 comparator_0.vinn.t37 5.5395
R11635 comparator_0.vinn.t30 comparator_0.vinn.n25 5.5395
R11636 comparator_0.vinn.n25 comparator_0.vinn.t35 5.5395
R11637 comparator_0.vinn.n29 comparator_0.vinn.t36 5.5395
R11638 comparator_0.vinn.n29 comparator_0.vinn.t34 5.5395
R11639 comparator_0.vinn.t34 comparator_0.vinn.n28 5.5395
R11640 comparator_0.vinn.n28 comparator_0.vinn.t11 5.5395
R11641 comparator_0.vinn.n32 comparator_0.vinn.t10 5.5395
R11642 comparator_0.vinn.n32 comparator_0.vinn.t29 5.5395
R11643 comparator_0.vinn.t29 comparator_0.vinn.n31 5.5395
R11644 comparator_0.vinn.n31 comparator_0.vinn.t21 5.5395
R11645 comparator_0.vinn.n35 comparator_0.vinn.t20 5.5395
R11646 comparator_0.vinn.t47 comparator_0.vinn.n35 5.5395
R11647 comparator_0.vinn.n36 comparator_0.vinn.t47 5.5395
R11648 comparator_0.vinn.n36 comparator_0.vinn.t40 5.5395
R11649 comparator_0.vinn.n10 comparator_0.vinn.t39 5.5395
R11650 comparator_0.vinn.n10 comparator_0.vinn.t33 5.5395
R11651 comparator_0.vinn.n23 comparator_0.vinn.t28 5.5395
R11652 comparator_0.vinn.n23 comparator_0.vinn.t46 5.5395
R11653 comparator_0.vinn.n12 comparator_0.vinn.t45 5.5395
R11654 comparator_0.vinn.n12 comparator_0.vinn.t32 5.5395
R11655 comparator_0.vinn.n21 comparator_0.vinn.t31 5.5395
R11656 comparator_0.vinn.n21 comparator_0.vinn.t4 5.5395
R11657 comparator_0.vinn.n22 comparator_0.vinn.t5 5.5395
R11658 comparator_0.vinn.t28 comparator_0.vinn.n22 5.5395
R11659 comparator_0.vinn.n20 comparator_0.vinn.t26 5.5395
R11660 comparator_0.vinn.t31 comparator_0.vinn.n20 5.5395
R11661 comparator_0.vinn.n26 comparator_0.vinn.t38 5.5395
R11662 comparator_0.vinn.n26 comparator_0.vinn.t30 5.5395
R11663 comparator_0.vinn.n34 comparator_0.vinn.n3 3.79433
R11664 comparator_0.vinn.n7 comparator_0.vinn.n5 3.79433
R11665 comparator_0.vinn.n2 comparator_0.vinn.n34 3.4105
R11666 comparator_0.vinn.n33 comparator_0.vinn.n1 3.4105
R11667 comparator_0.vinn.n30 comparator_0.vinn.n0 3.4105
R11668 comparator_0.vinn.n6 comparator_0.vinn.n5 3.4105
R11669 comparator_0.vinn.n24 comparator_0.vinn.n4 3.4105
R11670 comparator_0.vinn.n27 comparator_0.vinn.n8 3.4105
R11671 comparator_0.vinn.n65 comparator_0.vinn.t2 3.3065
R11672 comparator_0.vinn.n65 comparator_0.vinn.t15 3.3065
R11673 comparator_0.vinn.t15 comparator_0.vinn.n64 3.3065
R11674 comparator_0.vinn.n64 comparator_0.vinn.t7 3.3065
R11675 comparator_0.vinn.n62 comparator_0.vinn.t6 3.3065
R11676 comparator_0.vinn.n62 comparator_0.vinn.t18 3.3065
R11677 comparator_0.vinn.t18 comparator_0.vinn.n61 3.3065
R11678 comparator_0.vinn.n61 comparator_0.vinn.t43 3.3065
R11679 comparator_0.vinn.n59 comparator_0.vinn.t44 3.3065
R11680 comparator_0.vinn.n59 comparator_0.vinn.t16 3.3065
R11681 comparator_0.vinn.t16 comparator_0.vinn.n58 3.3065
R11682 comparator_0.vinn.n58 comparator_0.vinn.t1 3.3065
R11683 comparator_0.vinn.n56 comparator_0.vinn.t0 3.3065
R11684 comparator_0.vinn.n56 comparator_0.vinn.t14 3.3065
R11685 comparator_0.vinn.t14 comparator_0.vinn.n55 3.3065
R11686 comparator_0.vinn.n55 comparator_0.vinn.t42 3.3065
R11687 comparator_0.vinn.n37 comparator_0.vinn.t41 3.3065
R11688 comparator_0.vinn.n37 comparator_0.vinn.t12 3.3065
R11689 comparator_0.vinn.t17 comparator_0.vinn.n14 3.3065
R11690 comparator_0.vinn.n14 comparator_0.vinn.t23 3.3065
R11691 comparator_0.vinn.n9 comparator_0.vinn.t22 3.3065
R11692 comparator_0.vinn.t19 comparator_0.vinn.n9 3.3065
R11693 comparator_0.vinn.t13 comparator_0.vinn.n17 3.3065
R11694 comparator_0.vinn.n17 comparator_0.vinn.t9 3.3065
R11695 comparator_0.vinn.n15 comparator_0.vinn.t8 3.3065
R11696 comparator_0.vinn.n15 comparator_0.vinn.t17 3.3065
R11697 comparator_0.vinn.n18 comparator_0.vinn.t25 3.3065
R11698 comparator_0.vinn.n18 comparator_0.vinn.t13 3.3065
R11699 comparator_0.vinn.t19 comparator_0.vinn.n67 3.3065
R11700 comparator_0.vinn.n67 comparator_0.vinn.t3 3.3065
R11701 comparator_0.vinn.n66 comparator_0.vinn.n8 1.98488
R11702 comparator_0.vinn.n7 comparator_0.vinn.n19 1.98488
R11703 comparator_0.vinn.n6 comparator_0.vinn.n16 1.98488
R11704 comparator_0.vinn.n4 comparator_0.vinn.n13 1.98488
R11705 comparator_0.vinn.n54 comparator_0.vinn.n3 1.98488
R11706 comparator_0.vinn.n57 comparator_0.vinn.n2 1.98488
R11707 comparator_0.vinn.n60 comparator_0.vinn.n1 1.98488
R11708 comparator_0.vinn.n63 comparator_0.vinn.n0 1.98488
R11709 comparator_0.vinn.n51 comparator_0.vinn.n50 0.99106
R11710 comparator_0.vinn.n50 comparator_0.vinn.n49 0.99106
R11711 comparator_0.vinn.n49 comparator_0.vinn.n48 0.99106
R11712 comparator_0.vinn.n48 comparator_0.vinn.n47 0.99106
R11713 comparator_0.vinn.n47 comparator_0.vinn.n46 0.99106
R11714 comparator_0.vinn.n46 comparator_0.vinn.n45 0.99106
R11715 comparator_0.vinn.n44 comparator_0.vinn.n43 0.99093
R11716 comparator_0.vinn.n43 comparator_0.vinn.n42 0.99093
R11717 comparator_0.vinn.n42 comparator_0.vinn.n41 0.99093
R11718 comparator_0.vinn.n41 comparator_0.vinn.n40 0.99093
R11719 comparator_0.vinn.n40 comparator_0.vinn.n39 0.99093
R11720 comparator_0.vinn.n39 comparator_0.vinn.n38 0.99093
R11721 comparator_0.vinn.n34 comparator_0.vinn.n33 0.384333
R11722 comparator_0.vinn.n33 comparator_0.vinn.n30 0.384333
R11723 comparator_0.vinn.n30 comparator_0.vinn.n27 0.384333
R11724 comparator_0.vinn.n24 comparator_0.vinn.n5 0.384333
R11725 comparator_0.vinn.n27 comparator_0.vinn.n24 0.384333
R11726 comparator_0.vinn.n54 comparator_0.vinn.n53 0.0708125
R11727 rstring_mux_0.vtrip4.n5 rstring_mux_0.vtrip4.n3 50.7022
R11728 rstring_mux_0.vtrip4.n2 rstring_mux_0.vtrip4.n0 50.7022
R11729 rstring_mux_0.vtrip4.n7 rstring_mux_0.vtrip4.n6 24.0569
R11730 rstring_mux_0.vtrip4.n6 rstring_mux_0.vtrip4.n2 14.0584
R11731 rstring_mux_0.vtrip4.n5 rstring_mux_0.vtrip4.n4 13.8791
R11732 rstring_mux_0.vtrip4.n2 rstring_mux_0.vtrip4.n1 13.8791
R11733 rstring_mux_0.vtrip4 rstring_mux_0.vtrip4.t7 10.5739
R11734 rstring_mux_0.vtrip4.n3 rstring_mux_0.vtrip4.t3 5.5395
R11735 rstring_mux_0.vtrip4.n3 rstring_mux_0.vtrip4.t4 5.5395
R11736 rstring_mux_0.vtrip4.n0 rstring_mux_0.vtrip4.t9 5.5395
R11737 rstring_mux_0.vtrip4.n0 rstring_mux_0.vtrip4.t8 5.5395
R11738 rstring_mux_0.vtrip4.n6 rstring_mux_0.vtrip4.n5 3.33746
R11739 rstring_mux_0.vtrip4.n4 rstring_mux_0.vtrip4.t6 3.3065
R11740 rstring_mux_0.vtrip4.n4 rstring_mux_0.vtrip4.t5 3.3065
R11741 rstring_mux_0.vtrip4.n1 rstring_mux_0.vtrip4.t1 3.3065
R11742 rstring_mux_0.vtrip4.n1 rstring_mux_0.vtrip4.t2 3.3065
R11743 rstring_mux_0.vtrip4.n7 rstring_mux_0.vtrip4.t0 0.826075
R11744 rstring_mux_0.vtrip4 rstring_mux_0.vtrip4.n7 0.0563195
R11745 avdd.n1705 avdd.n1661 99969.2
R11746 avdd.n1705 avdd.n1704 83663.1
R11747 avdd.n1689 avdd.n1662 66867
R11748 avdd.n1690 avdd.n1663 60783.5
R11749 avdd.n1689 avdd.n1688 60384.8
R11750 avdd.n1678 avdd.n1661 58787
R11751 avdd.n1702 avdd.n1663 52810.3
R11752 avdd.n1703 avdd.n1662 50831
R11753 avdd.n1706 avdd.n1659 49200
R11754 avdd.n1688 avdd.n1687 47131.3
R11755 avdd.n1706 avdd.n1660 41239.5
R11756 avdd.n1690 avdd.n1668 29875.1
R11757 avdd.n1679 avdd.n1659 29132.4
R11758 avdd.n1704 avdd.n1703 27601.7
R11759 avdd.n1678 avdd.n1669 27058.6
R11760 avdd.n1179 avdd.n1052 25108.6
R11761 avdd.n1177 avdd.n1052 25108.6
R11762 avdd.n1601 avdd.n1298 25108.6
R11763 avdd.n1599 avdd.n1298 25108.6
R11764 avdd.n1179 avdd.n1178 25105.2
R11765 avdd.n1178 avdd.n1177 25105.2
R11766 avdd.n1601 avdd.n1600 25105.2
R11767 avdd.n1600 avdd.n1599 25105.2
R11768 avdd.n1686 avdd.n1668 22957.3
R11769 avdd.n1687 avdd.n1669 17438.8
R11770 avdd.n1757 avdd.n1750 15077.5
R11771 avdd.n1757 avdd.n1751 15077.5
R11772 avdd.n1794 avdd.n1751 15077.5
R11773 avdd.n1794 avdd.n1750 15077.5
R11774 avdd.n1702 avdd.n1660 13877.8
R11775 avdd.n1679 avdd.n1670 13642.7
R11776 avdd.n1180 avdd.n1050 12653.5
R11777 avdd.n1176 avdd.n1050 12653.5
R11778 avdd.n1602 avdd.n1296 12653.5
R11779 avdd.n1598 avdd.n1296 12653.5
R11780 avdd.n1180 avdd.n1051 12651.9
R11781 avdd.n1176 avdd.n1051 12651.9
R11782 avdd.n1602 avdd.n1297 12651.9
R11783 avdd.n1598 avdd.n1297 12651.9
R11784 avdd.n1200 avdd.n997 11582.8
R11785 avdd.n1160 avdd.n997 11582.8
R11786 avdd.n1622 avdd.n1243 11582.8
R11787 avdd.n1582 avdd.n1243 11582.8
R11788 avdd.n1202 avdd.n994 10507.7
R11789 avdd.n1162 avdd.n994 10507.7
R11790 avdd.n1624 avdd.n1240 10507.7
R11791 avdd.n1584 avdd.n1240 10507.7
R11792 avdd.n1194 avdd.n1014 10039.9
R11793 avdd.n1194 avdd.n993 10039.9
R11794 avdd.n1196 avdd.n1013 10039.9
R11795 avdd.n1196 avdd.n998 10039.9
R11796 avdd.n1616 avdd.n1260 10039.9
R11797 avdd.n1616 avdd.n1239 10039.9
R11798 avdd.n1618 avdd.n1259 10039.9
R11799 avdd.n1618 avdd.n1244 10039.9
R11800 avdd.n1858 avdd.n727 9739.14
R11801 avdd.n1858 avdd.n728 9739.14
R11802 avdd.n1857 avdd.n728 9739.14
R11803 avdd.n1857 avdd.n727 9739.14
R11804 avdd.n1686 avdd.n1670 8461.62
R11805 avdd.n1692 avdd.n1664 8070.02
R11806 avdd.n1691 avdd.n1667 6943.25
R11807 avdd.n1677 avdd.n1676 6761.04
R11808 avdd.n1701 avdd.n1664 6168.09
R11809 avdd.n1684 avdd.n1672 5303.72
R11810 avdd.n1697 avdd.n1696 4892.23
R11811 avdd.n1708 avdd.n1657 4681.79
R11812 avdd.n1674 avdd.n1657 4335.44
R11813 avdd.n1842 avdd.n1841 4316.28
R11814 avdd.n1844 avdd.n1841 4316.28
R11815 avdd.n1842 avdd.n1838 4316.28
R11816 avdd.n1844 avdd.n1838 4316.28
R11817 avdd.n1700 avdd.n1665 3225.22
R11818 avdd.n1681 avdd.n1680 3163.48
R11819 avdd.n1809 avdd.n1722 3160.55
R11820 avdd.n1810 avdd.n1722 3160.55
R11821 avdd.n1181 avdd.n1049 2933.46
R11822 avdd.n1603 avdd.n1295 2933.46
R11823 avdd.n1175 avdd.n1053 2922.54
R11824 avdd.n1597 avdd.n1299 2922.54
R11825 avdd.n1793 avdd.n1752 2890.84
R11826 avdd.n1758 avdd.n1752 2890.84
R11827 avdd.n1174 avdd.n1054 2865.69
R11828 avdd.n1596 avdd.n1300 2865.69
R11829 avdd.n1759 avdd.n1753 2860.42
R11830 avdd.n1792 avdd.n1753 2860.42
R11831 avdd.n1182 avdd.n1048 2841.22
R11832 avdd.n1604 avdd.n1294 2841.22
R11833 avdd.n1158 avdd.n1013 2620.03
R11834 avdd.n1158 avdd.n1014 2620.03
R11835 avdd.n998 avdd.n995 2620.03
R11836 avdd.n995 avdd.n993 2620.03
R11837 avdd.n1580 avdd.n1259 2620.03
R11838 avdd.n1580 avdd.n1260 2620.03
R11839 avdd.n1244 avdd.n1241 2620.03
R11840 avdd.n1241 avdd.n1239 2620.03
R11841 avdd.n1803 avdd.n1729 2513.9
R11842 avdd.n1803 avdd.n1721 2513.9
R11843 avdd.n1804 avdd.n1726 2513.9
R11844 avdd.n1804 avdd.n1723 2513.9
R11845 avdd.n1696 avdd.n1658 2495.62
R11846 avdd.n1156 avdd.n1071 2480.48
R11847 avdd.n1156 avdd.n1072 2480.48
R11848 avdd.n1071 avdd.n1070 2480.48
R11849 avdd.n1072 avdd.n1070 2480.48
R11850 avdd.n1578 avdd.n1317 2480.48
R11851 avdd.n1578 avdd.n1318 2480.48
R11852 avdd.n1317 avdd.n1316 2480.48
R11853 avdd.n1318 avdd.n1316 2480.48
R11854 avdd.n1708 avdd.n1707 2412.42
R11855 avdd.n1798 avdd.n1746 2346.83
R11856 avdd.n1797 avdd.n1746 2346.83
R11857 avdd.n1159 avdd.n999 2223.06
R11858 avdd.n1199 avdd.n999 2223.06
R11859 avdd.n1581 avdd.n1245 2223.06
R11860 avdd.n1621 avdd.n1245 2223.06
R11861 avdd.n1707 avdd.n1658 2115.76
R11862 avdd.n1007 avdd.n1006 2059.86
R11863 avdd.n1006 avdd.n1005 2059.86
R11864 avdd.n1005 avdd.n1002 2059.86
R11865 avdd.n1007 avdd.n1002 2059.86
R11866 avdd.n1253 avdd.n1252 2059.86
R11867 avdd.n1252 avdd.n1251 2059.86
R11868 avdd.n1251 avdd.n1248 2059.86
R11869 avdd.n1253 avdd.n1248 2059.86
R11870 avdd.n1203 avdd.n992 2000.19
R11871 avdd.n1163 avdd.n992 2000.19
R11872 avdd.n1625 avdd.n1238 2000.19
R11873 avdd.n1585 avdd.n1238 2000.19
R11874 avdd.n1685 avdd.n1671 1971.95
R11875 avdd.n1197 avdd.n1011 1923.01
R11876 avdd.n1198 avdd.n1197 1923.01
R11877 avdd.n1619 avdd.n1257 1923.01
R11878 avdd.n1620 avdd.n1619 1923.01
R11879 avdd.n1810 avdd.n1721 1837.76
R11880 avdd.n1809 avdd.n1723 1837.76
R11881 avdd.n729 avdd.n725 1616.56
R11882 avdd.n1855 avdd.n730 1616.56
R11883 avdd.n730 avdd.n726 1616.56
R11884 avdd.n1860 avdd.n725 1615.06
R11885 avdd.n1200 avdd.n998 1542.93
R11886 avdd.n1160 avdd.n1013 1542.93
R11887 avdd.n1622 avdd.n1244 1542.93
R11888 avdd.n1582 avdd.n1259 1542.93
R11889 avdd.n1748 avdd.n1726 1322.79
R11890 avdd.n1748 avdd.n1729 1322.79
R11891 avdd.n1727 avdd.n1723 1322.79
R11892 avdd.n1727 avdd.n1721 1322.79
R11893 avdd.n1193 avdd.n1015 1237.08
R11894 avdd.n1193 avdd.n990 1237.08
R11895 avdd.n1615 avdd.n1261 1237.08
R11896 avdd.n1615 avdd.n1236 1237.08
R11897 avdd.n1798 avdd.n1729 1024.03
R11898 avdd.n1797 avdd.n1726 1024.03
R11899 avdd.n1846 avdd.n1845 831.247
R11900 avdd.n1846 avdd.n1837 831.247
R11901 avdd.n107 avdd.t44 692.692
R11902 avdd.n444 avdd.t447 692.692
R11903 avdd avdd.t43 688.231
R11904 avdd avdd.t46 688.231
R11905 avdd.n1840 avdd.n1839 682.918
R11906 avdd.n1840 avdd.n1820 682.918
R11907 avdd.n32 avdd.t162 648.668
R11908 avdd.n368 avdd.t654 648.668
R11909 avdd.n340 avdd.t437 648.668
R11910 avdd.n312 avdd.t13 648.668
R11911 avdd.n284 avdd.t512 648.668
R11912 avdd.n256 avdd.t441 648.668
R11913 avdd.n228 avdd.t216 648.668
R11914 avdd.n200 avdd.t411 648.668
R11915 avdd.n172 avdd.t503 648.668
R11916 avdd.n144 avdd.t212 648.668
R11917 avdd.n705 avdd.t657 648.668
R11918 avdd.n677 avdd.t1 648.668
R11919 avdd.n649 avdd.t154 648.668
R11920 avdd.n621 avdd.t145 648.668
R11921 avdd.n593 avdd.t399 648.668
R11922 avdd.n565 avdd.t594 648.668
R11923 avdd.n537 avdd.t626 648.668
R11924 avdd.n509 avdd.t41 648.668
R11925 avdd.n481 avdd.t132 648.668
R11926 avdd.n957 avdd.n740 624.808
R11927 avdd.n955 avdd.n741 624.808
R11928 avdd.n944 avdd.n943 624.808
R11929 avdd.n932 avdd.n760 624.808
R11930 avdd.n930 avdd.n761 624.808
R11931 avdd.n919 avdd.n918 624.808
R11932 avdd.n907 avdd.n780 624.808
R11933 avdd.n905 avdd.n781 624.808
R11934 avdd.n894 avdd.n893 624.808
R11935 avdd.n882 avdd.n800 624.808
R11936 avdd.n880 avdd.n801 624.808
R11937 avdd.n869 avdd.n868 624.808
R11938 avdd.n857 avdd.n820 624.808
R11939 avdd.n855 avdd.n821 624.808
R11940 avdd.n844 avdd.n843 624.808
R11941 avdd.n1165 avdd.n1015 612.894
R11942 avdd.n1205 avdd.n990 612.894
R11943 avdd.n1587 avdd.n1261 612.894
R11944 avdd.n1627 avdd.n1236 612.894
R11945 avdd.n1808 avdd.n1719 609.883
R11946 avdd.n1812 avdd.n1811 555.672
R11947 avdd.t426 avdd.t424 511.356
R11948 avdd.t330 avdd.t432 511.356
R11949 avdd.t400 avdd.t330 511.356
R11950 avdd.t402 avdd.t400 511.356
R11951 avdd.t341 avdd.t402 511.356
R11952 avdd.t404 avdd.t341 511.356
R11953 avdd.t406 avdd.t404 511.356
R11954 avdd.t258 avdd.t406 511.356
R11955 avdd.n1164 avdd.n1069 506.353
R11956 avdd.n1586 avdd.n1315 506.353
R11957 avdd.n715 avdd.t513 499.882
R11958 avdd.t165 avdd.t169 484.288
R11959 avdd.t141 avdd.t167 484.288
R11960 avdd.t527 avdd.t519 484.288
R11961 avdd.t446 avdd.t525 484.288
R11962 avdd.n1802 avdd.n1800 481.507
R11963 avdd.n1805 avdd.n1725 481.507
R11964 avdd.n1076 avdd.n1075 479.625
R11965 avdd.n1075 avdd.n1074 479.625
R11966 avdd.n1322 avdd.n1321 479.625
R11967 avdd.n1321 avdd.n1320 479.625
R11968 avdd.t424 avdd.t428 475.098
R11969 avdd.n1202 avdd.n993 467.793
R11970 avdd.n1162 avdd.n1014 467.793
R11971 avdd.n1624 avdd.n1239 467.793
R11972 avdd.n1584 avdd.n1260 467.793
R11973 avdd.n1796 avdd.n1745 454.024
R11974 avdd.n1005 avdd.t141 437.699
R11975 avdd.n1251 avdd.t446 437.699
R11976 avdd.n1155 avdd.n1073 437.082
R11977 avdd.n1155 avdd.n1154 437.082
R11978 avdd.n1577 avdd.n1319 437.082
R11979 avdd.n1577 avdd.n1576 437.082
R11980 avdd.n1799 avdd.n1745 423.818
R11981 avdd.n1008 avdd.n1001 399.06
R11982 avdd.n1004 avdd.n1001 399.06
R11983 avdd.n1254 avdd.n1247 399.06
R11984 avdd.n1250 avdd.n1247 399.06
R11985 avdd.n1733 avdd.t337 397.264
R11986 avdd.n1734 avdd.t347 397.135
R11987 avdd.n1735 avdd.t227 397.135
R11988 avdd.n724 avdd.t247 388.149
R11989 avdd.n968 avdd.t359 388.149
R11990 avdd.n969 avdd.t394 388.149
R11991 avdd.n970 avdd.t390 388.149
R11992 avdd.n971 avdd.t296 388.149
R11993 avdd.n972 avdd.t378 388.149
R11994 avdd.n973 avdd.t367 388.149
R11995 avdd.n974 avdd.t380 388.149
R11996 avdd.n976 avdd.t392 388.149
R11997 avdd.n977 avdd.t261 388.149
R11998 avdd.n978 avdd.t374 388.149
R11999 avdd.n979 avdd.t274 388.149
R12000 avdd.n980 avdd.t332 388.149
R12001 avdd.n981 avdd.t242 388.149
R12002 avdd.n982 avdd.t303 388.149
R12003 avdd.n28 avdd.t7 372.885
R12004 avdd.n364 avdd.t160 372.885
R12005 avdd.n336 avdd.t152 372.885
R12006 avdd.n308 avdd.t493 372.885
R12007 avdd.n280 avdd.t150 372.885
R12008 avdd.n252 avdd.t423 372.885
R12009 avdd.n224 avdd.t100 372.885
R12010 avdd.n196 avdd.t104 372.885
R12011 avdd.n168 avdd.t124 372.885
R12012 avdd.n140 avdd.t136 372.885
R12013 avdd.n701 avdd.t589 372.885
R12014 avdd.n673 avdd.t92 372.885
R12015 avdd.n645 avdd.t174 372.885
R12016 avdd.n617 avdd.t143 372.885
R12017 avdd.n589 avdd.t35 372.885
R12018 avdd.n561 avdd.t620 372.885
R12019 avdd.n533 avdd.t37 372.885
R12020 avdd.n505 avdd.t587 372.885
R12021 avdd.n477 avdd.t571 372.885
R12022 avdd.t408 avdd.n732 354.904
R12023 avdd.n1811 avdd.n1720 352
R12024 avdd.n1808 avdd.n1807 352
R12025 avdd.n1757 avdd.t258 345.817
R12026 avdd.n1007 avdd.t165 343.495
R12027 avdd.n1253 avdd.t527 343.495
R12028 avdd.n1801 avdd.n1720 325.647
R12029 avdd.n1807 avdd.n1806 325.647
R12030 avdd.n1375 avdd.n1374 325.039
R12031 avdd.n1071 avdd.t53 323.445
R12032 avdd.n1072 avdd.t418 323.445
R12033 avdd.n1317 avdd.t24 323.445
R12034 avdd.n1318 avdd.t582 323.445
R12035 avdd.n21 avdd.n5 321.882
R12036 avdd.n11 avdd.n10 321.882
R12037 avdd.n23 avdd.n2 321.882
R12038 avdd.n357 avdd.n40 321.882
R12039 avdd.n343 avdd.n342 321.882
R12040 avdd.n38 avdd.n36 321.882
R12041 avdd.n329 avdd.n48 321.882
R12042 avdd.n315 avdd.n314 321.882
R12043 avdd.n46 avdd.n44 321.882
R12044 avdd.n301 avdd.n56 321.882
R12045 avdd.n287 avdd.n286 321.882
R12046 avdd.n54 avdd.n52 321.882
R12047 avdd.n273 avdd.n64 321.882
R12048 avdd.n259 avdd.n258 321.882
R12049 avdd.n62 avdd.n60 321.882
R12050 avdd.n245 avdd.n72 321.882
R12051 avdd.n231 avdd.n230 321.882
R12052 avdd.n70 avdd.n68 321.882
R12053 avdd.n217 avdd.n80 321.882
R12054 avdd.n203 avdd.n202 321.882
R12055 avdd.n78 avdd.n76 321.882
R12056 avdd.n189 avdd.n88 321.882
R12057 avdd.n175 avdd.n174 321.882
R12058 avdd.n86 avdd.n84 321.882
R12059 avdd.n161 avdd.n96 321.882
R12060 avdd.n147 avdd.n146 321.882
R12061 avdd.n94 avdd.n92 321.882
R12062 avdd.n109 avdd.n104 321.882
R12063 avdd.n126 avdd.n104 321.882
R12064 avdd.n126 avdd.n101 321.882
R12065 avdd.n130 avdd.n101 321.882
R12066 avdd.n131 avdd.n130 321.882
R12067 avdd.n131 avdd.n100 321.882
R12068 avdd.n135 avdd.n100 321.882
R12069 avdd.n694 avdd.n377 321.882
R12070 avdd.n680 avdd.n679 321.882
R12071 avdd.n375 avdd.n373 321.882
R12072 avdd.n666 avdd.n385 321.882
R12073 avdd.n652 avdd.n651 321.882
R12074 avdd.n383 avdd.n381 321.882
R12075 avdd.n638 avdd.n393 321.882
R12076 avdd.n624 avdd.n623 321.882
R12077 avdd.n391 avdd.n389 321.882
R12078 avdd.n610 avdd.n401 321.882
R12079 avdd.n596 avdd.n595 321.882
R12080 avdd.n399 avdd.n397 321.882
R12081 avdd.n582 avdd.n409 321.882
R12082 avdd.n568 avdd.n567 321.882
R12083 avdd.n407 avdd.n405 321.882
R12084 avdd.n554 avdd.n417 321.882
R12085 avdd.n540 avdd.n539 321.882
R12086 avdd.n415 avdd.n413 321.882
R12087 avdd.n526 avdd.n425 321.882
R12088 avdd.n512 avdd.n511 321.882
R12089 avdd.n423 avdd.n421 321.882
R12090 avdd.n498 avdd.n433 321.882
R12091 avdd.n484 avdd.n483 321.882
R12092 avdd.n431 avdd.n429 321.882
R12093 avdd.n446 avdd.n441 321.882
R12094 avdd.n463 avdd.n438 321.882
R12095 avdd.n467 avdd.n438 321.882
R12096 avdd.n468 avdd.n467 321.882
R12097 avdd.n468 avdd.n437 321.882
R12098 avdd.n472 avdd.n437 321.882
R12099 avdd.n714 avdd.n713 321.882
R12100 avdd.n1373 avdd.n1370 321.882
R12101 avdd.n1379 avdd.n1370 321.882
R12102 avdd.n1379 avdd.n1368 321.882
R12103 avdd.n1384 avdd.n1368 321.882
R12104 avdd.n1384 avdd.n1364 321.882
R12105 avdd.n1390 avdd.n1364 321.882
R12106 avdd.n1390 avdd.n1363 321.882
R12107 avdd.n1394 avdd.n1363 321.882
R12108 avdd.n1394 avdd.n1359 321.882
R12109 avdd.n1400 avdd.n1359 321.882
R12110 avdd.n1400 avdd.n1357 321.882
R12111 avdd.n1405 avdd.n1357 321.882
R12112 avdd.n1405 avdd.n1353 321.882
R12113 avdd.n1411 avdd.n1353 321.882
R12114 avdd.n1411 avdd.n1352 321.882
R12115 avdd.n1415 avdd.n1352 321.882
R12116 avdd.n1415 avdd.n1348 321.882
R12117 avdd.n1421 avdd.n1348 321.882
R12118 avdd.n1421 avdd.n1346 321.882
R12119 avdd.n1426 avdd.n1346 321.882
R12120 avdd.n1426 avdd.n1342 321.882
R12121 avdd.n1432 avdd.n1342 321.882
R12122 avdd.n1432 avdd.n1341 321.882
R12123 avdd.n1437 avdd.n1341 321.882
R12124 avdd.n1437 avdd.n1337 321.882
R12125 avdd.n1443 avdd.n1337 321.882
R12126 avdd.n1443 avdd.n1336 321.882
R12127 avdd.n1448 avdd.n1336 321.882
R12128 avdd.n1448 avdd.n1331 321.882
R12129 avdd.n1475 avdd.n1331 321.882
R12130 avdd.n1475 avdd.n1329 321.882
R12131 avdd.n1479 avdd.n1329 321.882
R12132 avdd.n1480 avdd.n1479 321.882
R12133 avdd.n1480 avdd.n1325 321.882
R12134 avdd.n1326 avdd.n1325 321.882
R12135 avdd.n1328 avdd.n1326 321.882
R12136 avdd.n842 avdd.n826 321.882
R12137 avdd.n847 avdd.n846 321.882
R12138 avdd.n846 avdd.n825 321.882
R12139 avdd.n858 avdd.n817 321.882
R12140 avdd.n854 avdd.n817 321.882
R12141 avdd.n867 avdd.n806 321.882
R12142 avdd.n819 avdd.n806 321.882
R12143 avdd.n872 avdd.n871 321.882
R12144 avdd.n871 avdd.n805 321.882
R12145 avdd.n883 avdd.n797 321.882
R12146 avdd.n879 avdd.n797 321.882
R12147 avdd.n892 avdd.n786 321.882
R12148 avdd.n799 avdd.n786 321.882
R12149 avdd.n897 avdd.n896 321.882
R12150 avdd.n896 avdd.n785 321.882
R12151 avdd.n908 avdd.n777 321.882
R12152 avdd.n904 avdd.n777 321.882
R12153 avdd.n917 avdd.n766 321.882
R12154 avdd.n779 avdd.n766 321.882
R12155 avdd.n922 avdd.n921 321.882
R12156 avdd.n921 avdd.n765 321.882
R12157 avdd.n933 avdd.n757 321.882
R12158 avdd.n929 avdd.n757 321.882
R12159 avdd.n942 avdd.n746 321.882
R12160 avdd.n759 avdd.n746 321.882
R12161 avdd.n947 avdd.n946 321.882
R12162 avdd.n946 avdd.n745 321.882
R12163 avdd.n958 avdd.n738 321.882
R12164 avdd.n954 avdd.n738 321.882
R12165 avdd.n733 avdd.n732 321.882
R12166 avdd.n734 avdd.n733 321.882
R12167 avdd.n1485 avdd.n1484 318.757
R12168 avdd.n834 avdd.n833 318.757
R12169 avdd.n463 avdd.n441 318.529
R12170 avdd.t240 avdd.t182 310.303
R12171 avdd.t182 avdd.t186 310.303
R12172 avdd.t179 avdd.t177 310.303
R12173 avdd.t177 avdd.t221 310.303
R12174 avdd.t234 avdd.t80 310.303
R12175 avdd.t80 avdd.t73 310.303
R12176 avdd.t65 avdd.t63 310.303
R12177 avdd.t63 avdd.t230 310.303
R12178 avdd.n1159 avdd.n1011 300.048
R12179 avdd.n1199 avdd.n1198 300.048
R12180 avdd.n1009 avdd.n1000 300.048
R12181 avdd.n1003 avdd.n1000 300.048
R12182 avdd.n1581 avdd.n1257 300.048
R12183 avdd.n1621 avdd.n1620 300.048
R12184 avdd.n1255 avdd.n1246 300.048
R12185 avdd.n1249 avdd.n1246 300.048
R12186 avdd.n1068 avdd.n1011 295.529
R12187 avdd.n1314 avdd.n1257 295.529
R12188 avdd.t169 avdd.n996 289.247
R12189 avdd.t519 avdd.n1242 289.247
R12190 avdd.n1204 avdd.n991 281.601
R12191 avdd.n1626 avdd.n1237 281.601
R12192 avdd.n1466 avdd.t541 280.161
R12193 avdd.n1459 avdd.t543 279.486
R12194 avdd.n360 avdd.n359 271.068
R12195 avdd.n332 avdd.n331 271.068
R12196 avdd.n304 avdd.n303 271.068
R12197 avdd.n276 avdd.n275 271.068
R12198 avdd.n248 avdd.n247 271.068
R12199 avdd.n220 avdd.n219 271.068
R12200 avdd.n192 avdd.n191 271.068
R12201 avdd.n164 avdd.n163 271.068
R12202 avdd.n697 avdd.n696 271.068
R12203 avdd.n669 avdd.n668 271.068
R12204 avdd.n641 avdd.n640 271.068
R12205 avdd.n613 avdd.n612 271.068
R12206 avdd.n585 avdd.n584 271.068
R12207 avdd.n557 avdd.n556 271.068
R12208 avdd.n529 avdd.n528 271.068
R12209 avdd.n501 avdd.n500 271.068
R12210 avdd.n717 avdd.n716 271.068
R12211 avdd.n1807 avdd.n1724 257.882
R12212 avdd.n1747 avdd.n1725 257.882
R12213 avdd.n1493 avdd.t591 257.603
R12214 avdd.n1467 avdd.t114 256.101
R12215 avdd.n1756 avdd.t426 255.679
R12216 avdd.t432 avdd.n1756 255.679
R12217 avdd.n721 avdd.t514 252.983
R12218 avdd.n1495 avdd.t120 252.983
R12219 avdd.n837 avdd.t501 252.983
R12220 avdd.n830 avdd.t487 252.983
R12221 avdd.n850 avdd.t537 252.983
R12222 avdd.n862 avdd.t219 252.983
R12223 avdd.n810 avdd.t112 252.983
R12224 avdd.n875 avdd.t623 252.983
R12225 avdd.n887 avdd.t495 252.983
R12226 avdd.n790 avdd.t126 252.983
R12227 avdd.n900 avdd.t573 252.983
R12228 avdd.n912 avdd.t9 252.983
R12229 avdd.n770 avdd.t575 252.983
R12230 avdd.n925 avdd.t106 252.983
R12231 avdd.n937 avdd.t17 252.983
R12232 avdd.n750 avdd.t206 252.983
R12233 avdd.n950 avdd.t122 252.983
R12234 avdd.n961 avdd.t409 252.983
R12235 avdd.n1860 avdd.n1859 241.459
R12236 avdd.n1856 avdd.n729 240.66
R12237 avdd.n1856 avdd.n1855 240.66
R12238 avdd.n1859 avdd.n726 240.66
R12239 avdd.t53 avdd.t47 233.565
R12240 avdd.t47 avdd.t57 233.565
R12241 avdd.t57 avdd.t55 233.565
R12242 avdd.t55 avdd.t49 233.565
R12243 avdd.t51 avdd.t59 233.565
R12244 avdd.t61 avdd.t51 233.565
R12245 avdd.t420 avdd.t61 233.565
R12246 avdd.t418 avdd.t420 233.565
R12247 avdd.t24 avdd.t28 233.565
R12248 avdd.t28 avdd.t32 233.565
R12249 avdd.t32 avdd.t18 233.565
R12250 avdd.t18 avdd.t22 233.565
R12251 avdd.t20 avdd.t30 233.565
R12252 avdd.t26 avdd.t20 233.565
R12253 avdd.t584 avdd.t26 233.565
R12254 avdd.t582 avdd.t584 233.565
R12255 avdd.n1230 avdd.t168 232.686
R12256 avdd.n1652 avdd.t526 232.686
R12257 avdd.n1144 avdd.t54 231.989
R12258 avdd.n1153 avdd.t419 231.989
R12259 avdd.n1566 avdd.t25 231.989
R12260 avdd.n1575 avdd.t583 231.989
R12261 avdd.n1231 avdd.t166 231.974
R12262 avdd.n1230 avdd.t170 231.974
R12263 avdd.n1653 avdd.t528 231.974
R12264 avdd.n1652 avdd.t520 231.974
R12265 avdd.n1227 avdd.t246 227.478
R12266 avdd.n1225 avdd.t256 227.478
R12267 avdd.n1223 avdd.t253 227.478
R12268 avdd.n1221 avdd.t290 227.478
R12269 avdd.n1219 avdd.t310 227.478
R12270 avdd.n1217 avdd.t313 227.478
R12271 avdd.n1215 avdd.t328 227.478
R12272 avdd.n1213 avdd.t323 227.478
R12273 avdd.n1211 avdd.t384 227.478
R12274 avdd.n1209 avdd.t336 227.478
R12275 avdd.n1207 avdd.t389 227.478
R12276 avdd.n1140 avdd.t277 227.478
R12277 avdd.t284 avdd.n1135 227.478
R12278 avdd.t282 avdd.n1132 227.478
R12279 avdd.n1129 avdd.t350 227.478
R12280 avdd.n1126 avdd.t364 227.478
R12281 avdd.t366 avdd.n1121 227.478
R12282 avdd.t377 avdd.n1118 227.478
R12283 avdd.n1115 avdd.t370 227.478
R12284 avdd.n1112 avdd.t241 227.478
R12285 avdd.t386 avdd.n1107 227.478
R12286 avdd.t250 avdd.n1104 227.478
R12287 avdd.n1649 avdd.t316 227.478
R12288 avdd.n1647 avdd.t293 227.478
R12289 avdd.n1645 avdd.t307 227.478
R12290 avdd.n1643 avdd.t287 227.478
R12291 avdd.n1641 avdd.t238 227.478
R12292 avdd.n1639 avdd.t280 227.478
R12293 avdd.n1637 avdd.t232 227.478
R12294 avdd.n1635 avdd.t373 227.478
R12295 avdd.n1633 avdd.t358 227.478
R12296 avdd.n1631 avdd.t355 227.478
R12297 avdd.n1629 avdd.t300 227.478
R12298 avdd.n1561 avdd.t362 227.478
R12299 avdd.t346 avdd.n1556 227.478
R12300 avdd.t352 avdd.n1553 227.478
R12301 avdd.n1550 avdd.t344 227.478
R12302 avdd.n1547 avdd.t270 227.478
R12303 avdd.t325 avdd.n1542 227.478
R12304 avdd.t266 avdd.n1539 227.478
R12305 avdd.n1536 avdd.t320 227.478
R12306 avdd.n1533 avdd.t302 227.478
R12307 avdd.t295 avdd.n1528 227.478
R12308 avdd.t264 avdd.n1525 227.478
R12309 avdd.n988 avdd.t223 227.345
R12310 avdd.t268 avdd.n1168 227.345
R12311 avdd.n1234 avdd.t273 227.345
R12312 avdd.t235 avdd.n1590 227.345
R12313 avdd.n22 avdd.t6 217.947
R12314 avdd.n1061 avdd.n991 211.953
R12315 avdd.n1307 avdd.n1237 211.953
R12316 avdd.n1799 avdd.t317 211.924
R12317 avdd.n1069 avdd.n1068 210.825
R12318 avdd.n1315 avdd.n1314 210.825
R12319 avdd.n1191 avdd.n1190 204.31
R12320 avdd.n1170 avdd.n1169 204.31
R12321 avdd.n1045 avdd.n1044 204.31
R12322 avdd.n1613 avdd.n1612 204.31
R12323 avdd.n1592 avdd.n1591 204.31
R12324 avdd.n1291 avdd.n1290 204.31
R12325 avdd.n1146 avdd.n1145 204.294
R12326 avdd.n1148 avdd.n1147 204.294
R12327 avdd.n1150 avdd.n1149 204.294
R12328 avdd.n1152 avdd.n1151 204.294
R12329 avdd.n1568 avdd.n1567 204.294
R12330 avdd.n1570 avdd.n1569 204.294
R12331 avdd.n1572 avdd.n1571 204.294
R12332 avdd.n1574 avdd.n1573 204.294
R12333 avdd.n1096 avdd.n1095 204.284
R12334 avdd.n1094 avdd.n1093 204.284
R12335 avdd.n1092 avdd.n1091 204.284
R12336 avdd.n1090 avdd.n1089 204.284
R12337 avdd.n1088 avdd.n1087 204.284
R12338 avdd.n1086 avdd.n1085 204.284
R12339 avdd.n1084 avdd.n1083 204.284
R12340 avdd.n1082 avdd.n1081 204.284
R12341 avdd.n1080 avdd.n1079 204.284
R12342 avdd.n1078 avdd.n1077 204.284
R12343 avdd.n1017 avdd.n1016 204.284
R12344 avdd.n1139 avdd.n1138 204.284
R12345 avdd.n1137 avdd.n1136 204.284
R12346 avdd.n1134 avdd.n1133 204.284
R12347 avdd.n1128 avdd.n1100 204.284
R12348 avdd.n1125 avdd.n1124 204.284
R12349 avdd.n1123 avdd.n1122 204.284
R12350 avdd.n1120 avdd.n1119 204.284
R12351 avdd.n1114 avdd.n1102 204.284
R12352 avdd.n1111 avdd.n1110 204.284
R12353 avdd.n1109 avdd.n1108 204.284
R12354 avdd.n1106 avdd.n1105 204.284
R12355 avdd.n1022 avdd.n1021 204.284
R12356 avdd.n1024 avdd.n1023 204.284
R12357 avdd.n1026 avdd.n1025 204.284
R12358 avdd.n1028 avdd.n1027 204.284
R12359 avdd.n1030 avdd.n1029 204.284
R12360 avdd.n1032 avdd.n1031 204.284
R12361 avdd.n1034 avdd.n1033 204.284
R12362 avdd.n1036 avdd.n1035 204.284
R12363 avdd.n1038 avdd.n1037 204.284
R12364 avdd.n1040 avdd.n1039 204.284
R12365 avdd.n1042 avdd.n1041 204.284
R12366 avdd.n1517 avdd.n1516 204.284
R12367 avdd.n1515 avdd.n1514 204.284
R12368 avdd.n1513 avdd.n1512 204.284
R12369 avdd.n1511 avdd.n1510 204.284
R12370 avdd.n1509 avdd.n1508 204.284
R12371 avdd.n1507 avdd.n1506 204.284
R12372 avdd.n1505 avdd.n1504 204.284
R12373 avdd.n1503 avdd.n1502 204.284
R12374 avdd.n1501 avdd.n1500 204.284
R12375 avdd.n1499 avdd.n1498 204.284
R12376 avdd.n1263 avdd.n1262 204.284
R12377 avdd.n1560 avdd.n1559 204.284
R12378 avdd.n1558 avdd.n1557 204.284
R12379 avdd.n1555 avdd.n1554 204.284
R12380 avdd.n1549 avdd.n1521 204.284
R12381 avdd.n1546 avdd.n1545 204.284
R12382 avdd.n1544 avdd.n1543 204.284
R12383 avdd.n1541 avdd.n1540 204.284
R12384 avdd.n1535 avdd.n1523 204.284
R12385 avdd.n1532 avdd.n1531 204.284
R12386 avdd.n1530 avdd.n1529 204.284
R12387 avdd.n1527 avdd.n1526 204.284
R12388 avdd.n1268 avdd.n1267 204.284
R12389 avdd.n1270 avdd.n1269 204.284
R12390 avdd.n1272 avdd.n1271 204.284
R12391 avdd.n1274 avdd.n1273 204.284
R12392 avdd.n1276 avdd.n1275 204.284
R12393 avdd.n1278 avdd.n1277 204.284
R12394 avdd.n1280 avdd.n1279 204.284
R12395 avdd.n1282 avdd.n1281 204.284
R12396 avdd.n1284 avdd.n1283 204.284
R12397 avdd.n1286 avdd.n1285 204.284
R12398 avdd.n1288 avdd.n1287 204.284
R12399 avdd.n1736 avdd.n1720 203.672
R12400 avdd.n1800 avdd.n1744 203.672
R12401 avdd.n1062 avdd.n1061 201.788
R12402 avdd.n1308 avdd.n1307 201.788
R12403 avdd.n1374 avdd.t542 201.107
R12404 avdd.n358 avdd.t159 197.562
R12405 avdd.n330 avdd.t151 197.562
R12406 avdd.n302 avdd.t492 197.562
R12407 avdd.n274 avdd.t149 197.562
R12408 avdd.n246 avdd.t422 197.562
R12409 avdd.n218 avdd.t99 197.562
R12410 avdd.n190 avdd.t103 197.562
R12411 avdd.n162 avdd.t123 197.562
R12412 avdd.n695 avdd.t588 197.562
R12413 avdd.n667 avdd.t91 197.562
R12414 avdd.n639 avdd.t173 197.562
R12415 avdd.n611 avdd.t142 197.562
R12416 avdd.n583 avdd.t34 197.562
R12417 avdd.n555 avdd.t619 197.562
R12418 avdd.n527 avdd.t36 197.562
R12419 avdd.n499 avdd.t586 197.562
R12420 avdd.n1796 avdd.n1725 196.142
R12421 avdd.t167 avdd.n996 195.042
R12422 avdd.t525 avdd.n1242 195.042
R12423 avdd.n109 avdd.t42 193.774
R12424 avdd.n446 avdd.t45 193.774
R12425 avdd.n1062 avdd.n1010 186.353
R12426 avdd.n1308 avdd.n1256 186.353
R12427 avdd.n21 avdd.n20 185
R12428 avdd.n22 avdd.n21 185
R12429 avdd.n6 avdd.n5 185
R12430 avdd.n12 avdd.n11 185
R12431 avdd.n10 avdd.n1 185
R12432 avdd.n25 avdd.n2 185
R12433 avdd.n24 avdd.n23 185
R12434 avdd.n23 avdd.n22 185
R12435 avdd.n357 avdd.n356 185
R12436 avdd.n358 avdd.n357 185
R12437 avdd.n41 avdd.n40 185
R12438 avdd.n352 avdd.n342 185
R12439 avdd.n351 avdd.n343 185
R12440 avdd.n38 avdd.n35 185
R12441 avdd.n361 avdd.n36 185
R12442 avdd.n329 avdd.n328 185
R12443 avdd.n330 avdd.n329 185
R12444 avdd.n49 avdd.n48 185
R12445 avdd.n324 avdd.n314 185
R12446 avdd.n323 avdd.n315 185
R12447 avdd.n46 avdd.n43 185
R12448 avdd.n333 avdd.n44 185
R12449 avdd.n301 avdd.n300 185
R12450 avdd.n302 avdd.n301 185
R12451 avdd.n57 avdd.n56 185
R12452 avdd.n296 avdd.n286 185
R12453 avdd.n295 avdd.n287 185
R12454 avdd.n54 avdd.n51 185
R12455 avdd.n305 avdd.n52 185
R12456 avdd.n273 avdd.n272 185
R12457 avdd.n274 avdd.n273 185
R12458 avdd.n65 avdd.n64 185
R12459 avdd.n268 avdd.n258 185
R12460 avdd.n267 avdd.n259 185
R12461 avdd.n62 avdd.n59 185
R12462 avdd.n277 avdd.n60 185
R12463 avdd.n245 avdd.n244 185
R12464 avdd.n246 avdd.n245 185
R12465 avdd.n73 avdd.n72 185
R12466 avdd.n240 avdd.n230 185
R12467 avdd.n239 avdd.n231 185
R12468 avdd.n70 avdd.n67 185
R12469 avdd.n249 avdd.n68 185
R12470 avdd.n217 avdd.n216 185
R12471 avdd.n218 avdd.n217 185
R12472 avdd.n81 avdd.n80 185
R12473 avdd.n212 avdd.n202 185
R12474 avdd.n211 avdd.n203 185
R12475 avdd.n78 avdd.n75 185
R12476 avdd.n221 avdd.n76 185
R12477 avdd.n189 avdd.n188 185
R12478 avdd.n190 avdd.n189 185
R12479 avdd.n89 avdd.n88 185
R12480 avdd.n184 avdd.n174 185
R12481 avdd.n183 avdd.n175 185
R12482 avdd.n86 avdd.n83 185
R12483 avdd.n193 avdd.n84 185
R12484 avdd.n161 avdd.n160 185
R12485 avdd.n162 avdd.n161 185
R12486 avdd.n97 avdd.n96 185
R12487 avdd.n156 avdd.n146 185
R12488 avdd.n155 avdd.n147 185
R12489 avdd.n94 avdd.n91 185
R12490 avdd.n165 avdd.n92 185
R12491 avdd.n110 avdd.n109 185
R12492 avdd.n105 avdd.n104 185
R12493 avdd.n104 avdd.n103 185
R12494 avdd.n126 avdd.n125 185
R12495 avdd.n127 avdd.n126 185
R12496 avdd.n106 avdd.n101 185
R12497 avdd.n128 avdd.n101 185
R12498 avdd.n130 avdd.n102 185
R12499 avdd.n130 avdd.n129 185
R12500 avdd.n131 avdd.n99 185
R12501 avdd.n132 avdd.n131 185
R12502 avdd.n137 avdd.n100 185
R12503 avdd.n133 avdd.n100 185
R12504 avdd.n136 avdd.n135 185
R12505 avdd.n135 avdd.n134 185
R12506 avdd.n694 avdd.n693 185
R12507 avdd.n695 avdd.n694 185
R12508 avdd.n378 avdd.n377 185
R12509 avdd.n689 avdd.n679 185
R12510 avdd.n688 avdd.n680 185
R12511 avdd.n375 avdd.n372 185
R12512 avdd.n698 avdd.n373 185
R12513 avdd.n666 avdd.n665 185
R12514 avdd.n667 avdd.n666 185
R12515 avdd.n386 avdd.n385 185
R12516 avdd.n661 avdd.n651 185
R12517 avdd.n660 avdd.n652 185
R12518 avdd.n383 avdd.n380 185
R12519 avdd.n670 avdd.n381 185
R12520 avdd.n638 avdd.n637 185
R12521 avdd.n639 avdd.n638 185
R12522 avdd.n394 avdd.n393 185
R12523 avdd.n633 avdd.n623 185
R12524 avdd.n632 avdd.n624 185
R12525 avdd.n391 avdd.n388 185
R12526 avdd.n642 avdd.n389 185
R12527 avdd.n610 avdd.n609 185
R12528 avdd.n611 avdd.n610 185
R12529 avdd.n402 avdd.n401 185
R12530 avdd.n605 avdd.n595 185
R12531 avdd.n604 avdd.n596 185
R12532 avdd.n399 avdd.n396 185
R12533 avdd.n614 avdd.n397 185
R12534 avdd.n582 avdd.n581 185
R12535 avdd.n583 avdd.n582 185
R12536 avdd.n410 avdd.n409 185
R12537 avdd.n577 avdd.n567 185
R12538 avdd.n576 avdd.n568 185
R12539 avdd.n407 avdd.n404 185
R12540 avdd.n586 avdd.n405 185
R12541 avdd.n554 avdd.n553 185
R12542 avdd.n555 avdd.n554 185
R12543 avdd.n418 avdd.n417 185
R12544 avdd.n549 avdd.n539 185
R12545 avdd.n548 avdd.n540 185
R12546 avdd.n415 avdd.n412 185
R12547 avdd.n558 avdd.n413 185
R12548 avdd.n526 avdd.n525 185
R12549 avdd.n527 avdd.n526 185
R12550 avdd.n426 avdd.n425 185
R12551 avdd.n521 avdd.n511 185
R12552 avdd.n520 avdd.n512 185
R12553 avdd.n423 avdd.n420 185
R12554 avdd.n530 avdd.n421 185
R12555 avdd.n498 avdd.n497 185
R12556 avdd.n499 avdd.n498 185
R12557 avdd.n434 avdd.n433 185
R12558 avdd.n493 avdd.n483 185
R12559 avdd.n492 avdd.n484 185
R12560 avdd.n431 avdd.n428 185
R12561 avdd.n502 avdd.n429 185
R12562 avdd.n447 avdd.n446 185
R12563 avdd.n442 avdd.n441 185
R12564 avdd.n441 avdd.n440 185
R12565 avdd.n463 avdd.n462 185
R12566 avdd.n464 avdd.n463 185
R12567 avdd.n443 avdd.n438 185
R12568 avdd.n465 avdd.n438 185
R12569 avdd.n467 avdd.n439 185
R12570 avdd.n467 avdd.n466 185
R12571 avdd.n468 avdd.n436 185
R12572 avdd.n469 avdd.n468 185
R12573 avdd.n474 avdd.n437 185
R12574 avdd.n470 avdd.n437 185
R12575 avdd.n473 avdd.n472 185
R12576 avdd.n472 avdd.n471 185
R12577 avdd.n714 avdd.n712 185
R12578 avdd.n715 avdd.n714 185
R12579 avdd.n718 avdd.n713 185
R12580 avdd.n1373 avdd.n1372 185
R12581 avdd.n1371 avdd.n1370 185
R12582 avdd.n1370 avdd.n1369 185
R12583 avdd.n1379 avdd.n1378 185
R12584 avdd.n1380 avdd.n1379 185
R12585 avdd.n1368 avdd.n1367 185
R12586 avdd.n1381 avdd.n1368 185
R12587 avdd.n1385 avdd.n1384 185
R12588 avdd.n1384 avdd.n1383 185
R12589 avdd.n1365 avdd.n1364 185
R12590 avdd.n1382 avdd.n1364 185
R12591 avdd.n1390 avdd.n1389 185
R12592 avdd.n1391 avdd.n1390 185
R12593 avdd.n1363 avdd.n1362 185
R12594 avdd.n1392 avdd.n1363 185
R12595 avdd.n1395 avdd.n1394 185
R12596 avdd.n1394 avdd.n1393 185
R12597 avdd.n1360 avdd.n1359 185
R12598 avdd.n1359 avdd.n1358 185
R12599 avdd.n1400 avdd.n1399 185
R12600 avdd.n1401 avdd.n1400 185
R12601 avdd.n1357 avdd.n1356 185
R12602 avdd.n1402 avdd.n1357 185
R12603 avdd.n1406 avdd.n1405 185
R12604 avdd.n1405 avdd.n1404 185
R12605 avdd.n1354 avdd.n1353 185
R12606 avdd.n1403 avdd.n1353 185
R12607 avdd.n1411 avdd.n1410 185
R12608 avdd.n1412 avdd.n1411 185
R12609 avdd.n1352 avdd.n1351 185
R12610 avdd.n1413 avdd.n1352 185
R12611 avdd.n1416 avdd.n1415 185
R12612 avdd.n1415 avdd.n1414 185
R12613 avdd.n1349 avdd.n1348 185
R12614 avdd.n1348 avdd.n1347 185
R12615 avdd.n1421 avdd.n1420 185
R12616 avdd.n1422 avdd.n1421 185
R12617 avdd.n1346 avdd.n1345 185
R12618 avdd.n1423 avdd.n1346 185
R12619 avdd.n1427 avdd.n1426 185
R12620 avdd.n1426 avdd.n1425 185
R12621 avdd.n1343 avdd.n1342 185
R12622 avdd.n1424 avdd.n1342 185
R12623 avdd.n1432 avdd.n1431 185
R12624 avdd.n1433 avdd.n1432 185
R12625 avdd.n1341 avdd.n1340 185
R12626 avdd.n1434 avdd.n1341 185
R12627 avdd.n1438 avdd.n1437 185
R12628 avdd.n1437 avdd.n1436 185
R12629 avdd.n1338 avdd.n1337 185
R12630 avdd.n1435 avdd.n1337 185
R12631 avdd.n1443 avdd.n1442 185
R12632 avdd.n1444 avdd.n1443 185
R12633 avdd.n1336 avdd.n1335 185
R12634 avdd.n1445 avdd.n1336 185
R12635 avdd.n1449 avdd.n1448 185
R12636 avdd.n1448 avdd.n1447 185
R12637 avdd.n1332 avdd.n1331 185
R12638 avdd.n1446 avdd.n1331 185
R12639 avdd.n1475 avdd.n1474 185
R12640 avdd.n1476 avdd.n1475 185
R12641 avdd.n1333 avdd.n1329 185
R12642 avdd.n1477 avdd.n1329 185
R12643 avdd.n1479 avdd.n1330 185
R12644 avdd.n1479 avdd.n1478 185
R12645 avdd.n1480 avdd.n1324 185
R12646 avdd.n1481 avdd.n1480 185
R12647 avdd.n1490 avdd.n1325 185
R12648 avdd.n1482 avdd.n1325 185
R12649 avdd.n1489 avdd.n1326 185
R12650 avdd.n1483 avdd.n1326 185
R12651 avdd.n1328 avdd.n1327 185
R12652 avdd.n959 avdd.n958 185
R12653 avdd.n958 avdd.n957 185
R12654 avdd.n738 avdd.n737 185
R12655 avdd.n956 avdd.n738 185
R12656 avdd.n954 avdd.n953 185
R12657 avdd.n955 avdd.n954 185
R12658 avdd.n948 avdd.n947 185
R12659 avdd.n947 avdd.n741 185
R12660 avdd.n946 avdd.n744 185
R12661 avdd.n946 avdd.n945 185
R12662 avdd.n747 avdd.n745 185
R12663 avdd.n944 avdd.n745 185
R12664 avdd.n942 avdd.n941 185
R12665 avdd.n943 avdd.n942 185
R12666 avdd.n940 avdd.n746 185
R12667 avdd.n758 avdd.n746 185
R12668 avdd.n759 avdd.n753 185
R12669 avdd.n760 avdd.n759 185
R12670 avdd.n934 avdd.n933 185
R12671 avdd.n933 avdd.n932 185
R12672 avdd.n757 avdd.n756 185
R12673 avdd.n931 avdd.n757 185
R12674 avdd.n929 avdd.n928 185
R12675 avdd.n930 avdd.n929 185
R12676 avdd.n923 avdd.n922 185
R12677 avdd.n922 avdd.n761 185
R12678 avdd.n921 avdd.n764 185
R12679 avdd.n921 avdd.n920 185
R12680 avdd.n767 avdd.n765 185
R12681 avdd.n919 avdd.n765 185
R12682 avdd.n917 avdd.n916 185
R12683 avdd.n918 avdd.n917 185
R12684 avdd.n915 avdd.n766 185
R12685 avdd.n778 avdd.n766 185
R12686 avdd.n779 avdd.n773 185
R12687 avdd.n780 avdd.n779 185
R12688 avdd.n909 avdd.n908 185
R12689 avdd.n908 avdd.n907 185
R12690 avdd.n777 avdd.n776 185
R12691 avdd.n906 avdd.n777 185
R12692 avdd.n904 avdd.n903 185
R12693 avdd.n905 avdd.n904 185
R12694 avdd.n898 avdd.n897 185
R12695 avdd.n897 avdd.n781 185
R12696 avdd.n896 avdd.n784 185
R12697 avdd.n896 avdd.n895 185
R12698 avdd.n787 avdd.n785 185
R12699 avdd.n894 avdd.n785 185
R12700 avdd.n892 avdd.n891 185
R12701 avdd.n893 avdd.n892 185
R12702 avdd.n890 avdd.n786 185
R12703 avdd.n798 avdd.n786 185
R12704 avdd.n799 avdd.n793 185
R12705 avdd.n800 avdd.n799 185
R12706 avdd.n884 avdd.n883 185
R12707 avdd.n883 avdd.n882 185
R12708 avdd.n797 avdd.n796 185
R12709 avdd.n881 avdd.n797 185
R12710 avdd.n879 avdd.n878 185
R12711 avdd.n880 avdd.n879 185
R12712 avdd.n873 avdd.n872 185
R12713 avdd.n872 avdd.n801 185
R12714 avdd.n871 avdd.n804 185
R12715 avdd.n871 avdd.n870 185
R12716 avdd.n807 avdd.n805 185
R12717 avdd.n869 avdd.n805 185
R12718 avdd.n867 avdd.n866 185
R12719 avdd.n868 avdd.n867 185
R12720 avdd.n865 avdd.n806 185
R12721 avdd.n818 avdd.n806 185
R12722 avdd.n819 avdd.n813 185
R12723 avdd.n820 avdd.n819 185
R12724 avdd.n859 avdd.n858 185
R12725 avdd.n858 avdd.n857 185
R12726 avdd.n817 avdd.n816 185
R12727 avdd.n856 avdd.n817 185
R12728 avdd.n854 avdd.n853 185
R12729 avdd.n855 avdd.n854 185
R12730 avdd.n848 avdd.n847 185
R12731 avdd.n847 avdd.n821 185
R12732 avdd.n846 avdd.n824 185
R12733 avdd.n846 avdd.n845 185
R12734 avdd.n827 avdd.n825 185
R12735 avdd.n844 avdd.n825 185
R12736 avdd.n842 avdd.n841 185
R12737 avdd.n843 avdd.n842 185
R12738 avdd.n840 avdd.n826 185
R12739 avdd.n966 avdd.n732 185
R12740 avdd.n965 avdd.n733 185
R12741 avdd.n739 avdd.n733 185
R12742 avdd.n964 avdd.n734 185
R12743 avdd.n740 avdd.n734 185
R12744 avdd.n1161 avdd.t240 180.231
R12745 avdd.n1201 avdd.t221 180.231
R12746 avdd.n1583 avdd.t234 180.231
R12747 avdd.n1623 avdd.t230 180.231
R12748 avdd.n1380 avdd.n1369 175.386
R12749 avdd.n1383 avdd.n1382 175.386
R12750 avdd.n1392 avdd.n1391 175.386
R12751 avdd.n1401 avdd.n1358 175.386
R12752 avdd.n1404 avdd.n1402 175.386
R12753 avdd.n1413 avdd.n1412 175.386
R12754 avdd.n1422 avdd.n1347 175.386
R12755 avdd.n1425 avdd.n1423 175.386
R12756 avdd.n1434 avdd.n1433 175.386
R12757 avdd.n1436 avdd.n1435 175.386
R12758 avdd.n1445 avdd.n1444 175.386
R12759 avdd.n1447 avdd.n1446 175.386
R12760 avdd.n1477 avdd.n1476 175.386
R12761 avdd.n1482 avdd.n1481 175.386
R12762 avdd.n1483 avdd.n1482 175.386
R12763 avdd.n740 avdd.n739 175.386
R12764 avdd.n956 avdd.n955 175.386
R12765 avdd.n945 avdd.n944 175.386
R12766 avdd.n760 avdd.n758 175.386
R12767 avdd.n931 avdd.n930 175.386
R12768 avdd.n920 avdd.n919 175.386
R12769 avdd.n780 avdd.n778 175.386
R12770 avdd.n906 avdd.n905 175.386
R12771 avdd.n895 avdd.n894 175.386
R12772 avdd.n800 avdd.n798 175.386
R12773 avdd.n881 avdd.n880 175.386
R12774 avdd.n870 avdd.n869 175.386
R12775 avdd.n820 avdd.n818 175.386
R12776 avdd.n856 avdd.n855 175.386
R12777 avdd.n845 avdd.n844 175.386
R12778 avdd.t590 avdd.n1483 169.905
R12779 avdd.n957 avdd.t121 169.905
R12780 avdd.t205 avdd.n741 169.905
R12781 avdd.n943 avdd.t16 169.905
R12782 avdd.n932 avdd.t105 169.905
R12783 avdd.t574 avdd.n761 169.905
R12784 avdd.n918 avdd.t8 169.905
R12785 avdd.n907 avdd.t572 169.905
R12786 avdd.t125 avdd.n781 169.905
R12787 avdd.n893 avdd.t494 169.905
R12788 avdd.n882 avdd.t622 169.905
R12789 avdd.t111 avdd.n801 169.905
R12790 avdd.n868 avdd.t218 169.905
R12791 avdd.n857 avdd.t536 169.905
R12792 avdd.t486 avdd.n821 169.905
R12793 avdd.n843 avdd.t500 169.905
R12794 avdd.t550 avdd.n1381 168.077
R12795 avdd.n1414 avdd.t544 168.077
R12796 avdd.t534 avdd.n1746 167.023
R12797 avdd.n1800 avdd.n1799 165.936
R12798 avdd.t113 avdd.n1445 162.596
R12799 avdd.t560 avdd.n1403 160.769
R12800 avdd.n1444 avdd.t540 160.769
R12801 avdd.n1802 avdd.n1801 155.859
R12802 avdd.n1806 avdd.n1805 155.859
R12803 avdd.n1195 avdd.t186 155.153
R12804 avdd.n1195 avdd.t179 155.153
R12805 avdd.n1617 avdd.t73 155.153
R12806 avdd.n1617 avdd.t65 155.153
R12807 avdd.n1465 avdd.n1452 154.113
R12808 avdd.n1464 avdd.n1453 154.113
R12809 avdd.n1463 avdd.n1454 154.113
R12810 avdd.n1462 avdd.n1455 154.113
R12811 avdd.n1461 avdd.n1456 154.113
R12812 avdd.n1460 avdd.n1457 154.113
R12813 avdd.n1459 avdd.n1458 154.113
R12814 avdd.n1469 avdd.n1468 154.042
R12815 avdd.t318 avdd.t534 153.764
R12816 avdd.n9 avdd.n8 153.571
R12817 avdd.n346 avdd.n345 153.571
R12818 avdd.n318 avdd.n317 153.571
R12819 avdd.n290 avdd.n289 153.571
R12820 avdd.n262 avdd.n261 153.571
R12821 avdd.n234 avdd.n233 153.571
R12822 avdd.n206 avdd.n205 153.571
R12823 avdd.n178 avdd.n177 153.571
R12824 avdd.n150 avdd.n149 153.571
R12825 avdd.n117 avdd.n116 153.571
R12826 avdd.n683 avdd.n682 153.571
R12827 avdd.n655 avdd.n654 153.571
R12828 avdd.n627 avdd.n626 153.571
R12829 avdd.n599 avdd.n598 153.571
R12830 avdd.n571 avdd.n570 153.571
R12831 avdd.n543 avdd.n542 153.571
R12832 avdd.n515 avdd.n514 153.571
R12833 avdd.n487 avdd.n486 153.571
R12834 avdd.n454 avdd.n453 153.571
R12835 avdd.t454 avdd.n1842 149.893
R12836 avdd.n1844 avdd.t474 149.893
R12837 avdd.t416 avdd.n1857 149.893
R12838 avdd.n1858 avdd.t140 149.893
R12839 avdd.n1393 avdd.t556 146.155
R12840 avdd.n1424 avdd.t548 146.155
R12841 avdd.n1478 avdd.t117 144.327
R12842 avdd.n1478 avdd.t119 140.673
R12843 avdd.n1393 avdd.t554 138.846
R12844 avdd.t568 avdd.n1424 138.846
R12845 avdd.n1845 avdd.n1839 125.742
R12846 avdd.n1837 avdd.n1820 125.742
R12847 avdd.n1403 avdd.t538 124.231
R12848 avdd.t523 avdd.t489 121.877
R12849 avdd.t515 avdd.t521 121.877
R12850 avdd.n127 avdd.n103 120.317
R12851 avdd.n129 avdd.n128 120.317
R12852 avdd.n133 avdd.n132 120.317
R12853 avdd.n134 avdd.n133 120.317
R12854 avdd.n466 avdd.n465 120.317
R12855 avdd.n470 avdd.n469 120.317
R12856 avdd.n471 avdd.n470 120.317
R12857 avdd.n464 avdd.n440 119.064
R12858 avdd.n22 avdd.t161 117.838
R12859 avdd.n1381 avdd.t558 116.924
R12860 avdd.n1414 avdd.t564 116.924
R12861 avdd.n1157 avdd.t49 116.782
R12862 avdd.n1157 avdd.t59 116.782
R12863 avdd.n1579 avdd.t22 116.782
R12864 avdd.n1579 avdd.t30 116.782
R12865 avdd.t161 avdd.t163 112.624
R12866 avdd.t468 avdd.t454 110.959
R12867 avdd.t484 avdd.t468 110.959
R12868 avdd.t464 avdd.t484 110.959
R12869 avdd.t480 avdd.t464 110.959
R12870 avdd.t476 avdd.t480 110.959
R12871 avdd.t458 avdd.t476 110.959
R12872 avdd.t472 avdd.t458 110.959
R12873 avdd.t470 avdd.t456 110.959
R12874 avdd.t466 avdd.t470 110.959
R12875 avdd.t482 avdd.t466 110.959
R12876 avdd.t462 avdd.t482 110.959
R12877 avdd.t478 avdd.t462 110.959
R12878 avdd.t460 avdd.t478 110.959
R12879 avdd.t474 avdd.t460 110.959
R12880 avdd.t415 avdd.t416 110.959
R12881 avdd.t304 avdd.t415 110.959
R12882 avdd.t94 avdd.t304 110.959
R12883 avdd.t93 avdd.t94 110.959
R12884 avdd.t243 avdd.t93 110.959
R12885 avdd.t579 avdd.t243 110.959
R12886 avdd.t578 avdd.t579 110.959
R12887 avdd.t333 avdd.t578 110.959
R12888 avdd.t497 avdd.t333 110.959
R12889 avdd.t496 avdd.t497 110.959
R12890 avdd.t275 avdd.t496 110.959
R12891 avdd.t444 avdd.t275 110.959
R12892 avdd.t445 avdd.t444 110.959
R12893 avdd.t375 avdd.t445 110.959
R12894 avdd.t138 avdd.t375 110.959
R12895 avdd.t137 avdd.t138 110.959
R12896 avdd.t262 avdd.t137 110.959
R12897 avdd.t176 avdd.t262 110.959
R12898 avdd.t175 avdd.t176 110.959
R12899 avdd.t393 avdd.t175 110.959
R12900 avdd.t508 avdd.t393 110.959
R12901 avdd.t507 avdd.t508 110.959
R12902 avdd.t381 avdd.t507 110.959
R12903 avdd.t4 avdd.t381 110.959
R12904 avdd.t5 avdd.t4 110.959
R12905 avdd.t368 avdd.t5 110.959
R12906 avdd.t451 avdd.t368 110.959
R12907 avdd.t450 avdd.t451 110.959
R12908 avdd.t379 avdd.t450 110.959
R12909 avdd.t157 avdd.t379 110.959
R12910 avdd.t158 avdd.t157 110.959
R12911 avdd.t297 avdd.t158 110.959
R12912 avdd.t109 avdd.t297 110.959
R12913 avdd.t110 avdd.t109 110.959
R12914 avdd.t391 avdd.t110 110.959
R12915 avdd.t171 avdd.t391 110.959
R12916 avdd.t172 avdd.t171 110.959
R12917 avdd.t395 avdd.t172 110.959
R12918 avdd.t627 avdd.t395 110.959
R12919 avdd.t628 avdd.t627 110.959
R12920 avdd.t360 avdd.t628 110.959
R12921 avdd.t414 avdd.t360 110.959
R12922 avdd.t413 avdd.t414 110.959
R12923 avdd.t248 avdd.t413 110.959
R12924 avdd.t139 avdd.t248 110.959
R12925 avdd.t140 avdd.t139 110.959
R12926 avdd.n358 avdd.t653 106.817
R12927 avdd.n330 avdd.t436 106.817
R12928 avdd.n302 avdd.t12 106.817
R12929 avdd.n274 avdd.t511 106.817
R12930 avdd.n246 avdd.t440 106.817
R12931 avdd.n218 avdd.t215 106.817
R12932 avdd.n190 avdd.t410 106.817
R12933 avdd.n162 avdd.t502 106.817
R12934 avdd.n695 avdd.t656 106.817
R12935 avdd.n667 avdd.t0 106.817
R12936 avdd.n639 avdd.t153 106.817
R12937 avdd.n611 avdd.t144 106.817
R12938 avdd.n583 avdd.t398 106.817
R12939 avdd.n555 avdd.t593 106.817
R12940 avdd.n527 avdd.t625 106.817
R12941 avdd.n499 avdd.t40 106.817
R12942 avdd.t209 avdd.n127 106.531
R12943 avdd.t129 avdd.n464 106.531
R12944 avdd.n1198 avdd.n1010 105.412
R12945 avdd.n1620 avdd.n1256 105.412
R12946 avdd.n1382 avdd.t552 102.308
R12947 avdd.t546 avdd.n1422 102.308
R12948 avdd.t653 avdd.t10 102.091
R12949 avdd.t436 avdd.t438 102.091
R12950 avdd.t12 avdd.t14 102.091
R12951 avdd.t511 avdd.t147 102.091
R12952 avdd.t440 avdd.t442 102.091
R12953 avdd.t215 avdd.t107 102.091
R12954 avdd.t410 avdd.t207 102.091
R12955 avdd.t502 avdd.t101 102.091
R12956 avdd.t656 avdd.t498 102.091
R12957 avdd.t0 avdd.t2 102.091
R12958 avdd.t153 avdd.t155 102.091
R12959 avdd.t144 avdd.t127 102.091
R12960 avdd.t398 avdd.t396 102.091
R12961 avdd.t593 avdd.t576 102.091
R12962 avdd.t625 avdd.t452 102.091
R12963 avdd.t40 avdd.t38 102.091
R12964 avdd.t42 avdd.n103 101.564
R12965 avdd.t45 avdd.n440 101.564
R12966 avdd.n1004 avdd.n1003 99.0123
R12967 avdd.n1009 avdd.n1008 99.0123
R12968 avdd.n1250 avdd.n1249 99.0123
R12969 avdd.n1255 avdd.n1254 99.0123
R12970 avdd.n134 avdd.t135 97.7578
R12971 avdd.n471 avdd.t570 97.7578
R12972 avdd.n1446 avdd.t115 96.8274
R12973 avdd.t529 avdd.n1728 96.5971
R12974 avdd.n1402 avdd.t566 95.0005
R12975 avdd.n1436 avdd.t562 95.0005
R12976 avdd.n1204 avdd.n1203 94.1181
R12977 avdd.n1164 avdd.n1163 94.1181
R12978 avdd.n1626 avdd.n1625 94.1181
R12979 avdd.n1586 avdd.n1585 94.1181
R12980 avdd.n1053 avdd.n1048 91.1064
R12981 avdd.n1299 avdd.n1294 91.1064
R12982 avdd.t430 avdd.t529 88.8801
R12983 avdd.n5 avdd.n3 86.068
R12984 avdd.n10 avdd.n4 86.068
R12985 avdd.n11 avdd.n3 86.068
R12986 avdd.n4 avdd.n2 86.068
R12987 avdd.n40 avdd.n37 86.068
R12988 avdd.n343 avdd.n39 86.068
R12989 avdd.n359 avdd.n36 86.068
R12990 avdd.n342 avdd.n37 86.068
R12991 avdd.n39 avdd.n38 86.068
R12992 avdd.n48 avdd.n45 86.068
R12993 avdd.n315 avdd.n47 86.068
R12994 avdd.n331 avdd.n44 86.068
R12995 avdd.n314 avdd.n45 86.068
R12996 avdd.n47 avdd.n46 86.068
R12997 avdd.n56 avdd.n53 86.068
R12998 avdd.n287 avdd.n55 86.068
R12999 avdd.n303 avdd.n52 86.068
R13000 avdd.n286 avdd.n53 86.068
R13001 avdd.n55 avdd.n54 86.068
R13002 avdd.n64 avdd.n61 86.068
R13003 avdd.n259 avdd.n63 86.068
R13004 avdd.n275 avdd.n60 86.068
R13005 avdd.n258 avdd.n61 86.068
R13006 avdd.n63 avdd.n62 86.068
R13007 avdd.n72 avdd.n69 86.068
R13008 avdd.n231 avdd.n71 86.068
R13009 avdd.n247 avdd.n68 86.068
R13010 avdd.n230 avdd.n69 86.068
R13011 avdd.n71 avdd.n70 86.068
R13012 avdd.n80 avdd.n77 86.068
R13013 avdd.n203 avdd.n79 86.068
R13014 avdd.n219 avdd.n76 86.068
R13015 avdd.n202 avdd.n77 86.068
R13016 avdd.n79 avdd.n78 86.068
R13017 avdd.n88 avdd.n85 86.068
R13018 avdd.n175 avdd.n87 86.068
R13019 avdd.n191 avdd.n84 86.068
R13020 avdd.n174 avdd.n85 86.068
R13021 avdd.n87 avdd.n86 86.068
R13022 avdd.n96 avdd.n93 86.068
R13023 avdd.n147 avdd.n95 86.068
R13024 avdd.n163 avdd.n92 86.068
R13025 avdd.n146 avdd.n93 86.068
R13026 avdd.n95 avdd.n94 86.068
R13027 avdd.n377 avdd.n374 86.068
R13028 avdd.n680 avdd.n376 86.068
R13029 avdd.n696 avdd.n373 86.068
R13030 avdd.n679 avdd.n374 86.068
R13031 avdd.n376 avdd.n375 86.068
R13032 avdd.n385 avdd.n382 86.068
R13033 avdd.n652 avdd.n384 86.068
R13034 avdd.n668 avdd.n381 86.068
R13035 avdd.n651 avdd.n382 86.068
R13036 avdd.n384 avdd.n383 86.068
R13037 avdd.n393 avdd.n390 86.068
R13038 avdd.n624 avdd.n392 86.068
R13039 avdd.n640 avdd.n389 86.068
R13040 avdd.n623 avdd.n390 86.068
R13041 avdd.n392 avdd.n391 86.068
R13042 avdd.n401 avdd.n398 86.068
R13043 avdd.n596 avdd.n400 86.068
R13044 avdd.n612 avdd.n397 86.068
R13045 avdd.n595 avdd.n398 86.068
R13046 avdd.n400 avdd.n399 86.068
R13047 avdd.n409 avdd.n406 86.068
R13048 avdd.n568 avdd.n408 86.068
R13049 avdd.n584 avdd.n405 86.068
R13050 avdd.n567 avdd.n406 86.068
R13051 avdd.n408 avdd.n407 86.068
R13052 avdd.n417 avdd.n414 86.068
R13053 avdd.n540 avdd.n416 86.068
R13054 avdd.n556 avdd.n413 86.068
R13055 avdd.n539 avdd.n414 86.068
R13056 avdd.n416 avdd.n415 86.068
R13057 avdd.n425 avdd.n422 86.068
R13058 avdd.n512 avdd.n424 86.068
R13059 avdd.n528 avdd.n421 86.068
R13060 avdd.n511 avdd.n422 86.068
R13061 avdd.n424 avdd.n423 86.068
R13062 avdd.n433 avdd.n430 86.068
R13063 avdd.n484 avdd.n432 86.068
R13064 avdd.n500 avdd.n429 86.068
R13065 avdd.n483 avdd.n430 86.068
R13066 avdd.n432 avdd.n431 86.068
R13067 avdd.n716 avdd.n713 86.068
R13068 avdd.n1484 avdd.t590 82.3568
R13069 avdd.n833 avdd.t500 82.3568
R13070 avdd.t566 avdd.n1401 80.3851
R13071 avdd.t562 avdd.n1434 80.3851
R13072 avdd.n1476 avdd.t115 78.5582
R13073 avdd.t515 avdd.t434 73.4459
R13074 avdd.n1391 avdd.t552 73.0774
R13075 avdd.n1423 avdd.t546 73.0774
R13076 avdd.n129 avdd.t213 72.6918
R13077 avdd.n466 avdd.t133 72.6918
R13078 avdd.n1003 avdd.n991 71.5299
R13079 avdd.n1010 avdd.n1009 71.5299
R13080 avdd.n1249 avdd.n1237 71.5299
R13081 avdd.n1256 avdd.n1255 71.5299
R13082 avdd.t517 avdd.n1749 69.9865
R13083 avdd.n1374 avdd.n1373 68.6629
R13084 avdd.n1484 avdd.n1328 68.6629
R13085 avdd.n833 avdd.n826 68.6629
R13086 avdd.n1755 avdd.t506 59.3422
R13087 avdd.t558 avdd.n1380 58.462
R13088 avdd.t564 avdd.n1413 58.462
R13089 avdd.t225 avdd.t523 58.0117
R13090 avdd.n1843 avdd.t472 55.4795
R13091 avdd.t456 avdd.n1843 55.4795
R13092 avdd.n1835 avdd.t475 54.6604
R13093 avdd.n1818 avdd.t455 54.6604
R13094 avdd.n1738 avdd.t530 53.8832
R13095 avdd.n1732 avdd.t518 53.8832
R13096 avdd.n1731 avdd.t535 53.8832
R13097 avdd.t542 avdd.n1369 51.1543
R13098 avdd.n1412 avdd.t538 51.1543
R13099 avdd.n1716 avdd.n1715 50.4475
R13100 avdd.n1778 avdd.t329 49.5908
R13101 avdd.n1762 avdd.t329 49.5908
R13102 avdd.n22 avdd.n3 49.4675
R13103 avdd.n22 avdd.n4 49.4675
R13104 avdd.n358 avdd.n37 49.4675
R13105 avdd.n358 avdd.n39 49.4675
R13106 avdd.n359 avdd.n358 49.4675
R13107 avdd.n330 avdd.n45 49.4675
R13108 avdd.n330 avdd.n47 49.4675
R13109 avdd.n331 avdd.n330 49.4675
R13110 avdd.n302 avdd.n53 49.4675
R13111 avdd.n302 avdd.n55 49.4675
R13112 avdd.n303 avdd.n302 49.4675
R13113 avdd.n274 avdd.n61 49.4675
R13114 avdd.n274 avdd.n63 49.4675
R13115 avdd.n275 avdd.n274 49.4675
R13116 avdd.n246 avdd.n69 49.4675
R13117 avdd.n246 avdd.n71 49.4675
R13118 avdd.n247 avdd.n246 49.4675
R13119 avdd.n218 avdd.n77 49.4675
R13120 avdd.n218 avdd.n79 49.4675
R13121 avdd.n219 avdd.n218 49.4675
R13122 avdd.n190 avdd.n85 49.4675
R13123 avdd.n190 avdd.n87 49.4675
R13124 avdd.n191 avdd.n190 49.4675
R13125 avdd.n162 avdd.n93 49.4675
R13126 avdd.n162 avdd.n95 49.4675
R13127 avdd.n163 avdd.n162 49.4675
R13128 avdd.n695 avdd.n374 49.4675
R13129 avdd.n695 avdd.n376 49.4675
R13130 avdd.n696 avdd.n695 49.4675
R13131 avdd.n667 avdd.n382 49.4675
R13132 avdd.n667 avdd.n384 49.4675
R13133 avdd.n668 avdd.n667 49.4675
R13134 avdd.n639 avdd.n390 49.4675
R13135 avdd.n639 avdd.n392 49.4675
R13136 avdd.n640 avdd.n639 49.4675
R13137 avdd.n611 avdd.n398 49.4675
R13138 avdd.n611 avdd.n400 49.4675
R13139 avdd.n612 avdd.n611 49.4675
R13140 avdd.n583 avdd.n406 49.4675
R13141 avdd.n583 avdd.n408 49.4675
R13142 avdd.n584 avdd.n583 49.4675
R13143 avdd.n555 avdd.n414 49.4675
R13144 avdd.n555 avdd.n416 49.4675
R13145 avdd.n556 avdd.n555 49.4675
R13146 avdd.n527 avdd.n422 49.4675
R13147 avdd.n527 avdd.n424 49.4675
R13148 avdd.n528 avdd.n527 49.4675
R13149 avdd.n499 avdd.n430 49.4675
R13150 avdd.n499 avdd.n432 49.4675
R13151 avdd.n500 avdd.n499 49.4675
R13152 avdd.n716 avdd.n715 49.4675
R13153 avdd.n1834 avdd.n1833 49.1214
R13154 avdd.n1832 avdd.n1831 49.1214
R13155 avdd.n1830 avdd.n1829 49.1214
R13156 avdd.n1828 avdd.n1827 49.1214
R13157 avdd.n1826 avdd.n1825 49.1214
R13158 avdd.n1824 avdd.n1823 49.1214
R13159 avdd.n1822 avdd.n1821 49.1214
R13160 avdd.t489 avdd.t434 48.4319
R13161 avdd.n1740 avdd.n1739 48.3442
R13162 avdd.n1742 avdd.n1741 48.3442
R13163 avdd.n1767 avdd.n1766 48.2034
R13164 avdd.n1769 avdd.n1768 48.2034
R13165 avdd.n1775 avdd.n1774 48.2034
R13166 avdd.n1782 avdd.n1781 48.2034
R13167 avdd.n1784 avdd.n1783 48.2034
R13168 avdd.n1786 avdd.n1785 48.2034
R13169 avdd.n1788 avdd.n1787 48.2034
R13170 avdd.n1764 avdd.t260 48.0365
R13171 avdd.n1789 avdd.t226 48.0365
R13172 avdd.n132 avdd.t213 47.6258
R13173 avdd.n469 avdd.t133 47.6258
R13174 avdd.t505 avdd.t491 47.3674
R13175 avdd.t491 avdd.t228 47.3674
R13176 avdd.t228 avdd.t488 47.3674
R13177 avdd.t348 avdd.t488 47.3674
R13178 avdd.t338 avdd.t533 47.3674
R13179 avdd.t531 avdd.t338 47.3674
R13180 avdd.t506 avdd.t531 47.3674
R13181 avdd.n1205 avdd.n1204 44.8005
R13182 avdd.n1165 avdd.n1164 44.8005
R13183 avdd.n1627 avdd.n1626 44.8005
R13184 avdd.n1587 avdd.n1586 44.8005
R13185 avdd.n1054 avdd.n1049 43.2946
R13186 avdd.n1300 avdd.n1295 43.2946
R13187 avdd.n1728 avdd.t95 42.8436
R13188 avdd.n1771 avdd.n1770 42.4975
R13189 avdd.n1773 avdd.n1763 42.4505
R13190 avdd.n1795 avdd.t517 41.247
R13191 avdd.n1749 avdd.t225 38.5859
R13192 avdd.n1008 avdd.n1007 37.0005
R13193 avdd.n1005 avdd.n1004 37.0005
R13194 avdd.n1254 avdd.n1253 37.0005
R13195 avdd.n1251 avdd.n1250 37.0005
R13196 avdd.t554 avdd.n1392 36.539
R13197 avdd.n1425 avdd.t568 36.539
R13198 avdd.n1694 avdd.n1693 36.4934
R13199 avdd.n20 avdd.n6 36.1417
R13200 avdd.n12 avdd.n6 36.1417
R13201 avdd.n12 avdd.n1 36.1417
R13202 avdd.n25 avdd.n1 36.1417
R13203 avdd.n25 avdd.n24 36.1417
R13204 avdd.n356 avdd.n41 36.1417
R13205 avdd.n352 avdd.n41 36.1417
R13206 avdd.n352 avdd.n351 36.1417
R13207 avdd.n351 avdd.n35 36.1417
R13208 avdd.n361 avdd.n35 36.1417
R13209 avdd.n361 avdd.n360 36.1417
R13210 avdd.n328 avdd.n49 36.1417
R13211 avdd.n324 avdd.n49 36.1417
R13212 avdd.n324 avdd.n323 36.1417
R13213 avdd.n323 avdd.n43 36.1417
R13214 avdd.n333 avdd.n43 36.1417
R13215 avdd.n333 avdd.n332 36.1417
R13216 avdd.n300 avdd.n57 36.1417
R13217 avdd.n296 avdd.n57 36.1417
R13218 avdd.n296 avdd.n295 36.1417
R13219 avdd.n295 avdd.n51 36.1417
R13220 avdd.n305 avdd.n51 36.1417
R13221 avdd.n305 avdd.n304 36.1417
R13222 avdd.n272 avdd.n65 36.1417
R13223 avdd.n268 avdd.n65 36.1417
R13224 avdd.n268 avdd.n267 36.1417
R13225 avdd.n267 avdd.n59 36.1417
R13226 avdd.n277 avdd.n59 36.1417
R13227 avdd.n277 avdd.n276 36.1417
R13228 avdd.n244 avdd.n73 36.1417
R13229 avdd.n240 avdd.n73 36.1417
R13230 avdd.n240 avdd.n239 36.1417
R13231 avdd.n239 avdd.n67 36.1417
R13232 avdd.n249 avdd.n67 36.1417
R13233 avdd.n249 avdd.n248 36.1417
R13234 avdd.n216 avdd.n81 36.1417
R13235 avdd.n212 avdd.n81 36.1417
R13236 avdd.n212 avdd.n211 36.1417
R13237 avdd.n211 avdd.n75 36.1417
R13238 avdd.n221 avdd.n75 36.1417
R13239 avdd.n221 avdd.n220 36.1417
R13240 avdd.n188 avdd.n89 36.1417
R13241 avdd.n184 avdd.n89 36.1417
R13242 avdd.n184 avdd.n183 36.1417
R13243 avdd.n183 avdd.n83 36.1417
R13244 avdd.n193 avdd.n83 36.1417
R13245 avdd.n193 avdd.n192 36.1417
R13246 avdd.n160 avdd.n97 36.1417
R13247 avdd.n156 avdd.n97 36.1417
R13248 avdd.n156 avdd.n155 36.1417
R13249 avdd.n155 avdd.n91 36.1417
R13250 avdd.n165 avdd.n91 36.1417
R13251 avdd.n165 avdd.n164 36.1417
R13252 avdd.n110 avdd.n105 36.1417
R13253 avdd.n125 avdd.n105 36.1417
R13254 avdd.n125 avdd.n106 36.1417
R13255 avdd.n106 avdd.n102 36.1417
R13256 avdd.n102 avdd.n99 36.1417
R13257 avdd.n137 avdd.n99 36.1417
R13258 avdd.n137 avdd.n136 36.1417
R13259 avdd.n693 avdd.n378 36.1417
R13260 avdd.n689 avdd.n378 36.1417
R13261 avdd.n689 avdd.n688 36.1417
R13262 avdd.n688 avdd.n372 36.1417
R13263 avdd.n698 avdd.n372 36.1417
R13264 avdd.n698 avdd.n697 36.1417
R13265 avdd.n665 avdd.n386 36.1417
R13266 avdd.n661 avdd.n386 36.1417
R13267 avdd.n661 avdd.n660 36.1417
R13268 avdd.n660 avdd.n380 36.1417
R13269 avdd.n670 avdd.n380 36.1417
R13270 avdd.n670 avdd.n669 36.1417
R13271 avdd.n637 avdd.n394 36.1417
R13272 avdd.n633 avdd.n394 36.1417
R13273 avdd.n633 avdd.n632 36.1417
R13274 avdd.n632 avdd.n388 36.1417
R13275 avdd.n642 avdd.n388 36.1417
R13276 avdd.n642 avdd.n641 36.1417
R13277 avdd.n609 avdd.n402 36.1417
R13278 avdd.n605 avdd.n402 36.1417
R13279 avdd.n605 avdd.n604 36.1417
R13280 avdd.n604 avdd.n396 36.1417
R13281 avdd.n614 avdd.n396 36.1417
R13282 avdd.n614 avdd.n613 36.1417
R13283 avdd.n581 avdd.n410 36.1417
R13284 avdd.n577 avdd.n410 36.1417
R13285 avdd.n577 avdd.n576 36.1417
R13286 avdd.n576 avdd.n404 36.1417
R13287 avdd.n586 avdd.n404 36.1417
R13288 avdd.n586 avdd.n585 36.1417
R13289 avdd.n553 avdd.n418 36.1417
R13290 avdd.n549 avdd.n418 36.1417
R13291 avdd.n549 avdd.n548 36.1417
R13292 avdd.n548 avdd.n412 36.1417
R13293 avdd.n558 avdd.n412 36.1417
R13294 avdd.n558 avdd.n557 36.1417
R13295 avdd.n525 avdd.n426 36.1417
R13296 avdd.n521 avdd.n426 36.1417
R13297 avdd.n521 avdd.n520 36.1417
R13298 avdd.n520 avdd.n420 36.1417
R13299 avdd.n530 avdd.n420 36.1417
R13300 avdd.n530 avdd.n529 36.1417
R13301 avdd.n497 avdd.n434 36.1417
R13302 avdd.n493 avdd.n434 36.1417
R13303 avdd.n493 avdd.n492 36.1417
R13304 avdd.n492 avdd.n428 36.1417
R13305 avdd.n502 avdd.n428 36.1417
R13306 avdd.n502 avdd.n501 36.1417
R13307 avdd.n447 avdd.n442 36.1417
R13308 avdd.n462 avdd.n443 36.1417
R13309 avdd.n443 avdd.n439 36.1417
R13310 avdd.n439 avdd.n436 36.1417
R13311 avdd.n474 avdd.n436 36.1417
R13312 avdd.n474 avdd.n473 36.1417
R13313 avdd.n718 avdd.n712 36.1417
R13314 avdd.n718 avdd.n717 36.1417
R13315 avdd.n1372 avdd.n1371 36.1417
R13316 avdd.n1378 avdd.n1371 36.1417
R13317 avdd.n1378 avdd.n1367 36.1417
R13318 avdd.n1385 avdd.n1367 36.1417
R13319 avdd.n1385 avdd.n1365 36.1417
R13320 avdd.n1389 avdd.n1365 36.1417
R13321 avdd.n1389 avdd.n1362 36.1417
R13322 avdd.n1395 avdd.n1362 36.1417
R13323 avdd.n1395 avdd.n1360 36.1417
R13324 avdd.n1399 avdd.n1360 36.1417
R13325 avdd.n1399 avdd.n1356 36.1417
R13326 avdd.n1406 avdd.n1356 36.1417
R13327 avdd.n1406 avdd.n1354 36.1417
R13328 avdd.n1410 avdd.n1354 36.1417
R13329 avdd.n1410 avdd.n1351 36.1417
R13330 avdd.n1416 avdd.n1351 36.1417
R13331 avdd.n1416 avdd.n1349 36.1417
R13332 avdd.n1420 avdd.n1349 36.1417
R13333 avdd.n1420 avdd.n1345 36.1417
R13334 avdd.n1427 avdd.n1345 36.1417
R13335 avdd.n1427 avdd.n1343 36.1417
R13336 avdd.n1431 avdd.n1343 36.1417
R13337 avdd.n1431 avdd.n1340 36.1417
R13338 avdd.n1438 avdd.n1340 36.1417
R13339 avdd.n1438 avdd.n1338 36.1417
R13340 avdd.n1442 avdd.n1338 36.1417
R13341 avdd.n1442 avdd.n1335 36.1417
R13342 avdd.n1449 avdd.n1335 36.1417
R13343 avdd.n1449 avdd.n1332 36.1417
R13344 avdd.n1474 avdd.n1332 36.1417
R13345 avdd.n1474 avdd.n1333 36.1417
R13346 avdd.n1333 avdd.n1330 36.1417
R13347 avdd.n1330 avdd.n1324 36.1417
R13348 avdd.n1490 avdd.n1324 36.1417
R13349 avdd.n1490 avdd.n1489 36.1417
R13350 avdd.n1489 avdd.n1327 36.1417
R13351 avdd.n1485 avdd.n1327 36.1417
R13352 avdd.n841 avdd.n840 36.1417
R13353 avdd.n840 avdd.n834 36.1417
R13354 avdd.n848 avdd.n824 36.1417
R13355 avdd.n827 avdd.n824 36.1417
R13356 avdd.n859 avdd.n816 36.1417
R13357 avdd.n853 avdd.n816 36.1417
R13358 avdd.n866 avdd.n865 36.1417
R13359 avdd.n865 avdd.n813 36.1417
R13360 avdd.n873 avdd.n804 36.1417
R13361 avdd.n807 avdd.n804 36.1417
R13362 avdd.n884 avdd.n796 36.1417
R13363 avdd.n878 avdd.n796 36.1417
R13364 avdd.n891 avdd.n890 36.1417
R13365 avdd.n890 avdd.n793 36.1417
R13366 avdd.n898 avdd.n784 36.1417
R13367 avdd.n787 avdd.n784 36.1417
R13368 avdd.n909 avdd.n776 36.1417
R13369 avdd.n903 avdd.n776 36.1417
R13370 avdd.n916 avdd.n915 36.1417
R13371 avdd.n915 avdd.n773 36.1417
R13372 avdd.n923 avdd.n764 36.1417
R13373 avdd.n767 avdd.n764 36.1417
R13374 avdd.n934 avdd.n756 36.1417
R13375 avdd.n928 avdd.n756 36.1417
R13376 avdd.n941 avdd.n940 36.1417
R13377 avdd.n940 avdd.n753 36.1417
R13378 avdd.n948 avdd.n744 36.1417
R13379 avdd.n747 avdd.n744 36.1417
R13380 avdd.n959 avdd.n737 36.1417
R13381 avdd.n953 avdd.n737 36.1417
R13382 avdd.n966 avdd.n965 36.1417
R13383 avdd.n965 avdd.n964 36.1417
R13384 avdd.n462 avdd.n442 35.7652
R13385 avdd.n1481 avdd.t119 34.712
R13386 avdd.t521 avdd.t430 32.9977
R13387 avdd.n1736 avdd.n1724 31.624
R13388 avdd.n1747 avdd.n1744 31.624
R13389 avdd.n1812 avdd.n1719 31.624
R13390 avdd.n1154 avdd.n1076 31.2476
R13391 avdd.n1074 avdd.n1073 31.2476
R13392 avdd.n1576 avdd.n1322 31.2476
R13393 avdd.n1320 avdd.n1319 31.2476
R13394 avdd.n1693 avdd.n1666 31.2285
R13395 avdd.t117 avdd.n1477 31.0582
R13396 avdd.n1163 avdd.n1162 30.8338
R13397 avdd.n1162 avdd.n1161 30.8338
R13398 avdd.n1203 avdd.n1202 30.8338
R13399 avdd.n1202 avdd.n1201 30.8338
R13400 avdd.n1076 avdd.n1072 30.8338
R13401 avdd.n1074 avdd.n1071 30.8338
R13402 avdd.n1585 avdd.n1584 30.8338
R13403 avdd.n1584 avdd.n1583 30.8338
R13404 avdd.n1625 avdd.n1624 30.8338
R13405 avdd.n1624 avdd.n1623 30.8338
R13406 avdd.n1322 avdd.n1318 30.8338
R13407 avdd.n1320 avdd.n1317 30.8338
R13408 avdd.n1675 avdd.n1673 30.3029
R13409 avdd.t556 avdd.n1358 29.2313
R13410 avdd.n1433 avdd.t548 29.2313
R13411 avdd.n1699 avdd.n1694 27.9872
R13412 avdd.n1095 avdd.t187 27.6955
R13413 avdd.n1095 avdd.t595 27.6955
R13414 avdd.n1093 avdd.t190 27.6955
R13415 avdd.n1093 avdd.t597 27.6955
R13416 avdd.n1091 avdd.t188 27.6955
R13417 avdd.n1091 avdd.t596 27.6955
R13418 avdd.n1089 avdd.t196 27.6955
R13419 avdd.n1089 avdd.t606 27.6955
R13420 avdd.n1087 avdd.t613 27.6955
R13421 avdd.n1087 avdd.t191 27.6955
R13422 avdd.n1085 avdd.t614 27.6955
R13423 avdd.n1085 avdd.t192 27.6955
R13424 avdd.n1083 avdd.t617 27.6955
R13425 avdd.n1083 avdd.t194 27.6955
R13426 avdd.n1081 avdd.t615 27.6955
R13427 avdd.n1081 avdd.t193 27.6955
R13428 avdd.n1079 avdd.t598 27.6955
R13429 avdd.n1079 avdd.t197 27.6955
R13430 avdd.n1077 avdd.t618 27.6955
R13431 avdd.n1077 avdd.t195 27.6955
R13432 avdd.n1016 avdd.t599 27.6955
R13433 avdd.n1016 avdd.t199 27.6955
R13434 avdd.n1190 avdd.t604 27.6955
R13435 avdd.n1190 avdd.t180 27.6955
R13436 avdd.t277 avdd.n1139 27.6955
R13437 avdd.n1139 avdd.t198 27.6955
R13438 avdd.n1136 avdd.t284 27.6955
R13439 avdd.n1136 avdd.t201 27.6955
R13440 avdd.n1133 avdd.t282 27.6955
R13441 avdd.n1133 avdd.t200 27.6955
R13442 avdd.t350 avdd.n1128 27.6955
R13443 avdd.n1128 avdd.t183 27.6955
R13444 avdd.t364 avdd.n1125 27.6955
R13445 avdd.n1125 avdd.t600 27.6955
R13446 avdd.n1122 avdd.t366 27.6955
R13447 avdd.n1122 avdd.t601 27.6955
R13448 avdd.n1119 avdd.t377 27.6955
R13449 avdd.n1119 avdd.t603 27.6955
R13450 avdd.t370 avdd.n1114 27.6955
R13451 avdd.n1114 avdd.t602 27.6955
R13452 avdd.t241 avdd.n1111 27.6955
R13453 avdd.n1111 avdd.t609 27.6955
R13454 avdd.n1108 avdd.t386 27.6955
R13455 avdd.n1108 avdd.t605 27.6955
R13456 avdd.n1105 avdd.t250 27.6955
R13457 avdd.n1105 avdd.t611 27.6955
R13458 avdd.n1169 avdd.t268 27.6955
R13459 avdd.n1169 avdd.t612 27.6955
R13460 avdd.n1021 avdd.t607 27.6955
R13461 avdd.n1021 avdd.t245 27.6955
R13462 avdd.n1023 avdd.t610 27.6955
R13463 avdd.n1023 avdd.t255 27.6955
R13464 avdd.n1025 avdd.t608 27.6955
R13465 avdd.n1025 avdd.t252 27.6955
R13466 avdd.n1027 avdd.t616 27.6955
R13467 avdd.n1027 avdd.t289 27.6955
R13468 avdd.n1029 avdd.t202 27.6955
R13469 avdd.n1029 avdd.t309 27.6955
R13470 avdd.n1031 avdd.t203 27.6955
R13471 avdd.n1031 avdd.t312 27.6955
R13472 avdd.n1033 avdd.t178 27.6955
R13473 avdd.n1033 avdd.t327 27.6955
R13474 avdd.n1035 avdd.t204 27.6955
R13475 avdd.n1035 avdd.t322 27.6955
R13476 avdd.n1037 avdd.t184 27.6955
R13477 avdd.n1037 avdd.t383 27.6955
R13478 avdd.n1039 avdd.t181 27.6955
R13479 avdd.n1039 avdd.t335 27.6955
R13480 avdd.n1041 avdd.t185 27.6955
R13481 avdd.n1041 avdd.t388 27.6955
R13482 avdd.n1044 avdd.t189 27.6955
R13483 avdd.n1044 avdd.t222 27.6955
R13484 avdd.n1145 avdd.t48 27.6955
R13485 avdd.n1145 avdd.t58 27.6955
R13486 avdd.n1147 avdd.t56 27.6955
R13487 avdd.n1147 avdd.t50 27.6955
R13488 avdd.n1149 avdd.t60 27.6955
R13489 avdd.n1149 avdd.t52 27.6955
R13490 avdd.n1151 avdd.t62 27.6955
R13491 avdd.n1151 avdd.t421 27.6955
R13492 avdd.n1516 avdd.t77 27.6955
R13493 avdd.n1516 avdd.t651 27.6955
R13494 avdd.n1514 avdd.t75 27.6955
R13495 avdd.n1514 avdd.t649 27.6955
R13496 avdd.n1512 avdd.t76 27.6955
R13497 avdd.n1512 avdd.t650 27.6955
R13498 avdd.n1510 avdd.t74 27.6955
R13499 avdd.n1510 avdd.t648 27.6955
R13500 avdd.n1508 avdd.t633 27.6955
R13501 avdd.n1508 avdd.t71 27.6955
R13502 avdd.n1506 avdd.t643 27.6955
R13503 avdd.n1506 avdd.t79 27.6955
R13504 avdd.n1504 avdd.t631 27.6955
R13505 avdd.n1504 avdd.t70 27.6955
R13506 avdd.n1502 avdd.t642 27.6955
R13507 avdd.n1502 avdd.t69 27.6955
R13508 avdd.n1500 avdd.t641 27.6955
R13509 avdd.n1500 avdd.t68 27.6955
R13510 avdd.n1498 avdd.t640 27.6955
R13511 avdd.n1498 avdd.t66 27.6955
R13512 avdd.n1262 avdd.t630 27.6955
R13513 avdd.n1262 avdd.t88 27.6955
R13514 avdd.n1612 avdd.t652 27.6955
R13515 avdd.n1612 avdd.t82 27.6955
R13516 avdd.t362 avdd.n1560 27.6955
R13517 avdd.n1560 avdd.t85 27.6955
R13518 avdd.n1557 avdd.t346 27.6955
R13519 avdd.n1557 avdd.t83 27.6955
R13520 avdd.n1554 avdd.t352 27.6955
R13521 avdd.n1554 avdd.t84 27.6955
R13522 avdd.t344 avdd.n1549 27.6955
R13523 avdd.n1549 avdd.t81 27.6955
R13524 avdd.t270 avdd.n1546 27.6955
R13525 avdd.n1546 avdd.t639 27.6955
R13526 avdd.n1543 avdd.t325 27.6955
R13527 avdd.n1543 avdd.t647 27.6955
R13528 avdd.n1540 avdd.t266 27.6955
R13529 avdd.n1540 avdd.t638 27.6955
R13530 avdd.t320 avdd.n1535 27.6955
R13531 avdd.n1535 avdd.t646 27.6955
R13532 avdd.t302 avdd.n1532 27.6955
R13533 avdd.n1532 avdd.t645 27.6955
R13534 avdd.n1529 avdd.t295 27.6955
R13535 avdd.n1529 avdd.t644 27.6955
R13536 avdd.n1526 avdd.t264 27.6955
R13537 avdd.n1526 avdd.t635 27.6955
R13538 avdd.n1591 avdd.t235 27.6955
R13539 avdd.n1591 avdd.t629 27.6955
R13540 avdd.n1267 avdd.t637 27.6955
R13541 avdd.n1267 avdd.t315 27.6955
R13542 avdd.n1269 avdd.t634 27.6955
R13543 avdd.n1269 avdd.t292 27.6955
R13544 avdd.n1271 avdd.t636 27.6955
R13545 avdd.n1271 avdd.t306 27.6955
R13546 avdd.n1273 avdd.t632 27.6955
R13547 avdd.n1273 avdd.t286 27.6955
R13548 avdd.n1275 avdd.t87 27.6955
R13549 avdd.n1275 avdd.t237 27.6955
R13550 avdd.n1277 avdd.t67 27.6955
R13551 avdd.n1277 avdd.t279 27.6955
R13552 avdd.n1279 avdd.t86 27.6955
R13553 avdd.n1279 avdd.t231 27.6955
R13554 avdd.n1281 avdd.t64 27.6955
R13555 avdd.n1281 avdd.t372 27.6955
R13556 avdd.n1283 avdd.t90 27.6955
R13557 avdd.n1283 avdd.t357 27.6955
R13558 avdd.n1285 avdd.t89 27.6955
R13559 avdd.n1285 avdd.t354 27.6955
R13560 avdd.n1287 avdd.t78 27.6955
R13561 avdd.n1287 avdd.t299 27.6955
R13562 avdd.n1290 avdd.t72 27.6955
R13563 avdd.n1290 avdd.t272 27.6955
R13564 avdd.n1567 avdd.t29 27.6955
R13565 avdd.n1567 avdd.t33 27.6955
R13566 avdd.n1569 avdd.t19 27.6955
R13567 avdd.n1569 avdd.t23 27.6955
R13568 avdd.n1571 avdd.t31 27.6955
R13569 avdd.n1571 avdd.t21 27.6955
R13570 avdd.n1573 avdd.t27 27.6955
R13571 avdd.n1573 avdd.t585 27.6955
R13572 avdd.t318 avdd.n1795 26.7523
R13573 avdd.n1764 avdd.t257 25.5567
R13574 avdd.n1789 avdd.t224 25.5567
R13575 avdd.n1771 avdd.t340 25.4942
R13576 avdd.t533 avdd.t97 25.0145
R13577 avdd.n8 avdd.t164 23.5572
R13578 avdd.n345 avdd.t655 23.5572
R13579 avdd.n317 avdd.t439 23.5572
R13580 avdd.n289 avdd.t15 23.5572
R13581 avdd.n261 avdd.t510 23.5572
R13582 avdd.n233 avdd.t443 23.5572
R13583 avdd.n205 avdd.t217 23.5572
R13584 avdd.n177 avdd.t412 23.5572
R13585 avdd.n149 avdd.t504 23.5572
R13586 avdd.n116 avdd.t214 23.5572
R13587 avdd.n682 avdd.t658 23.5572
R13588 avdd.n654 avdd.t3 23.5572
R13589 avdd.n626 avdd.t156 23.5572
R13590 avdd.n598 avdd.t146 23.5572
R13591 avdd.n570 avdd.t397 23.5572
R13592 avdd.n542 avdd.t592 23.5572
R13593 avdd.n514 avdd.t624 23.5572
R13594 avdd.n486 avdd.t39 23.5572
R13595 avdd.n453 avdd.t134 23.5572
R13596 avdd.t348 avdd.t97 22.3534
R13597 avdd.n1698 avdd.n1695 21.9177
R13598 avdd.n1710 avdd.n1709 20.3986
R13599 avdd.n1709 avdd.n1656 20.2792
R13600 avdd.n108 avdd 20.0949
R13601 avdd.n445 avdd 20.0949
R13602 avdd.n1675 avdd.n1655 19.4414
R13603 avdd.n1685 avdd.n1684 18.824
R13604 avdd.n113 avdd 18.3657
R13605 avdd.n450 avdd 18.3657
R13606 avdd.n8 avdd.t581 17.8272
R13607 avdd.n345 avdd.t11 17.8272
R13608 avdd.n317 avdd.t449 17.8272
R13609 avdd.n289 avdd.t621 17.8272
R13610 avdd.n261 avdd.t148 17.8272
R13611 avdd.n233 avdd.t448 17.8272
R13612 avdd.n205 avdd.t108 17.8272
R13613 avdd.n177 avdd.t208 17.8272
R13614 avdd.n149 avdd.t102 17.8272
R13615 avdd.n116 avdd.t210 17.8272
R13616 avdd.n682 avdd.t499 17.8272
R13617 avdd.n654 avdd.t417 17.8272
R13618 avdd.n626 avdd.t659 17.8272
R13619 avdd.n598 avdd.t128 17.8272
R13620 avdd.n570 avdd.t580 17.8272
R13621 avdd.n542 avdd.t577 17.8272
R13622 avdd.n514 avdd.t453 17.8272
R13623 avdd.n486 avdd.t509 17.8272
R13624 avdd.n453 avdd.t130 17.8272
R13625 avdd.n1452 avdd.t549 17.8272
R13626 avdd.n1452 avdd.t563 17.8272
R13627 avdd.n1453 avdd.t547 17.8272
R13628 avdd.n1453 avdd.t569 17.8272
R13629 avdd.n1454 avdd.t565 17.8272
R13630 avdd.n1454 avdd.t545 17.8272
R13631 avdd.n1455 avdd.t561 17.8272
R13632 avdd.n1455 avdd.t539 17.8272
R13633 avdd.n1456 avdd.t557 17.8272
R13634 avdd.n1456 avdd.t567 17.8272
R13635 avdd.n1457 avdd.t553 17.8272
R13636 avdd.n1457 avdd.t555 17.8272
R13637 avdd.n1458 avdd.t559 17.8272
R13638 avdd.n1458 avdd.t551 17.8272
R13639 avdd.n1468 avdd.t116 17.8272
R13640 avdd.n1468 avdd.t118 17.8272
R13641 avdd.n1161 avdd.n1157 17.7802
R13642 avdd.n1201 avdd.n996 17.7802
R13643 avdd.n1583 avdd.n1579 17.7802
R13644 avdd.n1623 avdd.n1242 17.7802
R13645 avdd.n33 avdd.n32 17.7258
R13646 avdd.n369 avdd.n368 17.7258
R13647 avdd.n341 avdd.n340 17.7258
R13648 avdd.n313 avdd.n312 17.7258
R13649 avdd.n285 avdd.n284 17.7258
R13650 avdd.n257 avdd.n256 17.7258
R13651 avdd.n229 avdd.n228 17.7258
R13652 avdd.n201 avdd.n200 17.7258
R13653 avdd.n173 avdd.n172 17.7258
R13654 avdd.n145 avdd.n144 17.7258
R13655 avdd.n706 avdd.n705 17.7258
R13656 avdd.n678 avdd.n677 17.7258
R13657 avdd.n650 avdd.n649 17.7258
R13658 avdd.n622 avdd.n621 17.7258
R13659 avdd.n594 avdd.n593 17.7258
R13660 avdd.n566 avdd.n565 17.7258
R13661 avdd.n538 avdd.n537 17.7258
R13662 avdd.n510 avdd.n509 17.7258
R13663 avdd.n482 avdd.n481 17.7258
R13664 avdd.n113 avdd.n112 17.3701
R13665 avdd.n112 avdd.n107 17.3701
R13666 avdd.n450 avdd.n449 17.3701
R13667 avdd.n449 avdd.n444 17.3701
R13668 avdd.n370 avdd 16.7739
R13669 avdd.n1791 avdd.n1754 16.6169
R13670 avdd.t95 avdd.t505 16.4991
R13671 avdd.n1791 avdd.n1780 16.3798
R13672 avdd.n1737 avdd.n1736 14.9605
R13673 avdd.n1744 avdd.n1743 14.9605
R13674 avdd.n1672 avdd.n1667 14.6829
R13675 avdd.n1761 avdd.n1760 14.6449
R13676 avdd.n1404 avdd.t560 14.6159
R13677 avdd.n1435 avdd.t540 14.6159
R13678 avdd.n988 avdd.t220 14.6083
R13679 avdd.n1168 avdd.t267 14.6083
R13680 avdd.n1234 avdd.t271 14.6083
R13681 avdd.n1590 avdd.t233 14.6083
R13682 avdd.n1699 avdd.n1698 14.4431
R13683 avdd.n1219 avdd.t308 14.4262
R13684 avdd.n1217 avdd.t311 14.4262
R13685 avdd.n1215 avdd.t326 14.4262
R13686 avdd.n1213 avdd.t321 14.4262
R13687 avdd.n1211 avdd.t382 14.4262
R13688 avdd.n1209 avdd.t334 14.4262
R13689 avdd.n1207 avdd.t387 14.4262
R13690 avdd.n1126 avdd.t363 14.4262
R13691 avdd.n1121 avdd.t365 14.4262
R13692 avdd.n1118 avdd.t376 14.4262
R13693 avdd.n1115 avdd.t369 14.4262
R13694 avdd.n1112 avdd.t239 14.4262
R13695 avdd.n1107 avdd.t385 14.4262
R13696 avdd.n1104 avdd.t249 14.4262
R13697 avdd.n1641 avdd.t236 14.4262
R13698 avdd.n1639 avdd.t278 14.4262
R13699 avdd.n1637 avdd.t229 14.4262
R13700 avdd.n1635 avdd.t371 14.4262
R13701 avdd.n1633 avdd.t356 14.4262
R13702 avdd.n1631 avdd.t353 14.4262
R13703 avdd.n1629 avdd.t298 14.4262
R13704 avdd.n1547 avdd.t269 14.4262
R13705 avdd.n1542 avdd.t324 14.4262
R13706 avdd.n1539 avdd.t265 14.4262
R13707 avdd.n1536 avdd.t319 14.4262
R13708 avdd.n1533 avdd.t301 14.4262
R13709 avdd.n1528 avdd.t294 14.4262
R13710 avdd.n1525 avdd.t263 14.4262
R13711 avdd.n1227 avdd.t244 14.4191
R13712 avdd.n1225 avdd.t254 14.4191
R13713 avdd.n1223 avdd.t251 14.4191
R13714 avdd.n1221 avdd.t288 14.4191
R13715 avdd.n1140 avdd.t276 14.4191
R13716 avdd.n1135 avdd.t283 14.4191
R13717 avdd.n1132 avdd.t281 14.4191
R13718 avdd.n1129 avdd.t349 14.4191
R13719 avdd.n1649 avdd.t314 14.4191
R13720 avdd.n1647 avdd.t291 14.4191
R13721 avdd.n1645 avdd.t305 14.4191
R13722 avdd.n1643 avdd.t285 14.4191
R13723 avdd.n1561 avdd.t361 14.4191
R13724 avdd.n1556 avdd.t345 14.4191
R13725 avdd.n1553 avdd.t351 14.4191
R13726 avdd.n1550 avdd.t343 14.4191
R13727 avdd.n1779 avdd.n1760 14.4078
R13728 avdd.n1797 avdd.n1796 14.2313
R13729 avdd.t318 avdd.n1797 14.2313
R13730 avdd.n1799 avdd.n1798 14.2313
R13731 avdd.n1798 avdd.t318 14.2313
R13732 avdd.n1682 avdd.n1673 14.1829
R13733 avdd.n1154 avdd.n1153 14.0622
R13734 avdd.n1576 avdd.n1575 14.0622
R13735 avdd.n1683 avdd.n709 13.9971
R13736 avdd.n1862 avdd.n1861 13.8347
R13737 avdd.n1852 avdd.n1851 13.8322
R13738 avdd.n984 avdd.n983 13.822
R13739 avdd.n1854 avdd.n985 13.822
R13740 avdd.n1206 avdd.n1205 13.8005
R13741 avdd.n1193 avdd.n1192 13.8005
R13742 avdd.n1059 avdd.n1015 13.8005
R13743 avdd.n1043 avdd.n990 13.8005
R13744 avdd.n1166 avdd.n1165 13.8005
R13745 avdd.n1143 avdd.n1073 13.8005
R13746 avdd.n1628 avdd.n1627 13.8005
R13747 avdd.n1615 avdd.n1614 13.8005
R13748 avdd.n1305 avdd.n1261 13.8005
R13749 avdd.n1289 avdd.n1236 13.8005
R13750 avdd.n1588 avdd.n1587 13.8005
R13751 avdd.n1565 avdd.n1319 13.8005
R13752 avdd.n128 avdd.t209 13.7868
R13753 avdd.n465 avdd.t129 13.7868
R13754 avdd.n1058 avdd.n1018 13.436
R13755 avdd.n1185 avdd.n1046 13.436
R13756 avdd.n1172 avdd.n1171 13.436
R13757 avdd.n1304 avdd.n1264 13.436
R13758 avdd.n1607 avdd.n1292 13.436
R13759 avdd.n1594 avdd.n1593 13.436
R13760 avdd.n1175 avdd.n1174 13.177
R13761 avdd.n1597 avdd.n1596 13.177
R13762 avdd.n1066 avdd.n1065 13.0943
R13763 avdd.n1065 avdd.n1064 13.0943
R13764 avdd.n1312 avdd.n1311 13.0943
R13765 avdd.n1311 avdd.n1310 13.0943
R13766 avdd.n1447 avdd.t113 12.789
R13767 avdd.n32 avdd.n31 12.541
R13768 avdd.n368 avdd.n367 12.541
R13769 avdd.n340 avdd.n339 12.541
R13770 avdd.n312 avdd.n311 12.541
R13771 avdd.n284 avdd.n283 12.541
R13772 avdd.n256 avdd.n255 12.541
R13773 avdd.n228 avdd.n227 12.541
R13774 avdd.n200 avdd.n199 12.541
R13775 avdd.n172 avdd.n171 12.541
R13776 avdd.n144 avdd.n143 12.541
R13777 avdd.n705 avdd.n704 12.541
R13778 avdd.n677 avdd.n676 12.541
R13779 avdd.n649 avdd.n648 12.541
R13780 avdd.n621 avdd.n620 12.541
R13781 avdd.n593 avdd.n592 12.541
R13782 avdd.n565 avdd.n564 12.541
R13783 avdd.n537 avdd.n536 12.541
R13784 avdd.n509 avdd.n508 12.541
R13785 avdd.n481 avdd.n480 12.541
R13786 avdd.n24 avdd 12.424
R13787 avdd.n360 avdd 12.424
R13788 avdd.n332 avdd 12.424
R13789 avdd.n304 avdd 12.424
R13790 avdd.n276 avdd 12.424
R13791 avdd.n248 avdd 12.424
R13792 avdd.n220 avdd 12.424
R13793 avdd.n192 avdd 12.424
R13794 avdd.n164 avdd 12.424
R13795 avdd.n136 avdd 12.424
R13796 avdd.n697 avdd 12.424
R13797 avdd.n669 avdd 12.424
R13798 avdd.n641 avdd 12.424
R13799 avdd.n613 avdd 12.424
R13800 avdd.n585 avdd 12.424
R13801 avdd.n557 avdd 12.424
R13802 avdd.n529 avdd 12.424
R13803 avdd.n501 avdd 12.424
R13804 avdd.n473 avdd 12.424
R13805 avdd.n1681 avdd.n1671 11.2946
R13806 avdd.n1695 avdd.n1656 11.1593
R13807 avdd.n1759 avdd.n1758 11.0005
R13808 avdd.n1793 avdd.n1792 11.0005
R13809 avdd.n1066 avdd.n1012 10.9402
R13810 avdd.n1064 avdd.n1012 10.9402
R13811 avdd.n1312 avdd.n1258 10.9402
R13812 avdd.n1310 avdd.n1258 10.9402
R13813 avdd.n1845 avdd.n1844 10.8829
R13814 avdd.n1842 avdd.n1837 10.8829
R13815 avdd.n1857 avdd.n1856 10.8829
R13816 avdd.n1859 avdd.n1858 10.8829
R13817 avdd.n1746 avdd.n1745 10.2783
R13818 avdd.n1748 avdd.n1747 10.2783
R13819 avdd.n1749 avdd.n1748 10.2783
R13820 avdd.n1727 avdd.n1724 10.2783
R13821 avdd.n1728 avdd.n1727 10.2783
R13822 avdd.n1722 avdd.n1719 10.2783
R13823 avdd.n1755 avdd.n1722 10.2783
R13824 avdd.n1758 avdd.n1757 10.2783
R13825 avdd.n1794 avdd.n1793 10.2783
R13826 avdd.n1795 avdd.n1794 10.2783
R13827 avdd.t135 avdd.t211 10.0269
R13828 avdd.t570 avdd.t131 10.0269
R13829 avdd.n1188 avdd.n1019 9.71534
R13830 avdd.n1610 avdd.n1265 9.71534
R13831 avdd.n29 avdd.n28 9.5406
R13832 avdd.n365 avdd.n364 9.5406
R13833 avdd.n337 avdd.n336 9.5406
R13834 avdd.n309 avdd.n308 9.5406
R13835 avdd.n281 avdd.n280 9.5406
R13836 avdd.n253 avdd.n252 9.5406
R13837 avdd.n225 avdd.n224 9.5406
R13838 avdd.n197 avdd.n196 9.5406
R13839 avdd.n169 avdd.n168 9.5406
R13840 avdd.n141 avdd.n140 9.5406
R13841 avdd.n702 avdd.n701 9.5406
R13842 avdd.n674 avdd.n673 9.5406
R13843 avdd.n646 avdd.n645 9.5406
R13844 avdd.n618 avdd.n617 9.5406
R13845 avdd.n590 avdd.n589 9.5406
R13846 avdd.n562 avdd.n561 9.5406
R13847 avdd.n534 avdd.n533 9.5406
R13848 avdd.n506 avdd.n505 9.5406
R13849 avdd.n478 avdd.n477 9.5406
R13850 avdd.n1666 avdd.n709 9.42955
R13851 avdd.n1692 avdd.n1691 9.41227
R13852 avdd.n30 avdd.n29 9.3005
R13853 avdd.n29 avdd.n27 9.3005
R13854 avdd.n16 avdd.n15 9.3005
R13855 avdd.n17 avdd.n16 9.3005
R13856 avdd.n20 avdd.n19 9.3005
R13857 avdd.n18 avdd.n6 9.3005
R13858 avdd.n13 avdd.n12 9.3005
R13859 avdd.n14 avdd.n1 9.3005
R13860 avdd.n26 avdd.n25 9.3005
R13861 avdd.n24 avdd.n0 9.3005
R13862 avdd.n114 avdd.n107 9.3005
R13863 avdd.n142 avdd.n141 9.3005
R13864 avdd.n141 avdd.n139 9.3005
R13865 avdd.n170 avdd.n169 9.3005
R13866 avdd.n169 avdd.n167 9.3005
R13867 avdd.n198 avdd.n197 9.3005
R13868 avdd.n197 avdd.n195 9.3005
R13869 avdd.n226 avdd.n225 9.3005
R13870 avdd.n225 avdd.n223 9.3005
R13871 avdd.n254 avdd.n253 9.3005
R13872 avdd.n253 avdd.n251 9.3005
R13873 avdd.n282 avdd.n281 9.3005
R13874 avdd.n281 avdd.n279 9.3005
R13875 avdd.n310 avdd.n309 9.3005
R13876 avdd.n309 avdd.n307 9.3005
R13877 avdd.n338 avdd.n337 9.3005
R13878 avdd.n337 avdd.n335 9.3005
R13879 avdd.n366 avdd.n365 9.3005
R13880 avdd.n365 avdd.n363 9.3005
R13881 avdd.n114 avdd.n113 9.3005
R13882 avdd.n121 avdd.n120 9.3005
R13883 avdd.n122 avdd.n121 9.3005
R13884 avdd.n153 avdd.n152 9.3005
R13885 avdd.n152 avdd.n151 9.3005
R13886 avdd.n181 avdd.n180 9.3005
R13887 avdd.n180 avdd.n179 9.3005
R13888 avdd.n209 avdd.n208 9.3005
R13889 avdd.n208 avdd.n207 9.3005
R13890 avdd.n237 avdd.n236 9.3005
R13891 avdd.n236 avdd.n235 9.3005
R13892 avdd.n265 avdd.n264 9.3005
R13893 avdd.n264 avdd.n263 9.3005
R13894 avdd.n293 avdd.n292 9.3005
R13895 avdd.n292 avdd.n291 9.3005
R13896 avdd.n321 avdd.n320 9.3005
R13897 avdd.n320 avdd.n319 9.3005
R13898 avdd.n349 avdd.n348 9.3005
R13899 avdd.n348 avdd.n347 9.3005
R13900 avdd.n111 avdd.n110 9.3005
R13901 avdd.n115 avdd.n105 9.3005
R13902 avdd.n125 avdd.n124 9.3005
R13903 avdd.n123 avdd.n106 9.3005
R13904 avdd.n118 avdd.n102 9.3005
R13905 avdd.n119 avdd.n99 9.3005
R13906 avdd.n138 avdd.n137 9.3005
R13907 avdd.n136 avdd.n98 9.3005
R13908 avdd.n160 avdd.n159 9.3005
R13909 avdd.n158 avdd.n97 9.3005
R13910 avdd.n157 avdd.n156 9.3005
R13911 avdd.n155 avdd.n154 9.3005
R13912 avdd.n148 avdd.n91 9.3005
R13913 avdd.n166 avdd.n165 9.3005
R13914 avdd.n164 avdd.n90 9.3005
R13915 avdd.n188 avdd.n187 9.3005
R13916 avdd.n186 avdd.n89 9.3005
R13917 avdd.n185 avdd.n184 9.3005
R13918 avdd.n183 avdd.n182 9.3005
R13919 avdd.n176 avdd.n83 9.3005
R13920 avdd.n194 avdd.n193 9.3005
R13921 avdd.n192 avdd.n82 9.3005
R13922 avdd.n216 avdd.n215 9.3005
R13923 avdd.n214 avdd.n81 9.3005
R13924 avdd.n213 avdd.n212 9.3005
R13925 avdd.n211 avdd.n210 9.3005
R13926 avdd.n204 avdd.n75 9.3005
R13927 avdd.n222 avdd.n221 9.3005
R13928 avdd.n220 avdd.n74 9.3005
R13929 avdd.n244 avdd.n243 9.3005
R13930 avdd.n242 avdd.n73 9.3005
R13931 avdd.n241 avdd.n240 9.3005
R13932 avdd.n239 avdd.n238 9.3005
R13933 avdd.n232 avdd.n67 9.3005
R13934 avdd.n250 avdd.n249 9.3005
R13935 avdd.n248 avdd.n66 9.3005
R13936 avdd.n272 avdd.n271 9.3005
R13937 avdd.n270 avdd.n65 9.3005
R13938 avdd.n269 avdd.n268 9.3005
R13939 avdd.n267 avdd.n266 9.3005
R13940 avdd.n260 avdd.n59 9.3005
R13941 avdd.n278 avdd.n277 9.3005
R13942 avdd.n276 avdd.n58 9.3005
R13943 avdd.n300 avdd.n299 9.3005
R13944 avdd.n298 avdd.n57 9.3005
R13945 avdd.n297 avdd.n296 9.3005
R13946 avdd.n295 avdd.n294 9.3005
R13947 avdd.n288 avdd.n51 9.3005
R13948 avdd.n306 avdd.n305 9.3005
R13949 avdd.n304 avdd.n50 9.3005
R13950 avdd.n328 avdd.n327 9.3005
R13951 avdd.n326 avdd.n49 9.3005
R13952 avdd.n325 avdd.n324 9.3005
R13953 avdd.n323 avdd.n322 9.3005
R13954 avdd.n316 avdd.n43 9.3005
R13955 avdd.n334 avdd.n333 9.3005
R13956 avdd.n332 avdd.n42 9.3005
R13957 avdd.n356 avdd.n355 9.3005
R13958 avdd.n354 avdd.n41 9.3005
R13959 avdd.n353 avdd.n352 9.3005
R13960 avdd.n351 avdd.n350 9.3005
R13961 avdd.n344 avdd.n35 9.3005
R13962 avdd.n362 avdd.n361 9.3005
R13963 avdd.n360 avdd.n34 9.3005
R13964 avdd.n451 avdd.n444 9.3005
R13965 avdd.n479 avdd.n478 9.3005
R13966 avdd.n478 avdd.n476 9.3005
R13967 avdd.n507 avdd.n506 9.3005
R13968 avdd.n506 avdd.n504 9.3005
R13969 avdd.n535 avdd.n534 9.3005
R13970 avdd.n534 avdd.n532 9.3005
R13971 avdd.n563 avdd.n562 9.3005
R13972 avdd.n562 avdd.n560 9.3005
R13973 avdd.n591 avdd.n590 9.3005
R13974 avdd.n590 avdd.n588 9.3005
R13975 avdd.n619 avdd.n618 9.3005
R13976 avdd.n618 avdd.n616 9.3005
R13977 avdd.n647 avdd.n646 9.3005
R13978 avdd.n646 avdd.n644 9.3005
R13979 avdd.n675 avdd.n674 9.3005
R13980 avdd.n674 avdd.n672 9.3005
R13981 avdd.n703 avdd.n702 9.3005
R13982 avdd.n702 avdd.n700 9.3005
R13983 avdd.n451 avdd.n450 9.3005
R13984 avdd.n458 avdd.n457 9.3005
R13985 avdd.n459 avdd.n458 9.3005
R13986 avdd.n490 avdd.n489 9.3005
R13987 avdd.n489 avdd.n488 9.3005
R13988 avdd.n518 avdd.n517 9.3005
R13989 avdd.n517 avdd.n516 9.3005
R13990 avdd.n546 avdd.n545 9.3005
R13991 avdd.n545 avdd.n544 9.3005
R13992 avdd.n574 avdd.n573 9.3005
R13993 avdd.n573 avdd.n572 9.3005
R13994 avdd.n602 avdd.n601 9.3005
R13995 avdd.n601 avdd.n600 9.3005
R13996 avdd.n630 avdd.n629 9.3005
R13997 avdd.n629 avdd.n628 9.3005
R13998 avdd.n658 avdd.n657 9.3005
R13999 avdd.n657 avdd.n656 9.3005
R14000 avdd.n686 avdd.n685 9.3005
R14001 avdd.n685 avdd.n684 9.3005
R14002 avdd.n448 avdd.n447 9.3005
R14003 avdd.n452 avdd.n442 9.3005
R14004 avdd.n462 avdd.n461 9.3005
R14005 avdd.n460 avdd.n443 9.3005
R14006 avdd.n455 avdd.n439 9.3005
R14007 avdd.n456 avdd.n436 9.3005
R14008 avdd.n475 avdd.n474 9.3005
R14009 avdd.n473 avdd.n435 9.3005
R14010 avdd.n497 avdd.n496 9.3005
R14011 avdd.n495 avdd.n434 9.3005
R14012 avdd.n494 avdd.n493 9.3005
R14013 avdd.n492 avdd.n491 9.3005
R14014 avdd.n485 avdd.n428 9.3005
R14015 avdd.n503 avdd.n502 9.3005
R14016 avdd.n501 avdd.n427 9.3005
R14017 avdd.n525 avdd.n524 9.3005
R14018 avdd.n523 avdd.n426 9.3005
R14019 avdd.n522 avdd.n521 9.3005
R14020 avdd.n520 avdd.n519 9.3005
R14021 avdd.n513 avdd.n420 9.3005
R14022 avdd.n531 avdd.n530 9.3005
R14023 avdd.n529 avdd.n419 9.3005
R14024 avdd.n553 avdd.n552 9.3005
R14025 avdd.n551 avdd.n418 9.3005
R14026 avdd.n550 avdd.n549 9.3005
R14027 avdd.n548 avdd.n547 9.3005
R14028 avdd.n541 avdd.n412 9.3005
R14029 avdd.n559 avdd.n558 9.3005
R14030 avdd.n557 avdd.n411 9.3005
R14031 avdd.n581 avdd.n580 9.3005
R14032 avdd.n579 avdd.n410 9.3005
R14033 avdd.n578 avdd.n577 9.3005
R14034 avdd.n576 avdd.n575 9.3005
R14035 avdd.n569 avdd.n404 9.3005
R14036 avdd.n587 avdd.n586 9.3005
R14037 avdd.n585 avdd.n403 9.3005
R14038 avdd.n609 avdd.n608 9.3005
R14039 avdd.n607 avdd.n402 9.3005
R14040 avdd.n606 avdd.n605 9.3005
R14041 avdd.n604 avdd.n603 9.3005
R14042 avdd.n597 avdd.n396 9.3005
R14043 avdd.n615 avdd.n614 9.3005
R14044 avdd.n613 avdd.n395 9.3005
R14045 avdd.n637 avdd.n636 9.3005
R14046 avdd.n635 avdd.n394 9.3005
R14047 avdd.n634 avdd.n633 9.3005
R14048 avdd.n632 avdd.n631 9.3005
R14049 avdd.n625 avdd.n388 9.3005
R14050 avdd.n643 avdd.n642 9.3005
R14051 avdd.n641 avdd.n387 9.3005
R14052 avdd.n665 avdd.n664 9.3005
R14053 avdd.n663 avdd.n386 9.3005
R14054 avdd.n662 avdd.n661 9.3005
R14055 avdd.n660 avdd.n659 9.3005
R14056 avdd.n653 avdd.n380 9.3005
R14057 avdd.n671 avdd.n670 9.3005
R14058 avdd.n669 avdd.n379 9.3005
R14059 avdd.n693 avdd.n692 9.3005
R14060 avdd.n691 avdd.n378 9.3005
R14061 avdd.n690 avdd.n689 9.3005
R14062 avdd.n688 avdd.n687 9.3005
R14063 avdd.n681 avdd.n372 9.3005
R14064 avdd.n699 avdd.n698 9.3005
R14065 avdd.n697 avdd.n371 9.3005
R14066 avdd.n1839 avdd.n1836 9.3005
R14067 avdd.n1848 avdd.n1820 9.3005
R14068 avdd.n721 avdd.n720 9.3005
R14069 avdd.n722 avdd.n721 9.3005
R14070 avdd.n712 avdd.n710 9.3005
R14071 avdd.n719 avdd.n718 9.3005
R14072 avdd.n717 avdd.n711 9.3005
R14073 avdd.n1813 avdd.n1812 9.3005
R14074 avdd.n1792 avdd.n1791 9.3005
R14075 avdd.n1760 avdd.n1759 9.3005
R14076 avdd.n1495 avdd.n1494 9.3005
R14077 avdd.n1491 avdd.n1490 9.3005
R14078 avdd.n1489 avdd.n1488 9.3005
R14079 avdd.n1487 avdd.n1327 9.3005
R14080 avdd.n1486 avdd.n1485 9.3005
R14081 avdd.n1376 avdd.n1371 9.3005
R14082 avdd.n1378 avdd.n1377 9.3005
R14083 avdd.n1367 avdd.n1366 9.3005
R14084 avdd.n1386 avdd.n1385 9.3005
R14085 avdd.n1387 avdd.n1365 9.3005
R14086 avdd.n1389 avdd.n1388 9.3005
R14087 avdd.n1362 avdd.n1361 9.3005
R14088 avdd.n1396 avdd.n1395 9.3005
R14089 avdd.n1397 avdd.n1360 9.3005
R14090 avdd.n1399 avdd.n1398 9.3005
R14091 avdd.n1356 avdd.n1355 9.3005
R14092 avdd.n1407 avdd.n1406 9.3005
R14093 avdd.n1408 avdd.n1354 9.3005
R14094 avdd.n1410 avdd.n1409 9.3005
R14095 avdd.n1351 avdd.n1350 9.3005
R14096 avdd.n1417 avdd.n1416 9.3005
R14097 avdd.n1418 avdd.n1349 9.3005
R14098 avdd.n1420 avdd.n1419 9.3005
R14099 avdd.n1345 avdd.n1344 9.3005
R14100 avdd.n1428 avdd.n1427 9.3005
R14101 avdd.n1429 avdd.n1343 9.3005
R14102 avdd.n1431 avdd.n1430 9.3005
R14103 avdd.n1340 avdd.n1339 9.3005
R14104 avdd.n1439 avdd.n1438 9.3005
R14105 avdd.n1440 avdd.n1338 9.3005
R14106 avdd.n1442 avdd.n1441 9.3005
R14107 avdd.n1335 avdd.n1334 9.3005
R14108 avdd.n1450 avdd.n1449 9.3005
R14109 avdd.n1451 avdd.n1332 9.3005
R14110 avdd.n1474 avdd.n1473 9.3005
R14111 avdd.n1472 avdd.n1333 9.3005
R14112 avdd.n1471 avdd.n1330 9.3005
R14113 avdd.n1496 avdd.n1495 9.3005
R14114 avdd.n1324 avdd.n1323 9.3005
R14115 avdd.n1855 avdd.n1854 9.3005
R14116 avdd.n1852 avdd.n726 9.3005
R14117 avdd.n1861 avdd.n1860 9.3005
R14118 avdd.n983 avdd.n729 9.3005
R14119 avdd.n961 avdd.n735 9.3005
R14120 avdd.n962 avdd.n961 9.3005
R14121 avdd.n950 avdd.n742 9.3005
R14122 avdd.n951 avdd.n950 9.3005
R14123 avdd.n750 avdd.n749 9.3005
R14124 avdd.n751 avdd.n750 9.3005
R14125 avdd.n938 avdd.n937 9.3005
R14126 avdd.n937 avdd.n936 9.3005
R14127 avdd.n925 avdd.n762 9.3005
R14128 avdd.n926 avdd.n925 9.3005
R14129 avdd.n770 avdd.n769 9.3005
R14130 avdd.n771 avdd.n770 9.3005
R14131 avdd.n913 avdd.n912 9.3005
R14132 avdd.n912 avdd.n911 9.3005
R14133 avdd.n900 avdd.n782 9.3005
R14134 avdd.n901 avdd.n900 9.3005
R14135 avdd.n790 avdd.n789 9.3005
R14136 avdd.n791 avdd.n790 9.3005
R14137 avdd.n888 avdd.n887 9.3005
R14138 avdd.n887 avdd.n886 9.3005
R14139 avdd.n875 avdd.n802 9.3005
R14140 avdd.n876 avdd.n875 9.3005
R14141 avdd.n810 avdd.n809 9.3005
R14142 avdd.n811 avdd.n810 9.3005
R14143 avdd.n863 avdd.n862 9.3005
R14144 avdd.n862 avdd.n861 9.3005
R14145 avdd.n850 avdd.n822 9.3005
R14146 avdd.n851 avdd.n850 9.3005
R14147 avdd.n830 avdd.n829 9.3005
R14148 avdd.n831 avdd.n830 9.3005
R14149 avdd.n838 avdd.n837 9.3005
R14150 avdd.n837 avdd.n836 9.3005
R14151 avdd.n967 avdd.n966 9.3005
R14152 avdd.n965 avdd.n731 9.3005
R14153 avdd.n964 avdd.n963 9.3005
R14154 avdd.n960 avdd.n959 9.3005
R14155 avdd.n737 avdd.n736 9.3005
R14156 avdd.n953 avdd.n952 9.3005
R14157 avdd.n949 avdd.n948 9.3005
R14158 avdd.n744 avdd.n743 9.3005
R14159 avdd.n748 avdd.n747 9.3005
R14160 avdd.n941 avdd.n752 9.3005
R14161 avdd.n940 avdd.n939 9.3005
R14162 avdd.n754 avdd.n753 9.3005
R14163 avdd.n935 avdd.n934 9.3005
R14164 avdd.n756 avdd.n755 9.3005
R14165 avdd.n928 avdd.n927 9.3005
R14166 avdd.n924 avdd.n923 9.3005
R14167 avdd.n764 avdd.n763 9.3005
R14168 avdd.n768 avdd.n767 9.3005
R14169 avdd.n916 avdd.n772 9.3005
R14170 avdd.n915 avdd.n914 9.3005
R14171 avdd.n774 avdd.n773 9.3005
R14172 avdd.n910 avdd.n909 9.3005
R14173 avdd.n776 avdd.n775 9.3005
R14174 avdd.n903 avdd.n902 9.3005
R14175 avdd.n899 avdd.n898 9.3005
R14176 avdd.n784 avdd.n783 9.3005
R14177 avdd.n788 avdd.n787 9.3005
R14178 avdd.n891 avdd.n792 9.3005
R14179 avdd.n890 avdd.n889 9.3005
R14180 avdd.n794 avdd.n793 9.3005
R14181 avdd.n885 avdd.n884 9.3005
R14182 avdd.n796 avdd.n795 9.3005
R14183 avdd.n878 avdd.n877 9.3005
R14184 avdd.n874 avdd.n873 9.3005
R14185 avdd.n804 avdd.n803 9.3005
R14186 avdd.n808 avdd.n807 9.3005
R14187 avdd.n866 avdd.n812 9.3005
R14188 avdd.n865 avdd.n864 9.3005
R14189 avdd.n814 avdd.n813 9.3005
R14190 avdd.n860 avdd.n859 9.3005
R14191 avdd.n816 avdd.n815 9.3005
R14192 avdd.n853 avdd.n852 9.3005
R14193 avdd.n849 avdd.n848 9.3005
R14194 avdd.n824 avdd.n823 9.3005
R14195 avdd.n828 avdd.n827 9.3005
R14196 avdd.n841 avdd.n832 9.3005
R14197 avdd.n840 avdd.n839 9.3005
R14198 avdd.n835 avdd.n834 9.3005
R14199 avdd.n1712 avdd.n1711 9.27144
R14200 avdd.n1853 avdd.n1852 9.2699
R14201 avdd.n1854 avdd.n1853 9.2699
R14202 avdd.n1683 avdd.n1682 8.94982
R14203 avdd.n1002 avdd.n1000 8.40959
R14204 avdd.n1002 avdd.n996 8.40959
R14205 avdd.n1006 avdd.n1001 8.40959
R14206 avdd.n1006 avdd.n996 8.40959
R14207 avdd.n1160 avdd.n1159 8.40959
R14208 avdd.n1161 avdd.n1160 8.40959
R14209 avdd.n1200 avdd.n1199 8.40959
R14210 avdd.n1201 avdd.n1200 8.40959
R14211 avdd.n1248 avdd.n1246 8.40959
R14212 avdd.n1248 avdd.n1242 8.40959
R14213 avdd.n1252 avdd.n1247 8.40959
R14214 avdd.n1252 avdd.n1242 8.40959
R14215 avdd.n1582 avdd.n1581 8.40959
R14216 avdd.n1583 avdd.n1582 8.40959
R14217 avdd.n1622 avdd.n1621 8.40959
R14218 avdd.n1623 avdd.n1622 8.40959
R14219 avdd.n1173 avdd.n1056 8.24855
R14220 avdd.n1595 avdd.n1302 8.24855
R14221 avdd.n1232 avdd.n1231 8.24253
R14222 avdd.n1654 avdd.n1653 8.24253
R14223 avdd.n1183 avdd.n1046 8.18605
R14224 avdd.n1605 avdd.n1292 8.18605
R14225 avdd.n1184 avdd.n1183 8.17238
R14226 avdd.n1606 avdd.n1605 8.17238
R14227 avdd.n1173 avdd.n1172 8.10988
R14228 avdd.n1595 avdd.n1594 8.10988
R14229 avdd.n1817 avdd.n1816 7.90948
R14230 avdd.n1143 avdd.n1142 7.90079
R14231 avdd.n1565 avdd.n1564 7.68198
R14232 avdd.n1813 avdd.n1717 7.55653
R14233 avdd.n1730 avdd.n1717 7.55653
R14234 avdd.n1809 avdd.n1808 7.4005
R14235 avdd.t348 avdd.n1809 7.4005
R14236 avdd.n1811 avdd.n1810 7.4005
R14237 avdd.n1810 avdd.t348 7.4005
R14238 avdd.n1383 avdd.t550 7.30819
R14239 avdd.t544 avdd.n1347 7.30819
R14240 avdd.n1057 avdd.n1046 7.29542
R14241 avdd.n1303 avdd.n1292 7.29542
R14242 avdd.n1817 avdd.n985 7.06613
R14243 avdd.n1730 avdd.n1718 7.06516
R14244 avdd.n1813 avdd.n1718 7.06516
R14245 avdd.n28 avdd 7.01471
R14246 avdd.n364 avdd 7.01471
R14247 avdd.n336 avdd 7.01471
R14248 avdd.n308 avdd 7.01471
R14249 avdd.n280 avdd 7.01471
R14250 avdd.n252 avdd 7.01471
R14251 avdd.n224 avdd 7.01471
R14252 avdd.n196 avdd 7.01471
R14253 avdd.n168 avdd 7.01471
R14254 avdd.n140 avdd 7.01471
R14255 avdd.n701 avdd 7.01471
R14256 avdd.n673 avdd 7.01471
R14257 avdd.n645 avdd 7.01471
R14258 avdd.n617 avdd 7.01471
R14259 avdd.n589 avdd 7.01471
R14260 avdd.n561 avdd 7.01471
R14261 avdd.n533 avdd 7.01471
R14262 avdd.n505 avdd 7.01471
R14263 avdd.n477 avdd 7.01471
R14264 avdd.n1172 avdd.n1058 6.77003
R14265 avdd.n1056 avdd.n1055 6.77003
R14266 avdd.n1594 avdd.n1304 6.77003
R14267 avdd.n1302 avdd.n1301 6.77003
R14268 avdd.n1075 avdd.n1070 6.60764
R14269 avdd.n1157 avdd.n1070 6.60764
R14270 avdd.n1156 avdd.n1155 6.60764
R14271 avdd.n1157 avdd.n1156 6.60764
R14272 avdd.n1321 avdd.n1316 6.60764
R14273 avdd.n1579 avdd.n1316 6.60764
R14274 avdd.n1578 avdd.n1577 6.60764
R14275 avdd.n1579 avdd.n1578 6.60764
R14276 avdd.n1184 avdd.n1047 6.59816
R14277 avdd.n1606 avdd.n1293 6.59816
R14278 avdd.n1188 avdd.n1187 6.47706
R14279 avdd.n1610 avdd.n1609 6.47706
R14280 avdd.n1375 avdd.n1372 6.11192
R14281 avdd.n7 avdd 5.7342
R14282 avdd.n1850 avdd.n1849 5.7183
R14283 avdd.n1765 avdd.n1764 5.70732
R14284 avdd.n1790 avdd.n1789 5.70732
R14285 avdd.n1772 avdd.n1771 5.70732
R14286 avdd.n1765 avdd.n1760 5.70369
R14287 avdd.n1836 avdd.n1835 5.70305
R14288 avdd.n1791 avdd.n1790 5.70274
R14289 avdd.n1731 avdd.n1730 5.70242
R14290 avdd.n1849 avdd.n1848 5.6605
R14291 avdd.n1814 avdd.n1813 5.6605
R14292 avdd.n1777 avdd.n1776 5.6605
R14293 avdd.n1833 avdd.t479 5.5395
R14294 avdd.n1833 avdd.t461 5.5395
R14295 avdd.n1831 avdd.t483 5.5395
R14296 avdd.n1831 avdd.t463 5.5395
R14297 avdd.n1829 avdd.t471 5.5395
R14298 avdd.n1829 avdd.t467 5.5395
R14299 avdd.n1827 avdd.t473 5.5395
R14300 avdd.n1827 avdd.t457 5.5395
R14301 avdd.n1825 avdd.t477 5.5395
R14302 avdd.n1825 avdd.t459 5.5395
R14303 avdd.n1823 avdd.t465 5.5395
R14304 avdd.n1823 avdd.t481 5.5395
R14305 avdd.n1821 avdd.t469 5.5395
R14306 avdd.n1821 avdd.t485 5.5395
R14307 avdd.n1773 avdd.t433 5.5395
R14308 avdd.t331 avdd.n1773 5.5395
R14309 avdd.n1715 avdd.t339 5.5395
R14310 avdd.n1715 avdd.t532 5.5395
R14311 avdd.n1739 avdd.t516 5.5395
R14312 avdd.n1739 avdd.t522 5.5395
R14313 avdd.n1741 avdd.t524 5.5395
R14314 avdd.n1741 avdd.t490 5.5395
R14315 avdd.n1770 avdd.t403 5.5395
R14316 avdd.n1770 avdd.t342 5.5395
R14317 avdd.n1766 avdd.t407 5.5395
R14318 avdd.n1766 avdd.t259 5.5395
R14319 avdd.t342 avdd.n1769 5.5395
R14320 avdd.n1769 avdd.t405 5.5395
R14321 avdd.n1774 avdd.t331 5.5395
R14322 avdd.n1774 avdd.t401 5.5395
R14323 avdd.n1781 avdd.t425 5.5395
R14324 avdd.n1781 avdd.t427 5.5395
R14325 avdd.n1783 avdd.t98 5.5395
R14326 avdd.n1783 avdd.t429 5.5395
R14327 avdd.n1785 avdd.t431 5.5395
R14328 avdd.n1785 avdd.t96 5.5395
R14329 avdd.t226 avdd.n1788 5.5395
R14330 avdd.n1788 avdd.t435 5.5395
R14331 avdd.n1847 avdd.n1836 5.48326
R14332 avdd.n1848 avdd.n1847 5.48326
R14333 avdd.n739 avdd.t408 5.48127
R14334 avdd.t121 avdd.n956 5.48127
R14335 avdd.n945 avdd.t205 5.48127
R14336 avdd.n758 avdd.t16 5.48127
R14337 avdd.t105 avdd.n931 5.48127
R14338 avdd.n920 avdd.t574 5.48127
R14339 avdd.n778 avdd.t8 5.48127
R14340 avdd.t572 avdd.n906 5.48127
R14341 avdd.n895 avdd.t125 5.48127
R14342 avdd.n798 avdd.t494 5.48127
R14343 avdd.t622 avdd.n881 5.48127
R14344 avdd.n870 avdd.t111 5.48127
R14345 avdd.n818 avdd.t218 5.48127
R14346 avdd.t536 avdd.n856 5.48127
R14347 avdd.n845 avdd.t486 5.48127
R14348 avdd.n1805 avdd.n1804 5.28621
R14349 avdd.n1804 avdd.t515 5.28621
R14350 avdd.n1803 avdd.n1802 5.28621
R14351 avdd.t515 avdd.n1803 5.28621
R14352 avdd.n1020 avdd.n989 5.22511
R14353 avdd.n1167 avdd.n1019 5.22511
R14354 avdd.n1266 avdd.n1235 5.22511
R14355 avdd.n1589 avdd.n1265 5.22511
R14356 avdd.n1171 avdd.n1170 5.11573
R14357 avdd.n1593 avdd.n1592 5.11573
R14358 avdd.n1067 avdd.n1019 4.98102
R14359 avdd.n1313 avdd.n1265 4.98102
R14360 avdd.n1063 avdd.n1020 4.94972
R14361 avdd.n1309 avdd.n1266 4.94972
R14362 avdd.n1680 avdd.n1677 4.89462
R14363 avdd.n1676 avdd.n1674 4.89462
R14364 avdd.n1158 avdd.n1069 4.86892
R14365 avdd.n1161 avdd.n1158 4.86892
R14366 avdd.n1061 avdd.n995 4.86892
R14367 avdd.n1201 avdd.n995 4.86892
R14368 avdd.n1580 avdd.n1315 4.86892
R14369 avdd.n1583 avdd.n1580 4.86892
R14370 avdd.n1307 avdd.n1241 4.86892
R14371 avdd.n1623 avdd.n1241 4.86892
R14372 avdd.n708 avdd.n707 4.7853
R14373 avdd.n1564 avdd.n1497 4.76569
R14374 avdd.n989 avdd.n988 4.66083
R14375 avdd.n1168 avdd.n1167 4.66083
R14376 avdd.n1235 avdd.n1234 4.66083
R14377 avdd.n1590 avdd.n1589 4.66083
R14378 avdd.n1208 avdd.n1207 4.5005
R14379 avdd.n1210 avdd.n1209 4.5005
R14380 avdd.n1212 avdd.n1211 4.5005
R14381 avdd.n1214 avdd.n1213 4.5005
R14382 avdd.n1216 avdd.n1215 4.5005
R14383 avdd.n1218 avdd.n1217 4.5005
R14384 avdd.n1220 avdd.n1219 4.5005
R14385 avdd.n1222 avdd.n1221 4.5005
R14386 avdd.n1224 avdd.n1223 4.5005
R14387 avdd.n1226 avdd.n1225 4.5005
R14388 avdd.n1228 avdd.n1227 4.5005
R14389 avdd.n1185 avdd.n1184 4.5005
R14390 avdd.n1055 avdd.n1018 4.5005
R14391 avdd.n1171 avdd.n1056 4.5005
R14392 avdd.n1104 avdd.n1060 4.5005
R14393 avdd.n1107 avdd.n1103 4.5005
R14394 avdd.n1113 avdd.n1112 4.5005
R14395 avdd.n1116 avdd.n1115 4.5005
R14396 avdd.n1118 avdd.n1117 4.5005
R14397 avdd.n1121 avdd.n1101 4.5005
R14398 avdd.n1127 avdd.n1126 4.5005
R14399 avdd.n1130 avdd.n1129 4.5005
R14400 avdd.n1132 avdd.n1131 4.5005
R14401 avdd.n1135 avdd.n1099 4.5005
R14402 avdd.n1141 avdd.n1140 4.5005
R14403 avdd.n1189 avdd.n1188 4.5005
R14404 avdd.n1187 avdd.n1186 4.5005
R14405 avdd.n1630 avdd.n1629 4.5005
R14406 avdd.n1632 avdd.n1631 4.5005
R14407 avdd.n1634 avdd.n1633 4.5005
R14408 avdd.n1636 avdd.n1635 4.5005
R14409 avdd.n1638 avdd.n1637 4.5005
R14410 avdd.n1640 avdd.n1639 4.5005
R14411 avdd.n1642 avdd.n1641 4.5005
R14412 avdd.n1644 avdd.n1643 4.5005
R14413 avdd.n1646 avdd.n1645 4.5005
R14414 avdd.n1648 avdd.n1647 4.5005
R14415 avdd.n1650 avdd.n1649 4.5005
R14416 avdd.n1607 avdd.n1606 4.5005
R14417 avdd.n1301 avdd.n1264 4.5005
R14418 avdd.n1593 avdd.n1302 4.5005
R14419 avdd.n1525 avdd.n1306 4.5005
R14420 avdd.n1528 avdd.n1524 4.5005
R14421 avdd.n1534 avdd.n1533 4.5005
R14422 avdd.n1537 avdd.n1536 4.5005
R14423 avdd.n1539 avdd.n1538 4.5005
R14424 avdd.n1542 avdd.n1522 4.5005
R14425 avdd.n1548 avdd.n1547 4.5005
R14426 avdd.n1551 avdd.n1550 4.5005
R14427 avdd.n1553 avdd.n1552 4.5005
R14428 avdd.n1556 avdd.n1520 4.5005
R14429 avdd.n1562 avdd.n1561 4.5005
R14430 avdd.n1611 avdd.n1610 4.5005
R14431 avdd.n1609 avdd.n1608 4.5005
R14432 avdd.n1816 avdd.n1713 4.4965
R14433 avdd.n113 avdd 4.46111
R14434 avdd.n113 avdd 4.46111
R14435 avdd.n450 avdd 4.46111
R14436 avdd.n450 avdd 4.46111
R14437 avdd.n1229 avdd.n1228 4.45347
R14438 avdd.n1097 avdd.n1096 4.45347
R14439 avdd.n1138 avdd.n1098 4.45347
R14440 avdd.n1022 avdd.n987 4.45347
R14441 avdd.n1142 avdd.n1141 4.45347
R14442 avdd.n1651 avdd.n1650 4.45347
R14443 avdd.n1518 avdd.n1517 4.45347
R14444 avdd.n1559 avdd.n1519 4.45347
R14445 avdd.n1268 avdd.n1233 4.45347
R14446 avdd.n1563 avdd.n1562 4.45347
R14447 avdd.n1186 avdd.n1185 4.39112
R14448 avdd.n1608 avdd.n1607 4.39112
R14449 avdd.n1846 avdd.n1838 4.20505
R14450 avdd.n1843 avdd.n1838 4.20505
R14451 avdd.n1841 avdd.n1840 4.20505
R14452 avdd.n1843 avdd.n1841 4.20505
R14453 avdd.n1189 avdd.n1018 4.16066
R14454 avdd.n1611 avdd.n1264 4.16066
R14455 avdd.n1816 avdd.n1815 4.15861
R14456 avdd.n1701 avdd.n1700 4.14168
R14457 avdd.n1815 avdd.n1814 4.01324
R14458 avdd.n1848 avdd.n1819 3.91429
R14459 avdd.n1836 avdd.n1819 3.91429
R14460 avdd.n9 avdd 3.7406
R14461 avdd.n346 avdd 3.7406
R14462 avdd.n318 avdd 3.7406
R14463 avdd.n290 avdd 3.7406
R14464 avdd.n262 avdd 3.7406
R14465 avdd.n234 avdd 3.7406
R14466 avdd.n206 avdd 3.7406
R14467 avdd.n178 avdd 3.7406
R14468 avdd.n150 avdd 3.7406
R14469 avdd.n117 avdd 3.7406
R14470 avdd.n683 avdd 3.7406
R14471 avdd.n655 avdd 3.7406
R14472 avdd.n627 avdd 3.7406
R14473 avdd.n599 avdd 3.7406
R14474 avdd.n571 avdd 3.7406
R14475 avdd.n543 avdd 3.7406
R14476 avdd.n515 avdd 3.7406
R14477 avdd.n487 avdd 3.7406
R14478 avdd.n454 avdd 3.7406
R14479 avdd.n7 avdd 3.56469
R14480 avdd.n7 avdd 3.56469
R14481 avdd.n1671 avdd.n1670 3.55819
R14482 avdd.n1670 avdd.n1669 3.55819
R14483 avdd.n1187 avdd.n1020 3.23878
R14484 avdd.n1609 avdd.n1266 3.23878
R14485 avdd.n1702 avdd.n1701 2.93701
R14486 avdd.n1703 avdd.n1702 2.93701
R14487 avdd.n1176 avdd.n1175 2.80353
R14488 avdd.n1177 avdd.n1176 2.80353
R14489 avdd.n1181 avdd.n1180 2.80353
R14490 avdd.n1180 avdd.n1179 2.80353
R14491 avdd.n1598 avdd.n1597 2.80353
R14492 avdd.n1599 avdd.n1598 2.80353
R14493 avdd.n1603 avdd.n1602 2.80353
R14494 avdd.n1602 avdd.n1601 2.80353
R14495 avdd.n1686 avdd.n1685 2.28445
R14496 avdd.n1687 avdd.n1686 2.28445
R14497 avdd.n1711 avdd.n1710 2.27397
R14498 avdd.n1815 avdd.n1714 1.97988
R14499 avdd.n1761 avdd.n1754 1.97248
R14500 avdd.n1780 avdd.n1779 1.97248
R14501 avdd.n1376 avdd.n1375 1.87847
R14502 avdd.t428 avdd.n1755 1.86325
R14503 avdd.n707 avdd.n370 1.69386
R14504 avdd.n1712 avdd 1.67975
R14505 avdd.n1064 avdd.n1063 1.61378
R14506 avdd.n1310 avdd.n1309 1.61378
R14507 avdd.n1067 avdd.n1066 1.55875
R14508 avdd.n1313 avdd.n1312 1.55875
R14509 avdd.n1657 avdd.n1655 1.5505
R14510 avdd.n1763 avdd.n1762 1.52433
R14511 avdd.n1182 avdd.n1181 1.50638
R14512 avdd.n1604 avdd.n1603 1.50638
R14513 avdd.n727 avdd.n725 1.4805
R14514 avdd.t381 avdd.n727 1.4805
R14515 avdd.n730 avdd.n728 1.4805
R14516 avdd.t381 avdd.n728 1.4805
R14517 avdd.n1778 avdd.n1777 1.31832
R14518 avdd.n983 avdd.n982 1.28283
R14519 avdd.n999 avdd.n997 1.2505
R14520 avdd.n1195 avdd.n997 1.2505
R14521 avdd.n1197 avdd.n1196 1.2505
R14522 avdd.n1196 avdd.n1195 1.2505
R14523 avdd.n1194 avdd.n1193 1.2505
R14524 avdd.n1195 avdd.n1194 1.2505
R14525 avdd.n994 avdd.n992 1.2505
R14526 avdd.n1195 avdd.n994 1.2505
R14527 avdd.n1245 avdd.n1243 1.2505
R14528 avdd.n1617 avdd.n1243 1.2505
R14529 avdd.n1619 avdd.n1618 1.2505
R14530 avdd.n1618 avdd.n1617 1.2505
R14531 avdd.n1616 avdd.n1615 1.2505
R14532 avdd.n1617 avdd.n1616 1.2505
R14533 avdd.n1240 avdd.n1238 1.2505
R14534 avdd.n1617 avdd.n1240 1.2505
R14535 avdd.n984 avdd.n967 1.16964
R14536 avdd.n982 avdd.n981 1.15136
R14537 avdd.n981 avdd.n980 1.15136
R14538 avdd.n980 avdd.n979 1.15136
R14539 avdd.n979 avdd.n978 1.15136
R14540 avdd.n978 avdd.n977 1.15136
R14541 avdd.n977 avdd.n976 1.15136
R14542 avdd.n974 avdd.n973 1.15136
R14543 avdd.n973 avdd.n972 1.15136
R14544 avdd.n972 avdd.n971 1.15136
R14545 avdd.n971 avdd.n970 1.15136
R14546 avdd.n970 avdd.n969 1.15136
R14547 avdd.n969 avdd.n968 1.15136
R14548 avdd.n968 avdd.n724 1.15136
R14549 avdd.n1053 avdd.n1050 1.14248
R14550 avdd.n1052 avdd.n1050 1.14248
R14551 avdd.n1051 avdd.n1049 1.14248
R14552 avdd.n1178 avdd.n1051 1.14248
R14553 avdd.n1299 avdd.n1296 1.14248
R14554 avdd.n1298 avdd.n1296 1.14248
R14555 avdd.n1297 avdd.n1295 1.14248
R14556 avdd.n1600 avdd.n1297 1.14248
R14557 avdd.n1861 avdd.n724 1.13628
R14558 avdd.n1697 avdd.n1665 1.12991
R14559 avdd.n976 avdd.n975 1.0824
R14560 avdd.n1098 avdd.n1097 1.05355
R14561 avdd.n1097 avdd.n987 1.05355
R14562 avdd.n1519 avdd.n1518 1.05355
R14563 avdd.n1518 avdd.n1233 1.05355
R14564 avdd.n1222 avdd.n1220 1.04347
R14565 avdd.n1090 avdd.n1088 1.04347
R14566 avdd.n1030 avdd.n1028 1.04347
R14567 avdd.n1124 avdd.n1100 1.04347
R14568 avdd.n1130 avdd.n1127 1.04347
R14569 avdd.n1644 avdd.n1642 1.04347
R14570 avdd.n1511 avdd.n1509 1.04347
R14571 avdd.n1276 avdd.n1274 1.04347
R14572 avdd.n1545 avdd.n1521 1.04347
R14573 avdd.n1551 avdd.n1548 1.04347
R14574 avdd.n1658 avdd.n986 1.03383
R14575 avdd.n1665 avdd.n1660 0.989805
R14576 avdd.n1704 avdd.n1660 0.989805
R14577 avdd.n370 avdd 0.983
R14578 avdd.n707 avdd 0.983
R14579 avdd.n1680 avdd.n1679 0.954108
R14580 avdd.n1679 avdd.n1678 0.954108
R14581 avdd.n1752 avdd.n1750 0.907363
R14582 avdd.n1756 avdd.n1750 0.907363
R14583 avdd.n1753 avdd.n1751 0.907363
R14584 avdd.n1756 avdd.n1751 0.907363
R14585 avdd.n1850 avdd.n1817 0.90425
R14586 avdd.n1691 avdd.n1690 0.877277
R14587 avdd.n1690 avdd.n1689 0.877277
R14588 avdd avdd.n709 0.876125
R14589 avdd.n985 avdd.n984 0.83425
R14590 avdd.n1055 avdd.n1047 0.773938
R14591 avdd.n1301 avdd.n1293 0.773938
R14592 avdd.n159 avdd 0.755
R14593 avdd.n187 avdd 0.755
R14594 avdd.n215 avdd 0.755
R14595 avdd.n243 avdd 0.755
R14596 avdd.n271 avdd 0.755
R14597 avdd.n299 avdd 0.755
R14598 avdd.n327 avdd 0.755
R14599 avdd.n355 avdd 0.755
R14600 avdd.n496 avdd 0.755
R14601 avdd.n524 avdd 0.755
R14602 avdd.n552 avdd 0.755
R14603 avdd.n580 avdd 0.755
R14604 avdd.n608 avdd 0.755
R14605 avdd.n636 avdd 0.755
R14606 avdd.n664 avdd 0.755
R14607 avdd.n692 avdd 0.755
R14608 avdd.n1186 avdd.n1045 0.725109
R14609 avdd.n1608 avdd.n1291 0.725109
R14610 avdd.n1231 avdd.n1230 0.713391
R14611 avdd.n1228 avdd.n1226 0.713391
R14612 avdd.n1226 avdd.n1224 0.713391
R14613 avdd.n1224 avdd.n1222 0.713391
R14614 avdd.n1220 avdd.n1218 0.713391
R14615 avdd.n1218 avdd.n1216 0.713391
R14616 avdd.n1216 avdd.n1214 0.713391
R14617 avdd.n1214 avdd.n1212 0.713391
R14618 avdd.n1212 avdd.n1210 0.713391
R14619 avdd.n1210 avdd.n1208 0.713391
R14620 avdd.n1096 avdd.n1094 0.713391
R14621 avdd.n1094 avdd.n1092 0.713391
R14622 avdd.n1092 avdd.n1090 0.713391
R14623 avdd.n1088 avdd.n1086 0.713391
R14624 avdd.n1086 avdd.n1084 0.713391
R14625 avdd.n1084 avdd.n1082 0.713391
R14626 avdd.n1082 avdd.n1080 0.713391
R14627 avdd.n1080 avdd.n1078 0.713391
R14628 avdd.n1078 avdd.n1017 0.713391
R14629 avdd.n1024 avdd.n1022 0.713391
R14630 avdd.n1026 avdd.n1024 0.713391
R14631 avdd.n1028 avdd.n1026 0.713391
R14632 avdd.n1032 avdd.n1030 0.713391
R14633 avdd.n1034 avdd.n1032 0.713391
R14634 avdd.n1036 avdd.n1034 0.713391
R14635 avdd.n1038 avdd.n1036 0.713391
R14636 avdd.n1040 avdd.n1038 0.713391
R14637 avdd.n1042 avdd.n1040 0.713391
R14638 avdd.n1138 avdd.n1137 0.713391
R14639 avdd.n1137 avdd.n1134 0.713391
R14640 avdd.n1134 avdd.n1100 0.713391
R14641 avdd.n1124 avdd.n1123 0.713391
R14642 avdd.n1123 avdd.n1120 0.713391
R14643 avdd.n1120 avdd.n1102 0.713391
R14644 avdd.n1110 avdd.n1102 0.713391
R14645 avdd.n1110 avdd.n1109 0.713391
R14646 avdd.n1109 avdd.n1106 0.713391
R14647 avdd.n1141 avdd.n1099 0.713391
R14648 avdd.n1131 avdd.n1099 0.713391
R14649 avdd.n1131 avdd.n1130 0.713391
R14650 avdd.n1127 avdd.n1101 0.713391
R14651 avdd.n1117 avdd.n1101 0.713391
R14652 avdd.n1117 avdd.n1116 0.713391
R14653 avdd.n1116 avdd.n1113 0.713391
R14654 avdd.n1113 avdd.n1103 0.713391
R14655 avdd.n1103 avdd.n1060 0.713391
R14656 avdd.n1653 avdd.n1652 0.713391
R14657 avdd.n1650 avdd.n1648 0.713391
R14658 avdd.n1648 avdd.n1646 0.713391
R14659 avdd.n1646 avdd.n1644 0.713391
R14660 avdd.n1642 avdd.n1640 0.713391
R14661 avdd.n1640 avdd.n1638 0.713391
R14662 avdd.n1638 avdd.n1636 0.713391
R14663 avdd.n1636 avdd.n1634 0.713391
R14664 avdd.n1634 avdd.n1632 0.713391
R14665 avdd.n1632 avdd.n1630 0.713391
R14666 avdd.n1517 avdd.n1515 0.713391
R14667 avdd.n1515 avdd.n1513 0.713391
R14668 avdd.n1513 avdd.n1511 0.713391
R14669 avdd.n1509 avdd.n1507 0.713391
R14670 avdd.n1507 avdd.n1505 0.713391
R14671 avdd.n1505 avdd.n1503 0.713391
R14672 avdd.n1503 avdd.n1501 0.713391
R14673 avdd.n1501 avdd.n1499 0.713391
R14674 avdd.n1499 avdd.n1263 0.713391
R14675 avdd.n1270 avdd.n1268 0.713391
R14676 avdd.n1272 avdd.n1270 0.713391
R14677 avdd.n1274 avdd.n1272 0.713391
R14678 avdd.n1278 avdd.n1276 0.713391
R14679 avdd.n1280 avdd.n1278 0.713391
R14680 avdd.n1282 avdd.n1280 0.713391
R14681 avdd.n1284 avdd.n1282 0.713391
R14682 avdd.n1286 avdd.n1284 0.713391
R14683 avdd.n1288 avdd.n1286 0.713391
R14684 avdd.n1559 avdd.n1558 0.713391
R14685 avdd.n1558 avdd.n1555 0.713391
R14686 avdd.n1555 avdd.n1521 0.713391
R14687 avdd.n1545 avdd.n1544 0.713391
R14688 avdd.n1544 avdd.n1541 0.713391
R14689 avdd.n1541 avdd.n1523 0.713391
R14690 avdd.n1531 avdd.n1523 0.713391
R14691 avdd.n1531 avdd.n1530 0.713391
R14692 avdd.n1530 avdd.n1527 0.713391
R14693 avdd.n1562 avdd.n1520 0.713391
R14694 avdd.n1552 avdd.n1520 0.713391
R14695 avdd.n1552 avdd.n1551 0.713391
R14696 avdd.n1548 avdd.n1522 0.713391
R14697 avdd.n1538 avdd.n1522 0.713391
R14698 avdd.n1538 avdd.n1537 0.713391
R14699 avdd.n1537 avdd.n1534 0.713391
R14700 avdd.n1534 avdd.n1524 0.713391
R14701 avdd.n1524 avdd.n1306 0.713391
R14702 avdd.n1146 avdd.n1144 0.695812
R14703 avdd.n1148 avdd.n1146 0.695812
R14704 avdd.n1150 avdd.n1148 0.695812
R14705 avdd.n1152 avdd.n1150 0.695812
R14706 avdd.n1153 avdd.n1152 0.695812
R14707 avdd.n1568 avdd.n1566 0.695812
R14708 avdd.n1570 avdd.n1568 0.695812
R14709 avdd.n1572 avdd.n1570 0.695812
R14710 avdd.n1574 avdd.n1572 0.695812
R14711 avdd.n1575 avdd.n1574 0.695812
R14712 avdd.n111 avdd 0.664
R14713 avdd.n448 avdd 0.664
R14714 avdd.n1191 avdd.n1189 0.662609
R14715 avdd.n1613 avdd.n1611 0.662609
R14716 avdd.n1863 avdd.n1862 0.624875
R14717 avdd.n1470 avdd 0.576587
R14718 avdd.n708 avdd 0.563625
R14719 avdd.n1668 avdd.n1667 0.56281
R14720 avdd.n1688 avdd.n1668 0.56281
R14721 avdd.n1674 avdd.n1659 0.559412
R14722 avdd.n1661 avdd.n1659 0.559412
R14723 avdd.n1851 avdd.n723 0.55425
R14724 avdd.n1787 avdd.n1786 0.545446
R14725 avdd.n1786 avdd.n1784 0.545446
R14726 avdd.n1784 avdd.n1782 0.545446
R14727 avdd.n1775 avdd.n1772 0.545446
R14728 avdd.n1768 avdd.n1767 0.545446
R14729 avdd.n1142 avdd.n1098 0.527027
R14730 avdd.n1229 avdd.n987 0.527027
R14731 avdd.n1563 avdd.n1519 0.527027
R14732 avdd.n1651 avdd.n1233 0.527027
R14733 avdd.n1460 avdd.n1459 0.526374
R14734 avdd.n1461 avdd.n1460 0.526374
R14735 avdd.n1462 avdd.n1461 0.526374
R14736 avdd.n1463 avdd.n1462 0.526374
R14737 avdd.n1464 avdd.n1463 0.526374
R14738 avdd.n1465 avdd.n1464 0.526374
R14739 avdd.n1466 avdd.n1465 0.49141
R14740 avdd.n1208 avdd.n1206 0.477062
R14741 avdd.n1192 avdd.n1017 0.477062
R14742 avdd.n1043 avdd.n1042 0.477062
R14743 avdd.n1106 avdd.n1059 0.477062
R14744 avdd.n1166 avdd.n1060 0.477062
R14745 avdd.n1630 avdd.n1628 0.477062
R14746 avdd.n1614 avdd.n1263 0.477062
R14747 avdd.n1289 avdd.n1288 0.477062
R14748 avdd.n1527 avdd.n1305 0.477062
R14749 avdd.n1588 avdd.n1306 0.477062
R14750 avdd.n1469 avdd.n1467 0.469796
R14751 avdd.n1664 avdd.n1663 0.444145
R14752 avdd.n1663 avdd.n1662 0.444145
R14753 avdd.n1710 avdd.n1655 0.418878
R14754 avdd.n1713 avdd.n986 0.4145
R14755 avdd.n709 avdd.n708 0.407375
R14756 avdd.n1470 avdd 0.358608
R14757 avdd avdd.n1493 0.357024
R14758 avdd.n1707 avdd.n1706 0.330857
R14759 avdd.n1706 avdd.n1705 0.330857
R14760 avdd.n1470 avdd.n1469 0.325765
R14761 avdd.n1863 avdd 0.32398
R14762 avdd.n1206 avdd.n989 0.318859
R14763 avdd.n1192 avdd.n1191 0.318859
R14764 avdd.n1045 avdd.n1043 0.318859
R14765 avdd.n1170 avdd.n1059 0.318859
R14766 avdd.n1167 avdd.n1166 0.318859
R14767 avdd.n1628 avdd.n1235 0.318859
R14768 avdd.n1614 avdd.n1613 0.318859
R14769 avdd.n1291 avdd.n1289 0.318859
R14770 avdd.n1592 avdd.n1305 0.318859
R14771 avdd.n1589 avdd.n1588 0.318859
R14772 avdd.n1776 avdd.n1714 0.316162
R14773 avdd.n1742 avdd.n1740 0.291392
R14774 avdd.n1740 avdd.n1738 0.291392
R14775 avdd.n1762 avdd.n1761 0.284354
R14776 avdd.n1779 avdd.n1778 0.284354
R14777 avdd.n1862 avdd.n723 0.2805
R14778 avdd.n1776 avdd.n1775 0.273291
R14779 avdd.n1790 avdd.n1787 0.272973
R14780 avdd.n1772 avdd.n1768 0.272973
R14781 avdd.n1767 avdd.n1765 0.272973
R14782 avdd.n1144 avdd.n1143 0.262219
R14783 avdd.n1566 avdd.n1565 0.262219
R14784 avdd.n1488 avdd.n1487 0.26137
R14785 avdd.n1487 avdd.n1486 0.26137
R14786 avdd.n1377 avdd.n1376 0.26137
R14787 avdd.n1377 avdd.n1366 0.26137
R14788 avdd.n1386 avdd.n1366 0.26137
R14789 avdd.n1387 avdd.n1386 0.26137
R14790 avdd.n1388 avdd.n1387 0.26137
R14791 avdd.n1388 avdd.n1361 0.26137
R14792 avdd.n1396 avdd.n1361 0.26137
R14793 avdd.n1397 avdd.n1396 0.26137
R14794 avdd.n1398 avdd.n1397 0.26137
R14795 avdd.n1398 avdd.n1355 0.26137
R14796 avdd.n1407 avdd.n1355 0.26137
R14797 avdd.n1409 avdd.n1408 0.26137
R14798 avdd.n1409 avdd.n1350 0.26137
R14799 avdd.n1417 avdd.n1350 0.26137
R14800 avdd.n1418 avdd.n1417 0.26137
R14801 avdd.n1419 avdd.n1418 0.26137
R14802 avdd.n1419 avdd.n1344 0.26137
R14803 avdd.n1428 avdd.n1344 0.26137
R14804 avdd.n1429 avdd.n1428 0.26137
R14805 avdd.n1430 avdd.n1429 0.26137
R14806 avdd.n1430 avdd.n1339 0.26137
R14807 avdd.n1439 avdd.n1339 0.26137
R14808 avdd.n1440 avdd.n1439 0.26137
R14809 avdd.n1441 avdd.n1440 0.26137
R14810 avdd.n1450 avdd.n1334 0.26137
R14811 avdd.n1451 avdd.n1450 0.26137
R14812 avdd.n1473 avdd.n1451 0.26137
R14813 avdd.n1473 avdd.n1472 0.26137
R14814 avdd.n1472 avdd.n1471 0.26137
R14815 avdd.n1713 avdd.n1712 0.2505
R14816 avdd avdd.n960 0.248811
R14817 avdd avdd.n949 0.248811
R14818 avdd.n752 avdd 0.248811
R14819 avdd avdd.n935 0.248811
R14820 avdd avdd.n924 0.248811
R14821 avdd.n772 avdd 0.248811
R14822 avdd avdd.n910 0.248811
R14823 avdd avdd.n899 0.248811
R14824 avdd.n792 avdd 0.248811
R14825 avdd avdd.n885 0.248811
R14826 avdd avdd.n874 0.248811
R14827 avdd.n812 avdd 0.248811
R14828 avdd avdd.n860 0.248811
R14829 avdd avdd.n849 0.248811
R14830 avdd.n832 avdd 0.248811
R14831 avdd.n1732 avdd.n1731 0.246297
R14832 avdd.n1711 avdd 0.242804
R14833 avdd.n1851 avdd.n1850 0.238625
R14834 avdd.n1782 avdd.n1714 0.229784
R14835 avdd.n1232 avdd.n1229 0.227878
R14836 avdd.n1654 avdd.n1651 0.227878
R14837 avdd.n1840 avdd.n1819 0.227329
R14838 avdd.n1847 avdd.n1846 0.227329
R14839 avdd.n1564 avdd.n1563 0.219304
R14840 avdd.n1743 avdd.n1742 0.1885
R14841 avdd.n1682 avdd.n1681 0.1865
R14842 avdd.n1737 avdd.n1735 0.183736
R14843 avdd.n723 avdd.n722 0.175331
R14844 avdd.n1814 avdd.n1716 0.156108
R14845 avdd.n1183 avdd.n1182 0.152959
R14846 avdd.n1174 avdd.n1173 0.152959
R14847 avdd.n1605 avdd.n1604 0.152959
R14848 avdd.n1596 avdd.n1595 0.152959
R14849 avdd.n1700 avdd.n1699 0.152959
R14850 avdd.n1467 avdd 0.144186
R14851 avdd.n1068 avdd.n1067 0.143577
R14852 avdd.n1314 avdd.n1313 0.143577
R14853 avdd.n1063 avdd.n1062 0.141409
R14854 avdd.n1309 avdd.n1308 0.141409
R14855 avdd avdd.n1466 0.132362
R14856 avdd.n1491 avdd 0.130935
R14857 avdd.n1488 avdd 0.130935
R14858 avdd.n1486 avdd 0.130935
R14859 avdd avdd.n1407 0.130935
R14860 avdd.n1408 avdd 0.130935
R14861 avdd.n1441 avdd 0.130935
R14862 avdd avdd.n1334 0.130935
R14863 avdd.n1493 avdd 0.130673
R14864 avdd.n1801 avdd.n1718 0.126176
R14865 avdd.n1806 avdd.n1717 0.126176
R14866 avdd.n1684 avdd.n1683 0.119731
R14867 avdd.n1822 avdd.n1818 0.113554
R14868 avdd.n1824 avdd.n1822 0.113554
R14869 avdd.n1826 avdd.n1824 0.113554
R14870 avdd.n1828 avdd.n1826 0.113554
R14871 avdd.n1830 avdd.n1828 0.113554
R14872 avdd.n1832 avdd.n1830 0.113554
R14873 avdd.n1834 avdd.n1832 0.113554
R14874 avdd.n1835 avdd.n1834 0.113554
R14875 avdd.n1735 avdd.n1734 0.113554
R14876 avdd.n1734 avdd.n1733 0.113554
R14877 avdd.n1777 avdd.n1763 0.0934054
R14878 avdd.n719 avdd.n711 0.0815811
R14879 avdd.n967 avdd.n731 0.0815811
R14880 avdd.n960 avdd.n736 0.0815811
R14881 avdd.n949 avdd.n743 0.0815811
R14882 avdd.n939 avdd.n752 0.0815811
R14883 avdd.n935 avdd.n755 0.0815811
R14884 avdd.n924 avdd.n763 0.0815811
R14885 avdd.n914 avdd.n772 0.0815811
R14886 avdd.n910 avdd.n775 0.0815811
R14887 avdd.n899 avdd.n783 0.0815811
R14888 avdd.n889 avdd.n792 0.0815811
R14889 avdd.n885 avdd.n795 0.0815811
R14890 avdd.n874 avdd.n803 0.0815811
R14891 avdd.n864 avdd.n812 0.0815811
R14892 avdd.n860 avdd.n815 0.0815811
R14893 avdd.n849 avdd.n823 0.0815811
R14894 avdd.n839 avdd.n832 0.0815811
R14895 avdd.n1853 avdd.n730 0.0793136
R14896 avdd.n975 avdd.n725 0.0793136
R14897 avdd.n1058 avdd.n1057 0.0766719
R14898 avdd.n1304 avdd.n1303 0.0766719
R14899 avdd.n1471 avdd.n1470 0.076587
R14900 avdd.n1494 avdd 0.0697568
R14901 avdd.n975 avdd.n974 0.0694655
R14902 avdd.n1188 avdd.n992 0.0674065
R14903 avdd.n1610 avdd.n1238 0.0674065
R14904 avdd.n1197 avdd.n1012 0.0669286
R14905 avdd.n1065 avdd.n999 0.0669286
R14906 avdd.n1619 avdd.n1258 0.0669286
R14907 avdd.n1311 avdd.n1245 0.0669286
R14908 avdd.n1057 avdd.n1054 0.0650833
R14909 avdd.n1048 avdd.n1047 0.0650833
R14910 avdd.n1303 avdd.n1300 0.0650833
R14911 avdd.n1294 avdd.n1293 0.0650833
R14912 avdd.n16 avdd.n9 0.0579519
R14913 avdd.n348 avdd.n346 0.0579519
R14914 avdd.n320 avdd.n318 0.0579519
R14915 avdd.n292 avdd.n290 0.0579519
R14916 avdd.n264 avdd.n262 0.0579519
R14917 avdd.n236 avdd.n234 0.0579519
R14918 avdd.n208 avdd.n206 0.0579519
R14919 avdd.n180 avdd.n178 0.0579519
R14920 avdd.n152 avdd.n150 0.0579519
R14921 avdd.n121 avdd.n117 0.0579519
R14922 avdd.n685 avdd.n683 0.0579519
R14923 avdd.n657 avdd.n655 0.0579519
R14924 avdd.n629 avdd.n627 0.0579519
R14925 avdd.n601 avdd.n599 0.0579519
R14926 avdd.n573 avdd.n571 0.0579519
R14927 avdd.n545 avdd.n543 0.0579519
R14928 avdd.n517 avdd.n515 0.0579519
R14929 avdd.n489 avdd.n487 0.0579519
R14930 avdd.n458 avdd.n454 0.0579519
R14931 avdd.n1470 avdd.n1323 0.057547
R14932 avdd.n720 avdd.n710 0.0553986
R14933 avdd.n963 avdd.n735 0.0553986
R14934 avdd.n952 avdd.n742 0.0553986
R14935 avdd.n749 avdd.n748 0.0553986
R14936 avdd.n938 avdd.n754 0.0553986
R14937 avdd.n927 avdd.n762 0.0553986
R14938 avdd.n769 avdd.n768 0.0553986
R14939 avdd.n913 avdd.n774 0.0553986
R14940 avdd.n902 avdd.n782 0.0553986
R14941 avdd.n789 avdd.n788 0.0553986
R14942 avdd.n888 avdd.n794 0.0553986
R14943 avdd.n877 avdd.n802 0.0553986
R14944 avdd.n809 avdd.n808 0.0553986
R14945 avdd.n863 avdd.n814 0.0553986
R14946 avdd.n852 avdd.n822 0.0553986
R14947 avdd.n829 avdd.n828 0.0553986
R14948 avdd.n838 avdd.n835 0.0553986
R14949 avdd.n1698 avdd.n1697 0.0527472
R14950 avdd.n1496 avdd.n1492 0.0516745
R14951 avdd.n1696 avdd.n1695 0.0510435
R14952 avdd.n1677 avdd.n1673 0.0507703
R14953 avdd.n1754 avdd.n1752 0.0489375
R14954 avdd.n1780 avdd.n1753 0.0489375
R14955 avdd.n1693 avdd.n1692 0.0467687
R14956 avdd avdd.n1863 0.04675
R14957 avdd.n1492 avdd 0.0441242
R14958 avdd.n1738 avdd.n1737 0.0436892
R14959 avdd.n1849 avdd.n1818 0.0430541
R14960 avdd.n1743 avdd.n1732 0.0430541
R14961 avdd.n711 avdd 0.0410405
R14962 avdd avdd.n18 0.04
R14963 avdd avdd.n123 0.04
R14964 avdd avdd.n157 0.04
R14965 avdd avdd.n185 0.04
R14966 avdd avdd.n213 0.04
R14967 avdd avdd.n241 0.04
R14968 avdd avdd.n269 0.04
R14969 avdd avdd.n297 0.04
R14970 avdd avdd.n325 0.04
R14971 avdd avdd.n353 0.04
R14972 avdd avdd.n460 0.04
R14973 avdd avdd.n494 0.04
R14974 avdd avdd.n522 0.04
R14975 avdd avdd.n550 0.04
R14976 avdd avdd.n578 0.04
R14977 avdd avdd.n606 0.04
R14978 avdd avdd.n634 0.04
R14979 avdd avdd.n662 0.04
R14980 avdd avdd.n690 0.04
R14981 avdd.n1656 avdd.n986 0.0375
R14982 avdd avdd.n14 0.0365
R14983 avdd avdd.n119 0.0365
R14984 avdd avdd.n148 0.0365
R14985 avdd avdd.n176 0.0365
R14986 avdd avdd.n204 0.0365
R14987 avdd avdd.n232 0.0365
R14988 avdd avdd.n260 0.0365
R14989 avdd avdd.n288 0.0365
R14990 avdd avdd.n316 0.0365
R14991 avdd avdd.n344 0.0365
R14992 avdd avdd.n456 0.0365
R14993 avdd avdd.n485 0.0365
R14994 avdd avdd.n513 0.0365
R14995 avdd avdd.n541 0.0365
R14996 avdd avdd.n569 0.0365
R14997 avdd avdd.n597 0.0365
R14998 avdd avdd.n625 0.0365
R14999 avdd avdd.n653 0.0365
R15000 avdd avdd.n681 0.0365
R15001 avdd.n962 avdd 0.0351284
R15002 avdd.n951 avdd 0.0351284
R15003 avdd avdd.n751 0.0351284
R15004 avdd.n936 avdd 0.0351284
R15005 avdd.n926 avdd 0.0351284
R15006 avdd avdd.n771 0.0351284
R15007 avdd.n911 avdd 0.0351284
R15008 avdd.n901 avdd 0.0351284
R15009 avdd avdd.n791 0.0351284
R15010 avdd.n886 avdd 0.0351284
R15011 avdd.n876 avdd 0.0351284
R15012 avdd avdd.n811 0.0351284
R15013 avdd.n861 avdd 0.0351284
R15014 avdd.n851 avdd 0.0351284
R15015 avdd avdd.n831 0.0351284
R15016 avdd.n836 avdd 0.0351284
R15017 avdd.n108 avdd 0.0335784
R15018 avdd.n445 avdd 0.0335784
R15019 avdd.n27 avdd 0.032
R15020 avdd.n139 avdd 0.032
R15021 avdd.n167 avdd 0.032
R15022 avdd.n195 avdd 0.032
R15023 avdd.n223 avdd 0.032
R15024 avdd.n251 avdd 0.032
R15025 avdd.n279 avdd 0.032
R15026 avdd.n307 avdd 0.032
R15027 avdd.n335 avdd 0.032
R15028 avdd.n363 avdd 0.032
R15029 avdd.n476 avdd 0.032
R15030 avdd.n504 avdd 0.032
R15031 avdd.n532 avdd 0.032
R15032 avdd.n560 avdd 0.032
R15033 avdd.n588 avdd 0.032
R15034 avdd.n616 avdd 0.032
R15035 avdd.n644 avdd 0.032
R15036 avdd.n672 avdd 0.032
R15037 avdd.n700 avdd 0.032
R15038 avdd.n1672 avdd.n1666 0.0301178
R15039 avdd.n1676 avdd.n1675 0.0300238
R15040 avdd.n1733 avdd.n1716 0.0287635
R15041 avdd.n1709 avdd.n1708 0.0283443
R15042 avdd.n114 avdd 0.028
R15043 avdd.n451 avdd 0.028
R15044 avdd.n720 avdd.n719 0.0266824
R15045 avdd.n735 avdd.n731 0.0266824
R15046 avdd.n742 avdd.n736 0.0266824
R15047 avdd.n749 avdd.n743 0.0266824
R15048 avdd.n939 avdd.n938 0.0266824
R15049 avdd.n762 avdd.n755 0.0266824
R15050 avdd.n769 avdd.n763 0.0266824
R15051 avdd.n914 avdd.n913 0.0266824
R15052 avdd.n782 avdd.n775 0.0266824
R15053 avdd.n789 avdd.n783 0.0266824
R15054 avdd.n889 avdd.n888 0.0266824
R15055 avdd.n802 avdd.n795 0.0266824
R15056 avdd.n809 avdd.n803 0.0266824
R15057 avdd.n864 avdd.n863 0.0266824
R15058 avdd.n822 avdd.n815 0.0266824
R15059 avdd.n829 avdd.n823 0.0266824
R15060 avdd.n839 avdd.n838 0.0266824
R15061 avdd.n13 avdd 0.0245
R15062 avdd.n124 avdd 0.0245
R15063 avdd.n118 avdd 0.0245
R15064 avdd avdd.n158 0.0245
R15065 avdd.n154 avdd 0.0245
R15066 avdd avdd.n186 0.0245
R15067 avdd.n182 avdd 0.0245
R15068 avdd avdd.n214 0.0245
R15069 avdd.n210 avdd 0.0245
R15070 avdd avdd.n242 0.0245
R15071 avdd.n238 avdd 0.0245
R15072 avdd avdd.n270 0.0245
R15073 avdd.n266 avdd 0.0245
R15074 avdd avdd.n298 0.0245
R15075 avdd.n294 avdd 0.0245
R15076 avdd avdd.n326 0.0245
R15077 avdd.n322 avdd 0.0245
R15078 avdd avdd.n354 0.0245
R15079 avdd.n350 avdd 0.0245
R15080 avdd.n455 avdd 0.0245
R15081 avdd avdd.n495 0.0245
R15082 avdd.n491 avdd 0.0245
R15083 avdd avdd.n523 0.0245
R15084 avdd.n519 avdd 0.0245
R15085 avdd avdd.n551 0.0245
R15086 avdd.n547 avdd 0.0245
R15087 avdd avdd.n579 0.0245
R15088 avdd.n575 avdd 0.0245
R15089 avdd avdd.n607 0.0245
R15090 avdd.n603 avdd 0.0245
R15091 avdd avdd.n635 0.0245
R15092 avdd.n631 avdd 0.0245
R15093 avdd avdd.n663 0.0245
R15094 avdd.n659 avdd 0.0245
R15095 avdd avdd.n691 0.0245
R15096 avdd.n687 avdd 0.0245
R15097 avdd.n1694 avdd.n1664 0.0240443
R15098 avdd.n461 avdd 0.024
R15099 avdd.n19 avdd.n7 0.0235
R15100 avdd.n1494 avdd.n1492 0.0190811
R15101 avdd.n1497 avdd.n1496 0.0164396
R15102 avdd avdd.n108 0.0163924
R15103 avdd avdd.n445 0.0163924
R15104 avdd avdd.n1232 0.01225
R15105 avdd avdd.n1654 0.01225
R15106 avdd avdd.n0 0.012
R15107 avdd avdd.n98 0.012
R15108 avdd avdd.n90 0.012
R15109 avdd avdd.n82 0.012
R15110 avdd avdd.n74 0.012
R15111 avdd avdd.n66 0.012
R15112 avdd avdd.n58 0.012
R15113 avdd avdd.n50 0.012
R15114 avdd avdd.n42 0.012
R15115 avdd avdd.n34 0.012
R15116 avdd avdd.n435 0.012
R15117 avdd avdd.n427 0.012
R15118 avdd avdd.n419 0.012
R15119 avdd avdd.n411 0.012
R15120 avdd avdd.n403 0.012
R15121 avdd avdd.n395 0.012
R15122 avdd avdd.n387 0.012
R15123 avdd avdd.n379 0.012
R15124 avdd avdd.n371 0.012
R15125 avdd.n1492 avdd.n1491 0.0113696
R15126 avdd.n1497 avdd.n1323 0.0105671
R15127 avdd.n19 avdd 0.009
R15128 avdd.n18 avdd 0.009
R15129 avdd.n17 avdd 0.009
R15130 avdd.n14 avdd 0.009
R15131 avdd.n31 avdd 0.009
R15132 avdd.n31 avdd 0.009
R15133 avdd.n30 avdd 0.009
R15134 avdd avdd.n111 0.009
R15135 avdd.n112 avdd 0.009
R15136 avdd.n124 avdd 0.009
R15137 avdd.n123 avdd 0.009
R15138 avdd.n122 avdd 0.009
R15139 avdd.n119 avdd 0.009
R15140 avdd.n143 avdd 0.009
R15141 avdd.n143 avdd 0.009
R15142 avdd.n142 avdd 0.009
R15143 avdd.n159 avdd 0.009
R15144 avdd.n158 avdd 0.009
R15145 avdd.n157 avdd 0.009
R15146 avdd.n151 avdd 0.009
R15147 avdd.n148 avdd 0.009
R15148 avdd.n171 avdd 0.009
R15149 avdd.n171 avdd 0.009
R15150 avdd.n170 avdd 0.009
R15151 avdd.n187 avdd 0.009
R15152 avdd.n186 avdd 0.009
R15153 avdd.n185 avdd 0.009
R15154 avdd.n179 avdd 0.009
R15155 avdd.n176 avdd 0.009
R15156 avdd.n199 avdd 0.009
R15157 avdd.n199 avdd 0.009
R15158 avdd.n198 avdd 0.009
R15159 avdd.n215 avdd 0.009
R15160 avdd.n214 avdd 0.009
R15161 avdd.n213 avdd 0.009
R15162 avdd.n207 avdd 0.009
R15163 avdd.n204 avdd 0.009
R15164 avdd.n227 avdd 0.009
R15165 avdd.n227 avdd 0.009
R15166 avdd.n226 avdd 0.009
R15167 avdd.n243 avdd 0.009
R15168 avdd.n242 avdd 0.009
R15169 avdd.n241 avdd 0.009
R15170 avdd.n235 avdd 0.009
R15171 avdd.n232 avdd 0.009
R15172 avdd.n255 avdd 0.009
R15173 avdd.n255 avdd 0.009
R15174 avdd.n254 avdd 0.009
R15175 avdd.n271 avdd 0.009
R15176 avdd.n270 avdd 0.009
R15177 avdd.n269 avdd 0.009
R15178 avdd.n263 avdd 0.009
R15179 avdd.n260 avdd 0.009
R15180 avdd.n283 avdd 0.009
R15181 avdd.n283 avdd 0.009
R15182 avdd.n282 avdd 0.009
R15183 avdd.n299 avdd 0.009
R15184 avdd.n298 avdd 0.009
R15185 avdd.n297 avdd 0.009
R15186 avdd.n291 avdd 0.009
R15187 avdd.n288 avdd 0.009
R15188 avdd.n311 avdd 0.009
R15189 avdd.n311 avdd 0.009
R15190 avdd.n310 avdd 0.009
R15191 avdd.n327 avdd 0.009
R15192 avdd.n326 avdd 0.009
R15193 avdd.n325 avdd 0.009
R15194 avdd.n319 avdd 0.009
R15195 avdd.n316 avdd 0.009
R15196 avdd.n339 avdd 0.009
R15197 avdd.n339 avdd 0.009
R15198 avdd.n338 avdd 0.009
R15199 avdd.n355 avdd 0.009
R15200 avdd.n354 avdd 0.009
R15201 avdd.n353 avdd 0.009
R15202 avdd.n347 avdd 0.009
R15203 avdd.n344 avdd 0.009
R15204 avdd.n367 avdd 0.009
R15205 avdd.n367 avdd 0.009
R15206 avdd.n366 avdd 0.009
R15207 avdd avdd.n448 0.009
R15208 avdd.n449 avdd 0.009
R15209 avdd.n461 avdd 0.009
R15210 avdd.n460 avdd 0.009
R15211 avdd.n459 avdd 0.009
R15212 avdd.n456 avdd 0.009
R15213 avdd.n480 avdd 0.009
R15214 avdd.n480 avdd 0.009
R15215 avdd.n479 avdd 0.009
R15216 avdd.n496 avdd 0.009
R15217 avdd.n495 avdd 0.009
R15218 avdd.n494 avdd 0.009
R15219 avdd.n488 avdd 0.009
R15220 avdd.n485 avdd 0.009
R15221 avdd.n508 avdd 0.009
R15222 avdd.n508 avdd 0.009
R15223 avdd.n507 avdd 0.009
R15224 avdd.n524 avdd 0.009
R15225 avdd.n523 avdd 0.009
R15226 avdd.n522 avdd 0.009
R15227 avdd.n516 avdd 0.009
R15228 avdd.n513 avdd 0.009
R15229 avdd.n536 avdd 0.009
R15230 avdd.n536 avdd 0.009
R15231 avdd.n535 avdd 0.009
R15232 avdd.n552 avdd 0.009
R15233 avdd.n551 avdd 0.009
R15234 avdd.n550 avdd 0.009
R15235 avdd.n544 avdd 0.009
R15236 avdd.n541 avdd 0.009
R15237 avdd.n564 avdd 0.009
R15238 avdd.n564 avdd 0.009
R15239 avdd.n563 avdd 0.009
R15240 avdd.n580 avdd 0.009
R15241 avdd.n579 avdd 0.009
R15242 avdd.n578 avdd 0.009
R15243 avdd.n572 avdd 0.009
R15244 avdd.n569 avdd 0.009
R15245 avdd.n592 avdd 0.009
R15246 avdd.n592 avdd 0.009
R15247 avdd.n591 avdd 0.009
R15248 avdd.n608 avdd 0.009
R15249 avdd.n607 avdd 0.009
R15250 avdd.n606 avdd 0.009
R15251 avdd.n600 avdd 0.009
R15252 avdd.n597 avdd 0.009
R15253 avdd.n620 avdd 0.009
R15254 avdd.n620 avdd 0.009
R15255 avdd.n619 avdd 0.009
R15256 avdd.n636 avdd 0.009
R15257 avdd.n635 avdd 0.009
R15258 avdd.n634 avdd 0.009
R15259 avdd.n628 avdd 0.009
R15260 avdd.n625 avdd 0.009
R15261 avdd.n648 avdd 0.009
R15262 avdd.n648 avdd 0.009
R15263 avdd.n647 avdd 0.009
R15264 avdd.n664 avdd 0.009
R15265 avdd.n663 avdd 0.009
R15266 avdd.n662 avdd 0.009
R15267 avdd.n656 avdd 0.009
R15268 avdd.n653 avdd 0.009
R15269 avdd.n676 avdd 0.009
R15270 avdd.n676 avdd 0.009
R15271 avdd.n675 avdd 0.009
R15272 avdd.n692 avdd 0.009
R15273 avdd.n691 avdd 0.009
R15274 avdd.n690 avdd 0.009
R15275 avdd.n684 avdd 0.009
R15276 avdd.n681 avdd 0.009
R15277 avdd.n704 avdd 0.009
R15278 avdd.n704 avdd 0.009
R15279 avdd.n703 avdd 0.009
R15280 avdd.n27 avdd.n26 0.0085
R15281 avdd avdd.n115 0.0085
R15282 avdd.n139 avdd.n138 0.0085
R15283 avdd.n167 avdd.n166 0.0085
R15284 avdd.n195 avdd.n194 0.0085
R15285 avdd.n223 avdd.n222 0.0085
R15286 avdd.n251 avdd.n250 0.0085
R15287 avdd.n279 avdd.n278 0.0085
R15288 avdd.n307 avdd.n306 0.0085
R15289 avdd.n335 avdd.n334 0.0085
R15290 avdd.n363 avdd.n362 0.0085
R15291 avdd avdd.n452 0.0085
R15292 avdd.n476 avdd.n475 0.0085
R15293 avdd.n504 avdd.n503 0.0085
R15294 avdd.n532 avdd.n531 0.0085
R15295 avdd.n560 avdd.n559 0.0085
R15296 avdd.n588 avdd.n587 0.0085
R15297 avdd.n616 avdd.n615 0.0085
R15298 avdd.n644 avdd.n643 0.0085
R15299 avdd.n672 avdd.n671 0.0085
R15300 avdd.n700 avdd.n699 0.0085
R15301 avdd avdd.n17 0.0075
R15302 avdd avdd.n122 0.0075
R15303 avdd.n151 avdd 0.0075
R15304 avdd.n179 avdd 0.0075
R15305 avdd.n207 avdd 0.0075
R15306 avdd.n235 avdd 0.0075
R15307 avdd.n263 avdd 0.0075
R15308 avdd.n291 avdd 0.0075
R15309 avdd.n319 avdd 0.0075
R15310 avdd.n347 avdd 0.0075
R15311 avdd avdd.n459 0.0075
R15312 avdd.n488 avdd 0.0075
R15313 avdd.n516 avdd 0.0075
R15314 avdd.n544 avdd 0.0075
R15315 avdd.n572 avdd 0.0075
R15316 avdd.n600 avdd 0.0075
R15317 avdd.n628 avdd 0.0075
R15318 avdd.n656 avdd 0.0075
R15319 avdd.n684 avdd 0.0075
R15320 avdd.n722 avdd.n710 0.00641216
R15321 avdd.n963 avdd.n962 0.00641216
R15322 avdd.n952 avdd.n951 0.00641216
R15323 avdd.n751 avdd.n748 0.00641216
R15324 avdd.n936 avdd.n754 0.00641216
R15325 avdd.n927 avdd.n926 0.00641216
R15326 avdd.n771 avdd.n768 0.00641216
R15327 avdd.n911 avdd.n774 0.00641216
R15328 avdd.n902 avdd.n901 0.00641216
R15329 avdd.n791 avdd.n788 0.00641216
R15330 avdd.n886 avdd.n794 0.00641216
R15331 avdd.n877 avdd.n876 0.00641216
R15332 avdd.n811 avdd.n808 0.00641216
R15333 avdd.n861 avdd.n814 0.00641216
R15334 avdd.n852 avdd.n851 0.00641216
R15335 avdd.n831 avdd.n828 0.00641216
R15336 avdd.n836 avdd.n835 0.00641216
R15337 avdd.n15 avdd 0.0055
R15338 avdd.n33 avdd.n0 0.0055
R15339 avdd.n120 avdd 0.0055
R15340 avdd.n145 avdd.n98 0.0055
R15341 avdd.n153 avdd 0.0055
R15342 avdd.n173 avdd.n90 0.0055
R15343 avdd.n181 avdd 0.0055
R15344 avdd.n201 avdd.n82 0.0055
R15345 avdd.n209 avdd 0.0055
R15346 avdd.n229 avdd.n74 0.0055
R15347 avdd.n237 avdd 0.0055
R15348 avdd.n257 avdd.n66 0.0055
R15349 avdd.n265 avdd 0.0055
R15350 avdd.n285 avdd.n58 0.0055
R15351 avdd.n293 avdd 0.0055
R15352 avdd.n313 avdd.n50 0.0055
R15353 avdd.n321 avdd 0.0055
R15354 avdd.n341 avdd.n42 0.0055
R15355 avdd.n349 avdd 0.0055
R15356 avdd.n369 avdd.n34 0.0055
R15357 avdd.n457 avdd 0.0055
R15358 avdd.n482 avdd.n435 0.0055
R15359 avdd.n490 avdd 0.0055
R15360 avdd.n510 avdd.n427 0.0055
R15361 avdd.n518 avdd 0.0055
R15362 avdd.n538 avdd.n419 0.0055
R15363 avdd.n546 avdd 0.0055
R15364 avdd.n566 avdd.n411 0.0055
R15365 avdd.n574 avdd 0.0055
R15366 avdd.n594 avdd.n403 0.0055
R15367 avdd.n602 avdd 0.0055
R15368 avdd.n622 avdd.n395 0.0055
R15369 avdd.n630 avdd 0.0055
R15370 avdd.n650 avdd.n387 0.0055
R15371 avdd.n658 avdd 0.0055
R15372 avdd.n678 avdd.n379 0.0055
R15373 avdd.n686 avdd 0.0055
R15374 avdd.n706 avdd.n371 0.0055
R15375 avdd.n15 avdd.n13 0.004
R15376 avdd avdd.n33 0.004
R15377 avdd.n120 avdd.n118 0.004
R15378 avdd avdd.n145 0.004
R15379 avdd.n154 avdd.n153 0.004
R15380 avdd avdd.n173 0.004
R15381 avdd.n182 avdd.n181 0.004
R15382 avdd avdd.n201 0.004
R15383 avdd.n210 avdd.n209 0.004
R15384 avdd avdd.n229 0.004
R15385 avdd.n238 avdd.n237 0.004
R15386 avdd avdd.n257 0.004
R15387 avdd.n266 avdd.n265 0.004
R15388 avdd avdd.n285 0.004
R15389 avdd.n294 avdd.n293 0.004
R15390 avdd avdd.n313 0.004
R15391 avdd.n322 avdd.n321 0.004
R15392 avdd avdd.n341 0.004
R15393 avdd.n350 avdd.n349 0.004
R15394 avdd avdd.n369 0.004
R15395 avdd.n457 avdd.n455 0.004
R15396 avdd avdd.n482 0.004
R15397 avdd.n491 avdd.n490 0.004
R15398 avdd avdd.n510 0.004
R15399 avdd.n519 avdd.n518 0.004
R15400 avdd avdd.n538 0.004
R15401 avdd.n547 avdd.n546 0.004
R15402 avdd avdd.n566 0.004
R15403 avdd.n575 avdd.n574 0.004
R15404 avdd avdd.n594 0.004
R15405 avdd.n603 avdd.n602 0.004
R15406 avdd avdd.n622 0.004
R15407 avdd.n631 avdd.n630 0.004
R15408 avdd avdd.n650 0.004
R15409 avdd.n659 avdd.n658 0.004
R15410 avdd avdd.n678 0.004
R15411 avdd.n687 avdd.n686 0.004
R15412 avdd avdd.n706 0.004
R15413 avdd.n112 avdd 0.0035
R15414 avdd.n449 avdd 0.0035
R15415 avdd avdd.n30 0.003
R15416 avdd avdd.n142 0.003
R15417 avdd avdd.n170 0.003
R15418 avdd avdd.n198 0.003
R15419 avdd avdd.n226 0.003
R15420 avdd avdd.n254 0.003
R15421 avdd avdd.n282 0.003
R15422 avdd avdd.n310 0.003
R15423 avdd avdd.n338 0.003
R15424 avdd avdd.n366 0.003
R15425 avdd avdd.n479 0.003
R15426 avdd avdd.n507 0.003
R15427 avdd avdd.n535 0.003
R15428 avdd avdd.n563 0.003
R15429 avdd avdd.n591 0.003
R15430 avdd avdd.n619 0.003
R15431 avdd avdd.n647 0.003
R15432 avdd avdd.n675 0.003
R15433 avdd avdd.n703 0.003
R15434 avdd.n26 avdd 0.001
R15435 avdd.n115 avdd.n114 0.001
R15436 avdd.n138 avdd 0.001
R15437 avdd.n166 avdd 0.001
R15438 avdd.n194 avdd 0.001
R15439 avdd.n222 avdd 0.001
R15440 avdd.n250 avdd 0.001
R15441 avdd.n278 avdd 0.001
R15442 avdd.n306 avdd 0.001
R15443 avdd.n334 avdd 0.001
R15444 avdd.n362 avdd 0.001
R15445 avdd.n452 avdd.n451 0.001
R15446 avdd.n475 avdd 0.001
R15447 avdd.n503 avdd 0.001
R15448 avdd.n531 avdd 0.001
R15449 avdd.n559 avdd 0.001
R15450 avdd.n587 avdd 0.001
R15451 avdd.n615 avdd 0.001
R15452 avdd.n643 avdd 0.001
R15453 avdd.n671 avdd 0.001
R15454 avdd.n699 avdd 0.001
R15455 porb.n2 porb.n0 243.458
R15456 porb.n2 porb.n1 205.059
R15457 porb.n4 porb.n3 205.059
R15458 porb.n6 porb.n5 205.059
R15459 porb.n8 porb.n7 205.059
R15460 porb.n10 porb.n9 205.059
R15461 porb.n12 porb.n11 205.059
R15462 porb.n14 porb.n13 205.059
R15463 porb.n17 porb.n15 133.534
R15464 porb.n17 porb.n16 99.1759
R15465 porb.n19 porb.n18 99.1759
R15466 porb.n21 porb.n20 99.1759
R15467 porb.n23 porb.n22 99.1759
R15468 porb.n25 porb.n24 99.1759
R15469 porb.n27 porb.n26 99.1759
R15470 porb porb.n28 97.4305
R15471 porb.n4 porb.n2 38.4005
R15472 porb.n6 porb.n4 38.4005
R15473 porb.n8 porb.n6 38.4005
R15474 porb.n10 porb.n8 38.4005
R15475 porb.n12 porb.n10 38.4005
R15476 porb.n14 porb.n12 38.4005
R15477 porb.n19 porb.n17 34.3584
R15478 porb.n21 porb.n19 34.3584
R15479 porb.n23 porb.n21 34.3584
R15480 porb.n25 porb.n23 34.3584
R15481 porb.n27 porb.n25 34.3584
R15482 porb.n29 porb.n27 34.3584
R15483 porb.n13 porb.t17 26.5955
R15484 porb.n13 porb.t22 26.5955
R15485 porb.n0 porb.t31 26.5955
R15486 porb.n0 porb.t26 26.5955
R15487 porb.n1 porb.t30 26.5955
R15488 porb.n1 porb.t24 26.5955
R15489 porb.n3 porb.t21 26.5955
R15490 porb.n3 porb.t23 26.5955
R15491 porb.n5 porb.t20 26.5955
R15492 porb.n5 porb.t28 26.5955
R15493 porb.n7 porb.t16 26.5955
R15494 porb.n7 porb.t27 26.5955
R15495 porb.n9 porb.t19 26.5955
R15496 porb.n9 porb.t25 26.5955
R15497 porb.n11 porb.t18 26.5955
R15498 porb.n11 porb.t29 26.5955
R15499 porb.n28 porb.t13 24.9236
R15500 porb.n28 porb.t2 24.9236
R15501 porb.n15 porb.t11 24.9236
R15502 porb.n15 porb.t6 24.9236
R15503 porb.n16 porb.t10 24.9236
R15504 porb.n16 porb.t4 24.9236
R15505 porb.n18 porb.t1 24.9236
R15506 porb.n18 porb.t3 24.9236
R15507 porb.n20 porb.t0 24.9236
R15508 porb.n20 porb.t8 24.9236
R15509 porb.n22 porb.t12 24.9236
R15510 porb.n22 porb.t7 24.9236
R15511 porb.n24 porb.t15 24.9236
R15512 porb.n24 porb.t5 24.9236
R15513 porb.n26 porb.t14 24.9236
R15514 porb.n26 porb.t9 24.9236
R15515 porb porb.n14 18.4247
R15516 porb.n30 porb.n29 8.33989
R15517 porb.n30 porb 4.78765
R15518 porb porb.n30 3.10353
R15519 porb.n29 porb 1.74595
R15520 dvdd.n481 dvdd.n479 53399.3
R15521 dvdd.n483 dvdd.n479 53399.3
R15522 dvdd.n483 dvdd.n482 53399.3
R15523 dvdd.n482 dvdd.n481 53399.3
R15524 dvdd.n480 dvdd.n478 26464.9
R15525 dvdd.n484 dvdd.n478 26464.9
R15526 dvdd.n484 dvdd.n477 26464.9
R15527 dvdd.n480 dvdd.n477 26464.9
R15528 dvdd.n284 dvdd.n282 15977.3
R15529 dvdd.n286 dvdd.n282 15974
R15530 dvdd.n285 dvdd.n284 15974
R15531 dvdd.n286 dvdd.n285 15970.6
R15532 dvdd.n513 dvdd.n510 8474.12
R15533 dvdd.n515 dvdd.n510 8474.12
R15534 dvdd.n513 dvdd.n512 8470.59
R15535 dvdd.n515 dvdd.n512 8470.59
R15536 dvdd.n283 dvdd.n280 8195.68
R15537 dvdd.n283 dvdd.n281 8194.05
R15538 dvdd.n287 dvdd.n280 8194.05
R15539 dvdd.n287 dvdd.n281 8192.43
R15540 dvdd.n476 dvdd.n475 6151.53
R15541 dvdd.n486 dvdd.n476 6151.53
R15542 dvdd.n485 dvdd.n475 6151.53
R15543 dvdd.n486 dvdd.n485 6151.53
R15544 dvdd.n215 dvdd.n214 4782.35
R15545 dvdd.n216 dvdd.n214 4782.35
R15546 dvdd.n215 dvdd.n199 4782.35
R15547 dvdd.n216 dvdd.n199 4782.35
R15548 dvdd.n289 dvdd.n279 1910.21
R15549 dvdd.n279 dvdd.n278 1909.84
R15550 dvdd.n289 dvdd.n288 1909.84
R15551 dvdd.n288 dvdd.n278 1909.46
R15552 dvdd.n518 dvdd.n509 903.907
R15553 dvdd.n516 dvdd.n511 903.529
R15554 dvdd.n511 dvdd.n509 903.529
R15555 dvdd.n269 dvdd.t61 871.962
R15556 dvdd.n129 dvdd.t203 871.962
R15557 dvdd.n186 dvdd.t241 871.962
R15558 dvdd.n353 dvdd.t201 871.962
R15559 dvdd.n299 dvdd.t227 871.962
R15560 dvdd.n517 dvdd.n516 857.977
R15561 dvdd.n217 dvdd.n213 510.118
R15562 dvdd.n218 dvdd.n217 510.118
R15563 dvdd.n218 dvdd.n198 510.118
R15564 dvdd.n213 dvdd.n198 510.118
R15565 dvdd.t96 dvdd.n215 369.05
R15566 dvdd.n216 dvdd.t90 369.05
R15567 dvdd.n499 dvdd.t323 360.925
R15568 dvdd.n497 dvdd.t313 360.795
R15569 dvdd dvdd.t226 350
R15570 dvdd dvdd.t200 350
R15571 dvdd.n311 dvdd.t143 349.238
R15572 dvdd.n236 dvdd.t17 348.805
R15573 dvdd.n96 dvdd.t273 348.755
R15574 dvdd.n153 dvdd.t302 348.755
R15575 dvdd dvdd.t202 341.488
R15576 dvdd dvdd.t240 341.488
R15577 dvdd dvdd.t60 336.933
R15578 dvdd.n274 dvdd.n223 320.976
R15579 dvdd.n263 dvdd.n227 320.976
R15580 dvdd.n229 dvdd.n228 320.976
R15581 dvdd.n255 dvdd.n231 320.976
R15582 dvdd.n249 dvdd.n248 320.976
R15583 dvdd.n246 dvdd.n234 320.976
R15584 dvdd.n240 dvdd.n239 320.976
R15585 dvdd.n238 dvdd.n237 320.976
R15586 dvdd.n134 dvdd.n83 320.976
R15587 dvdd.n123 dvdd.n87 320.976
R15588 dvdd.n89 dvdd.n88 320.976
R15589 dvdd.n115 dvdd.n91 320.976
R15590 dvdd.n109 dvdd.n108 320.976
R15591 dvdd.n106 dvdd.n94 320.976
R15592 dvdd.n100 dvdd.n99 320.976
R15593 dvdd.n98 dvdd.n97 320.976
R15594 dvdd.n191 dvdd.n140 320.976
R15595 dvdd.n180 dvdd.n144 320.976
R15596 dvdd.n146 dvdd.n145 320.976
R15597 dvdd.n172 dvdd.n148 320.976
R15598 dvdd.n166 dvdd.n165 320.976
R15599 dvdd.n163 dvdd.n151 320.976
R15600 dvdd.n157 dvdd.n156 320.976
R15601 dvdd.n155 dvdd.n154 320.976
R15602 dvdd.n348 dvdd.n298 320.976
R15603 dvdd.n358 dvdd.n294 320.976
R15604 dvdd.n338 dvdd.n302 320.976
R15605 dvdd.n304 dvdd.n303 320.976
R15606 dvdd.n330 dvdd.n306 320.976
R15607 dvdd.n324 dvdd.n323 320.976
R15608 dvdd.n321 dvdd.n309 320.976
R15609 dvdd.n315 dvdd.n314 320.976
R15610 dvdd.n313 dvdd.n312 320.976
R15611 dvdd.n80 dvdd.n72 307.762
R15612 dvdd.n469 dvdd.n363 307.762
R15613 dvdd.n465 dvdd.n370 307.762
R15614 dvdd.n461 dvdd.n377 307.762
R15615 dvdd.n457 dvdd.n384 307.762
R15616 dvdd.n453 dvdd.n391 307.762
R15617 dvdd.n449 dvdd.n398 307.762
R15618 dvdd.n445 dvdd.n405 307.762
R15619 dvdd.n441 dvdd.n412 307.762
R15620 dvdd.n437 dvdd.n419 307.762
R15621 dvdd.n528 dvdd.n71 307.762
R15622 dvdd.n532 dvdd.n64 307.762
R15623 dvdd.n536 dvdd.n57 307.762
R15624 dvdd.n540 dvdd.n50 307.762
R15625 dvdd.n544 dvdd.n43 307.762
R15626 dvdd.n548 dvdd.n36 307.762
R15627 dvdd.n552 dvdd.n29 307.762
R15628 dvdd.n556 dvdd.n22 307.762
R15629 dvdd.n560 dvdd.n15 307.762
R15630 dvdd.t94 dvdd.t96 264.262
R15631 dvdd.t98 dvdd.t94 264.262
R15632 dvdd.t319 dvdd.t98 264.262
R15633 dvdd.t62 dvdd.t319 264.262
R15634 dvdd.t54 dvdd.t62 264.262
R15635 dvdd.t52 dvdd.t54 264.262
R15636 dvdd.t74 dvdd.t52 264.262
R15637 dvdd.t78 dvdd.t74 264.262
R15638 dvdd.t92 dvdd.t78 264.262
R15639 dvdd.t72 dvdd.t92 264.262
R15640 dvdd.t76 dvdd.t72 264.262
R15641 dvdd.t90 dvdd.t76 264.262
R15642 dvdd.n225 dvdd.t27 250.785
R15643 dvdd.n85 dvdd.t251 250.785
R15644 dvdd.n142 dvdd.t312 250.785
R15645 dvdd.n300 dvdd.t161 250.785
R15646 dvdd.n431 dvdd.t67 246.106
R15647 dvdd.n5 dvdd.t280 246.106
R15648 dvdd.n276 dvdd.t57 244.737
R15649 dvdd.n136 dvdd.t195 244.737
R15650 dvdd.n193 dvdd.t237 244.737
R15651 dvdd.n360 dvdd.t191 244.737
R15652 dvdd.n296 dvdd.t225 244.737
R15653 dvdd.n492 dvdd.t321 241.409
R15654 dvdd.n505 dvdd.t316 240.538
R15655 dvdd.n197 dvdd.t318 240.488
R15656 dvdd.n196 dvdd.t91 228.669
R15657 dvdd.t180 dvdd.n513 224.668
R15658 dvdd.t182 dvdd.t174 223.429
R15659 dvdd.t176 dvdd.t182 223.429
R15660 dvdd.t152 dvdd.t142 221.054
R15661 dvdd.t144 dvdd.t152 221.054
R15662 dvdd.t166 dvdd.t144 221.054
R15663 dvdd.t146 dvdd.t166 221.054
R15664 dvdd.t158 dvdd.t146 221.054
R15665 dvdd.t140 dvdd.t158 221.054
R15666 dvdd.t162 dvdd.t140 221.054
R15667 dvdd.t148 dvdd.t162 221.054
R15668 dvdd.t164 dvdd.t148 221.054
R15669 dvdd.t150 dvdd.t164 221.054
R15670 dvdd.t154 dvdd.t150 221.054
R15671 dvdd.t168 dvdd.t154 221.054
R15672 dvdd.t156 dvdd.t170 221.054
R15673 dvdd.t170 dvdd.t160 221.054
R15674 dvdd.t226 dvdd.t222 221.054
R15675 dvdd.t222 dvdd.t228 221.054
R15676 dvdd.t228 dvdd.t224 221.054
R15677 dvdd.t200 dvdd.t192 221.054
R15678 dvdd.t192 dvdd.t204 221.054
R15679 dvdd.t204 dvdd.t190 221.054
R15680 dvdd.t252 dvdd.t272 215.677
R15681 dvdd.t242 dvdd.t252 215.677
R15682 dvdd.t254 dvdd.t242 215.677
R15683 dvdd.t266 dvdd.t254 215.677
R15684 dvdd.t258 dvdd.t266 215.677
R15685 dvdd.t260 dvdd.t258 215.677
R15686 dvdd.t248 dvdd.t260 215.677
R15687 dvdd.t270 dvdd.t248 215.677
R15688 dvdd.t244 dvdd.t270 215.677
R15689 dvdd.t262 dvdd.t244 215.677
R15690 dvdd.t246 dvdd.t264 215.677
R15691 dvdd.t264 dvdd.t256 215.677
R15692 dvdd.t256 dvdd.t268 215.677
R15693 dvdd.t268 dvdd.t250 215.677
R15694 dvdd.t202 dvdd.t198 215.677
R15695 dvdd.t198 dvdd.t206 215.677
R15696 dvdd.t206 dvdd.t194 215.677
R15697 dvdd.t281 dvdd.t301 215.677
R15698 dvdd.t303 dvdd.t281 215.677
R15699 dvdd.t283 dvdd.t303 215.677
R15700 dvdd.t295 dvdd.t283 215.677
R15701 dvdd.t287 dvdd.t295 215.677
R15702 dvdd.t289 dvdd.t287 215.677
R15703 dvdd.t309 dvdd.t289 215.677
R15704 dvdd.t299 dvdd.t309 215.677
R15705 dvdd.t305 dvdd.t299 215.677
R15706 dvdd.t291 dvdd.t305 215.677
R15707 dvdd.t307 dvdd.t293 215.677
R15708 dvdd.t293 dvdd.t285 215.677
R15709 dvdd.t285 dvdd.t297 215.677
R15710 dvdd.t297 dvdd.t311 215.677
R15711 dvdd.t240 dvdd.t234 215.677
R15712 dvdd.t234 dvdd.t238 215.677
R15713 dvdd.t238 dvdd.t236 215.677
R15714 dvdd.t28 dvdd.t16 212.8
R15715 dvdd.t18 dvdd.t28 212.8
R15716 dvdd.t30 dvdd.t18 212.8
R15717 dvdd.t10 dvdd.t30 212.8
R15718 dvdd.t34 dvdd.t10 212.8
R15719 dvdd.t36 dvdd.t34 212.8
R15720 dvdd.t24 dvdd.t36 212.8
R15721 dvdd.t14 dvdd.t24 212.8
R15722 dvdd.t20 dvdd.t14 212.8
R15723 dvdd.t38 dvdd.t20 212.8
R15724 dvdd.t22 dvdd.t40 212.8
R15725 dvdd.t40 dvdd.t32 212.8
R15726 dvdd.t32 dvdd.t12 212.8
R15727 dvdd.t12 dvdd.t26 212.8
R15728 dvdd.t60 dvdd.t58 212.8
R15729 dvdd.t58 dvdd.t64 212.8
R15730 dvdd.t64 dvdd.t56 212.8
R15731 dvdd.n433 dvdd.n426 205.5
R15732 dvdd.n7 dvdd.n0 205.5
R15733 dvdd.t160 dvdd 205.263
R15734 dvdd.n494 dvdd.n488 200.31
R15735 dvdd.n503 dvdd.n500 200.31
R15736 dvdd.n502 dvdd.n501 200.31
R15737 dvdd.n493 dvdd.n489 200.31
R15738 dvdd.n491 dvdd.n490 200.31
R15739 dvdd.n473 dvdd.n472 200.31
R15740 dvdd.t250 dvdd 200.27
R15741 dvdd.t311 dvdd 200.27
R15742 dvdd.n524 dvdd.n523 200.173
R15743 dvdd.n497 dvdd.n496 200.115
R15744 dvdd.n209 dvdd.n208 200.105
R15745 dvdd.n210 dvdd.n207 200.105
R15746 dvdd.n211 dvdd.n206 200.105
R15747 dvdd.n205 dvdd.n200 200.105
R15748 dvdd.n204 dvdd.n201 200.105
R15749 dvdd.n203 dvdd.n202 200.105
R15750 dvdd.n497 dvdd.n495 200.095
R15751 dvdd.n499 dvdd.n498 200.034
R15752 dvdd.t26 dvdd 197.601
R15753 dvdd.t224 dvdd 197.369
R15754 dvdd.t190 dvdd 197.369
R15755 dvdd.t194 dvdd 192.569
R15756 dvdd.t236 dvdd 192.569
R15757 dvdd.t56 dvdd 190
R15758 dvdd.n77 dvdd.n74 185
R15759 dvdd.n74 dvdd.n73 185
R15760 dvdd.n367 dvdd.n364 185
R15761 dvdd.n368 dvdd.n367 185
R15762 dvdd.n374 dvdd.n371 185
R15763 dvdd.n375 dvdd.n374 185
R15764 dvdd.n381 dvdd.n378 185
R15765 dvdd.n382 dvdd.n381 185
R15766 dvdd.n388 dvdd.n385 185
R15767 dvdd.n389 dvdd.n388 185
R15768 dvdd.n395 dvdd.n392 185
R15769 dvdd.n396 dvdd.n395 185
R15770 dvdd.n402 dvdd.n399 185
R15771 dvdd.n403 dvdd.n402 185
R15772 dvdd.n409 dvdd.n406 185
R15773 dvdd.n410 dvdd.n409 185
R15774 dvdd.n416 dvdd.n413 185
R15775 dvdd.n417 dvdd.n416 185
R15776 dvdd.n423 dvdd.n420 185
R15777 dvdd.n424 dvdd.n423 185
R15778 dvdd.n68 dvdd.n65 185
R15779 dvdd.n69 dvdd.n68 185
R15780 dvdd.n61 dvdd.n58 185
R15781 dvdd.n62 dvdd.n61 185
R15782 dvdd.n54 dvdd.n51 185
R15783 dvdd.n55 dvdd.n54 185
R15784 dvdd.n47 dvdd.n44 185
R15785 dvdd.n48 dvdd.n47 185
R15786 dvdd.n40 dvdd.n37 185
R15787 dvdd.n41 dvdd.n40 185
R15788 dvdd.n33 dvdd.n30 185
R15789 dvdd.n34 dvdd.n33 185
R15790 dvdd.n26 dvdd.n23 185
R15791 dvdd.n27 dvdd.n26 185
R15792 dvdd.n19 dvdd.n16 185
R15793 dvdd.n20 dvdd.n19 185
R15794 dvdd.n12 dvdd.n9 185
R15795 dvdd.n13 dvdd.n12 185
R15796 dvdd.t174 dvdd.t322 180.129
R15797 dvdd.n515 dvdd.t138 175.306
R15798 dvdd.t214 dvdd.n514 174.066
R15799 dvdd.n336 dvdd.t168 171.054
R15800 dvdd.n430 dvdd.t66 157.446
R15801 dvdd.n4 dvdd.t278 157.446
R15802 dvdd.n117 dvdd.t246 146.351
R15803 dvdd.n174 dvdd.t307 146.351
R15804 dvdd.t136 dvdd.t317 145.488
R15805 dvdd.n257 dvdd.t22 141.868
R15806 dvdd.t178 dvdd.t180 136.828
R15807 dvdd.t184 dvdd.t178 136.828
R15808 dvdd.t44 dvdd.t184 136.828
R15809 dvdd.t46 dvdd.t44 136.828
R15810 dvdd.t48 dvdd.t46 136.828
R15811 dvdd.t322 dvdd.t48 136.828
R15812 dvdd.t216 dvdd.t214 136.828
R15813 dvdd.t212 dvdd.t216 136.828
R15814 dvdd.t218 dvdd.t212 136.828
R15815 dvdd.t208 dvdd.t218 136.828
R15816 dvdd.t210 dvdd.t208 136.828
R15817 dvdd.n75 dvdd.t172 129.546
R15818 dvdd.t232 dvdd.n366 129.546
R15819 dvdd.t81 dvdd.n373 129.546
R15820 dvdd.t122 dvdd.n380 129.546
R15821 dvdd.t230 dvdd.n387 129.546
R15822 dvdd.t130 dvdd.n394 129.546
R15823 dvdd.t8 dvdd.n401 129.546
R15824 dvdd.t120 dvdd.n408 129.546
R15825 dvdd.t220 dvdd.n415 129.546
R15826 dvdd.t83 dvdd.n422 129.546
R15827 dvdd.t274 dvdd.n67 129.546
R15828 dvdd.t124 dvdd.n60 129.546
R15829 dvdd.t128 dvdd.n53 129.546
R15830 dvdd.t118 dvdd.n46 129.546
R15831 dvdd.t42 dvdd.n39 129.546
R15832 dvdd.t132 dvdd.n32 129.546
R15833 dvdd.t88 dvdd.n25 129.546
R15834 dvdd.t126 dvdd.n18 129.546
R15835 dvdd.t50 dvdd.n11 129.546
R15836 dvdd.t85 dvdd.n427 127.638
R15837 dvdd.t276 dvdd.n1 127.638
R15838 dvdd.t314 dvdd.t136 117.776
R15839 dvdd.t324 dvdd.t210 109.983
R15840 dvdd.t317 dvdd.t80 109.983
R15841 dvdd.n78 dvdd.n73 101.644
R15842 dvdd.n369 dvdd.n364 101.644
R15843 dvdd.n376 dvdd.n371 101.644
R15844 dvdd.n383 dvdd.n378 101.644
R15845 dvdd.n390 dvdd.n385 101.644
R15846 dvdd.n397 dvdd.n392 101.644
R15847 dvdd.n404 dvdd.n399 101.644
R15848 dvdd.n411 dvdd.n406 101.644
R15849 dvdd.n418 dvdd.n413 101.644
R15850 dvdd.n425 dvdd.n420 101.644
R15851 dvdd.n70 dvdd.n65 101.644
R15852 dvdd.n63 dvdd.n58 101.644
R15853 dvdd.n56 dvdd.n51 101.644
R15854 dvdd.n49 dvdd.n44 101.644
R15855 dvdd.n42 dvdd.n37 101.644
R15856 dvdd.n35 dvdd.n30 101.644
R15857 dvdd.n28 dvdd.n23 101.644
R15858 dvdd.n21 dvdd.n16 101.644
R15859 dvdd.n14 dvdd.n9 101.644
R15860 dvdd.n432 dvdd.n427 95.8438
R15861 dvdd.n6 dvdd.n1 95.8438
R15862 dvdd.n78 dvdd.n77 92.5005
R15863 dvdd.n429 dvdd.n428 92.5005
R15864 dvdd.n369 dvdd.n368 92.5005
R15865 dvdd.n376 dvdd.n375 92.5005
R15866 dvdd.n383 dvdd.n382 92.5005
R15867 dvdd.n390 dvdd.n389 92.5005
R15868 dvdd.n397 dvdd.n396 92.5005
R15869 dvdd.n404 dvdd.n403 92.5005
R15870 dvdd.n411 dvdd.n410 92.5005
R15871 dvdd.n418 dvdd.n417 92.5005
R15872 dvdd.n425 dvdd.n424 92.5005
R15873 dvdd.n3 dvdd.n2 92.5005
R15874 dvdd.n70 dvdd.n69 92.5005
R15875 dvdd.n63 dvdd.n62 92.5005
R15876 dvdd.n56 dvdd.n55 92.5005
R15877 dvdd.n49 dvdd.n48 92.5005
R15878 dvdd.n42 dvdd.n41 92.5005
R15879 dvdd.n35 dvdd.n34 92.5005
R15880 dvdd.n28 dvdd.n27 92.5005
R15881 dvdd.n21 dvdd.n20 92.5005
R15882 dvdd.n14 dvdd.n13 92.5005
R15883 dvdd.t80 dvdd.t324 83.1363
R15884 dvdd.n429 dvdd.n427 82.3534
R15885 dvdd.n3 dvdd.n1 82.3534
R15886 dvdd.t138 dvdd.t314 78.8063
R15887 dvdd.n76 dvdd.n75 77.057
R15888 dvdd.n366 dvdd.n365 77.057
R15889 dvdd.n373 dvdd.n372 77.057
R15890 dvdd.n380 dvdd.n379 77.057
R15891 dvdd.n387 dvdd.n386 77.057
R15892 dvdd.n394 dvdd.n393 77.057
R15893 dvdd.n401 dvdd.n400 77.057
R15894 dvdd.n408 dvdd.n407 77.057
R15895 dvdd.n415 dvdd.n414 77.057
R15896 dvdd.n422 dvdd.n421 77.057
R15897 dvdd.n67 dvdd.n66 77.057
R15898 dvdd.n60 dvdd.n59 77.057
R15899 dvdd.n53 dvdd.n52 77.057
R15900 dvdd.n46 dvdd.n45 77.057
R15901 dvdd.n39 dvdd.n38 77.057
R15902 dvdd.n32 dvdd.n31 77.057
R15903 dvdd.n25 dvdd.n24 77.057
R15904 dvdd.n18 dvdd.n17 77.057
R15905 dvdd.n11 dvdd.n10 77.057
R15906 dvdd.n257 dvdd.t38 70.9338
R15907 dvdd.n117 dvdd.t262 69.3248
R15908 dvdd.n174 dvdd.t291 69.3248
R15909 dvdd.t172 dvdd.n74 67.8576
R15910 dvdd.n367 dvdd.t232 67.8576
R15911 dvdd.n374 dvdd.t81 67.8576
R15912 dvdd.n381 dvdd.t122 67.8576
R15913 dvdd.n388 dvdd.t230 67.8576
R15914 dvdd.n395 dvdd.t130 67.8576
R15915 dvdd.n402 dvdd.t8 67.8576
R15916 dvdd.n409 dvdd.t120 67.8576
R15917 dvdd.n416 dvdd.t220 67.8576
R15918 dvdd.n423 dvdd.t83 67.8576
R15919 dvdd.n68 dvdd.t274 67.8576
R15920 dvdd.n61 dvdd.t124 67.8576
R15921 dvdd.n54 dvdd.t128 67.8576
R15922 dvdd.n47 dvdd.t118 67.8576
R15923 dvdd.n40 dvdd.t42 67.8576
R15924 dvdd.n33 dvdd.t132 67.8576
R15925 dvdd.n26 dvdd.t88 67.8576
R15926 dvdd.n19 dvdd.t126 67.8576
R15927 dvdd.n12 dvdd.t50 67.8576
R15928 dvdd.n428 dvdd.t85 55.9594
R15929 dvdd.n428 dvdd.t66 55.9594
R15930 dvdd.n2 dvdd.t276 55.9594
R15931 dvdd.n2 dvdd.t278 55.9594
R15932 dvdd.n336 dvdd.t156 50.0005
R15933 dvdd.n75 dvdd.t196 47.2949
R15934 dvdd.n366 dvdd.t0 47.2949
R15935 dvdd.n373 dvdd.t2 47.2949
R15936 dvdd.n380 dvdd.t4 47.2949
R15937 dvdd.n387 dvdd.t70 47.2949
R15938 dvdd.n394 dvdd.t112 47.2949
R15939 dvdd.n401 dvdd.t114 47.2949
R15940 dvdd.n408 dvdd.t106 47.2949
R15941 dvdd.n415 dvdd.t104 47.2949
R15942 dvdd.n422 dvdd.t116 47.2949
R15943 dvdd.n67 dvdd.t188 47.2949
R15944 dvdd.n60 dvdd.t186 47.2949
R15945 dvdd.n53 dvdd.t68 47.2949
R15946 dvdd.n46 dvdd.t134 47.2949
R15947 dvdd.n39 dvdd.t108 47.2949
R15948 dvdd.n32 dvdd.t110 47.2949
R15949 dvdd.n25 dvdd.t102 47.2949
R15950 dvdd.n18 dvdd.t100 47.2949
R15951 dvdd.n11 dvdd.t6 47.2949
R15952 dvdd.n217 dvdd.n216 46.2505
R15953 dvdd.n215 dvdd.n198 46.2505
R15954 dvdd.n518 dvdd.n517 45.9299
R15955 dvdd.n431 dvdd.n430 33.4807
R15956 dvdd.n5 dvdd.n4 33.4807
R15957 dvdd.n72 dvdd.t173 32.8338
R15958 dvdd.n72 dvdd.t197 32.8338
R15959 dvdd.n363 dvdd.t233 32.8338
R15960 dvdd.n363 dvdd.t1 32.8338
R15961 dvdd.n370 dvdd.t82 32.8338
R15962 dvdd.n370 dvdd.t3 32.8338
R15963 dvdd.n377 dvdd.t123 32.8338
R15964 dvdd.n377 dvdd.t5 32.8338
R15965 dvdd.n384 dvdd.t231 32.8338
R15966 dvdd.n384 dvdd.t71 32.8338
R15967 dvdd.n391 dvdd.t131 32.8338
R15968 dvdd.n391 dvdd.t113 32.8338
R15969 dvdd.n398 dvdd.t9 32.8338
R15970 dvdd.n398 dvdd.t115 32.8338
R15971 dvdd.n405 dvdd.t121 32.8338
R15972 dvdd.n405 dvdd.t107 32.8338
R15973 dvdd.n412 dvdd.t221 32.8338
R15974 dvdd.n412 dvdd.t105 32.8338
R15975 dvdd.n419 dvdd.t84 32.8338
R15976 dvdd.n419 dvdd.t117 32.8338
R15977 dvdd.n71 dvdd.t275 32.8338
R15978 dvdd.n71 dvdd.t189 32.8338
R15979 dvdd.n64 dvdd.t125 32.8338
R15980 dvdd.n64 dvdd.t187 32.8338
R15981 dvdd.n57 dvdd.t129 32.8338
R15982 dvdd.n57 dvdd.t69 32.8338
R15983 dvdd.n50 dvdd.t119 32.8338
R15984 dvdd.n50 dvdd.t135 32.8338
R15985 dvdd.n43 dvdd.t43 32.8338
R15986 dvdd.n43 dvdd.t109 32.8338
R15987 dvdd.n36 dvdd.t133 32.8338
R15988 dvdd.n36 dvdd.t111 32.8338
R15989 dvdd.n29 dvdd.t89 32.8338
R15990 dvdd.n29 dvdd.t103 32.8338
R15991 dvdd.n22 dvdd.t127 32.8338
R15992 dvdd.n22 dvdd.t101 32.8338
R15993 dvdd.n15 dvdd.t51 32.8338
R15994 dvdd.n15 dvdd.t7 32.8338
R15995 dvdd.n76 dvdd.n73 30.8889
R15996 dvdd.n77 dvdd.n76 30.8889
R15997 dvdd.n368 dvdd.n365 30.8889
R15998 dvdd.n365 dvdd.n364 30.8889
R15999 dvdd.n375 dvdd.n372 30.8889
R16000 dvdd.n372 dvdd.n371 30.8889
R16001 dvdd.n382 dvdd.n379 30.8889
R16002 dvdd.n379 dvdd.n378 30.8889
R16003 dvdd.n389 dvdd.n386 30.8889
R16004 dvdd.n386 dvdd.n385 30.8889
R16005 dvdd.n396 dvdd.n393 30.8889
R16006 dvdd.n393 dvdd.n392 30.8889
R16007 dvdd.n403 dvdd.n400 30.8889
R16008 dvdd.n400 dvdd.n399 30.8889
R16009 dvdd.n410 dvdd.n407 30.8889
R16010 dvdd.n407 dvdd.n406 30.8889
R16011 dvdd.n417 dvdd.n414 30.8889
R16012 dvdd.n414 dvdd.n413 30.8889
R16013 dvdd.n424 dvdd.n421 30.8889
R16014 dvdd.n421 dvdd.n420 30.8889
R16015 dvdd.n69 dvdd.n66 30.8889
R16016 dvdd.n66 dvdd.n65 30.8889
R16017 dvdd.n62 dvdd.n59 30.8889
R16018 dvdd.n59 dvdd.n58 30.8889
R16019 dvdd.n55 dvdd.n52 30.8889
R16020 dvdd.n52 dvdd.n51 30.8889
R16021 dvdd.n48 dvdd.n45 30.8889
R16022 dvdd.n45 dvdd.n44 30.8889
R16023 dvdd.n41 dvdd.n38 30.8889
R16024 dvdd.n38 dvdd.n37 30.8889
R16025 dvdd.n34 dvdd.n31 30.8889
R16026 dvdd.n31 dvdd.n30 30.8889
R16027 dvdd.n27 dvdd.n24 30.8889
R16028 dvdd.n24 dvdd.n23 30.8889
R16029 dvdd.n20 dvdd.n17 30.8889
R16030 dvdd.n17 dvdd.n16 30.8889
R16031 dvdd.n13 dvdd.n10 30.8889
R16032 dvdd.n10 dvdd.n9 30.8889
R16033 dvdd.n498 dvdd.t325 29.5505
R16034 dvdd.n525 dvdd.n524 29.3154
R16035 dvdd.n208 dvdd.t73 28.5655
R16036 dvdd.n208 dvdd.t77 28.5655
R16037 dvdd.n207 dvdd.t79 28.5655
R16038 dvdd.n207 dvdd.t93 28.5655
R16039 dvdd.n206 dvdd.t53 28.5655
R16040 dvdd.n206 dvdd.t75 28.5655
R16041 dvdd.n200 dvdd.t63 28.5655
R16042 dvdd.n200 dvdd.t55 28.5655
R16043 dvdd.n201 dvdd.t99 28.5655
R16044 dvdd.n201 dvdd.t320 28.5655
R16045 dvdd.n202 dvdd.t97 28.5655
R16046 dvdd.n202 dvdd.t95 28.5655
R16047 dvdd.n488 dvdd.t177 28.5655
R16048 dvdd.n488 dvdd.t215 28.5655
R16049 dvdd.n496 dvdd.t315 28.5655
R16050 dvdd.n496 dvdd.t139 28.5655
R16051 dvdd.n495 dvdd.t137 28.5655
R16052 dvdd.t315 dvdd.n495 28.5655
R16053 dvdd.n498 dvdd.t211 28.5655
R16054 dvdd.n500 dvdd.t219 28.5655
R16055 dvdd.n500 dvdd.t209 28.5655
R16056 dvdd.n501 dvdd.t217 28.5655
R16057 dvdd.n501 dvdd.t213 28.5655
R16058 dvdd.n489 dvdd.t175 28.5655
R16059 dvdd.n489 dvdd.t183 28.5655
R16060 dvdd.n490 dvdd.t47 28.5655
R16061 dvdd.n490 dvdd.t49 28.5655
R16062 dvdd.n472 dvdd.t185 28.5655
R16063 dvdd.n472 dvdd.t45 28.5655
R16064 dvdd.n523 dvdd.t181 28.5655
R16065 dvdd.n523 dvdd.t179 28.5655
R16066 dvdd.n430 dvdd.n429 27.7986
R16067 dvdd.n4 dvdd.n3 27.7986
R16068 dvdd.n223 dvdd.t59 26.5955
R16069 dvdd.n223 dvdd.t65 26.5955
R16070 dvdd.n227 dvdd.t33 26.5955
R16071 dvdd.n227 dvdd.t13 26.5955
R16072 dvdd.n228 dvdd.t23 26.5955
R16073 dvdd.n228 dvdd.t41 26.5955
R16074 dvdd.n231 dvdd.t21 26.5955
R16075 dvdd.n231 dvdd.t39 26.5955
R16076 dvdd.n248 dvdd.t25 26.5955
R16077 dvdd.n248 dvdd.t15 26.5955
R16078 dvdd.n234 dvdd.t35 26.5955
R16079 dvdd.n234 dvdd.t37 26.5955
R16080 dvdd.n239 dvdd.t31 26.5955
R16081 dvdd.n239 dvdd.t11 26.5955
R16082 dvdd.n237 dvdd.t29 26.5955
R16083 dvdd.n237 dvdd.t19 26.5955
R16084 dvdd.n83 dvdd.t199 26.5955
R16085 dvdd.n83 dvdd.t207 26.5955
R16086 dvdd.n87 dvdd.t257 26.5955
R16087 dvdd.n87 dvdd.t269 26.5955
R16088 dvdd.n88 dvdd.t247 26.5955
R16089 dvdd.n88 dvdd.t265 26.5955
R16090 dvdd.n91 dvdd.t245 26.5955
R16091 dvdd.n91 dvdd.t263 26.5955
R16092 dvdd.n108 dvdd.t249 26.5955
R16093 dvdd.n108 dvdd.t271 26.5955
R16094 dvdd.n94 dvdd.t259 26.5955
R16095 dvdd.n94 dvdd.t261 26.5955
R16096 dvdd.n99 dvdd.t255 26.5955
R16097 dvdd.n99 dvdd.t267 26.5955
R16098 dvdd.n97 dvdd.t253 26.5955
R16099 dvdd.n97 dvdd.t243 26.5955
R16100 dvdd.n140 dvdd.t235 26.5955
R16101 dvdd.n140 dvdd.t239 26.5955
R16102 dvdd.n144 dvdd.t286 26.5955
R16103 dvdd.n144 dvdd.t298 26.5955
R16104 dvdd.n145 dvdd.t308 26.5955
R16105 dvdd.n145 dvdd.t294 26.5955
R16106 dvdd.n148 dvdd.t306 26.5955
R16107 dvdd.n148 dvdd.t292 26.5955
R16108 dvdd.n165 dvdd.t310 26.5955
R16109 dvdd.n165 dvdd.t300 26.5955
R16110 dvdd.n151 dvdd.t288 26.5955
R16111 dvdd.n151 dvdd.t290 26.5955
R16112 dvdd.n156 dvdd.t284 26.5955
R16113 dvdd.n156 dvdd.t296 26.5955
R16114 dvdd.n154 dvdd.t282 26.5955
R16115 dvdd.n154 dvdd.t304 26.5955
R16116 dvdd.n298 dvdd.t223 26.5955
R16117 dvdd.n298 dvdd.t229 26.5955
R16118 dvdd.n294 dvdd.t193 26.5955
R16119 dvdd.n294 dvdd.t205 26.5955
R16120 dvdd.n302 dvdd.t157 26.5955
R16121 dvdd.n302 dvdd.t171 26.5955
R16122 dvdd.n303 dvdd.t155 26.5955
R16123 dvdd.n303 dvdd.t169 26.5955
R16124 dvdd.n306 dvdd.t165 26.5955
R16125 dvdd.n306 dvdd.t151 26.5955
R16126 dvdd.n323 dvdd.t163 26.5955
R16127 dvdd.n323 dvdd.t149 26.5955
R16128 dvdd.n309 dvdd.t159 26.5955
R16129 dvdd.n309 dvdd.t141 26.5955
R16130 dvdd.n314 dvdd.t167 26.5955
R16131 dvdd.n314 dvdd.t147 26.5955
R16132 dvdd.n312 dvdd.t153 26.5955
R16133 dvdd.n312 dvdd.t145 26.5955
R16134 dvdd.n426 dvdd.t86 24.6255
R16135 dvdd.n426 dvdd.t87 24.6255
R16136 dvdd.n0 dvdd.t277 24.6255
R16137 dvdd.n0 dvdd.t279 24.6255
R16138 dvdd.n79 dvdd 22.5644
R16139 dvdd.n468 dvdd.n467 22.5272
R16140 dvdd.n464 dvdd.n463 22.5272
R16141 dvdd.n460 dvdd.n459 22.5272
R16142 dvdd.n456 dvdd.n455 22.5272
R16143 dvdd.n452 dvdd.n451 22.5272
R16144 dvdd.n448 dvdd.n447 22.5272
R16145 dvdd.n444 dvdd.n443 22.5272
R16146 dvdd.n440 dvdd.n439 22.5272
R16147 dvdd.n436 dvdd.n435 22.5272
R16148 dvdd.n530 dvdd.n529 22.5272
R16149 dvdd.n534 dvdd.n533 22.5272
R16150 dvdd.n538 dvdd.n537 22.5272
R16151 dvdd.n542 dvdd.n541 22.5272
R16152 dvdd.n546 dvdd.n545 22.5272
R16153 dvdd.n550 dvdd.n549 22.5272
R16154 dvdd.n554 dvdd.n553 22.5272
R16155 dvdd.n558 dvdd.n557 22.5272
R16156 dvdd.n562 dvdd.n561 22.5272
R16157 dvdd.n487 dvdd.n486 19.426
R16158 dvdd.n320 dvdd.n310 18.1174
R16159 dvdd.n325 dvdd.n322 18.1174
R16160 dvdd.n329 dvdd.n307 18.1174
R16161 dvdd.n332 dvdd.n331 18.1174
R16162 dvdd.n340 dvdd.n339 18.1174
R16163 dvdd.n344 dvdd.n343 18.1174
R16164 dvdd.n348 dvdd.n347 18.1174
R16165 dvdd.n349 dvdd.n348 18.1174
R16166 dvdd.n354 dvdd.n352 18.1174
R16167 dvdd.n358 dvdd.n295 18.1174
R16168 dvdd.n359 dvdd.n358 18.1174
R16169 dvdd.n316 dvdd.n313 17.9205
R16170 dvdd.n80 dvdd.n79 17.4938
R16171 dvdd.n469 dvdd.n468 17.4938
R16172 dvdd.n465 dvdd.n464 17.4938
R16173 dvdd.n461 dvdd.n460 17.4938
R16174 dvdd.n457 dvdd.n456 17.4938
R16175 dvdd.n453 dvdd.n452 17.4938
R16176 dvdd.n449 dvdd.n448 17.4938
R16177 dvdd.n445 dvdd.n444 17.4938
R16178 dvdd.n441 dvdd.n440 17.4938
R16179 dvdd.n437 dvdd.n436 17.4938
R16180 dvdd.n529 dvdd.n528 17.4938
R16181 dvdd.n533 dvdd.n532 17.4938
R16182 dvdd.n537 dvdd.n536 17.4938
R16183 dvdd.n541 dvdd.n540 17.4938
R16184 dvdd.n545 dvdd.n544 17.4938
R16185 dvdd.n549 dvdd.n548 17.4938
R16186 dvdd.n553 dvdd.n552 17.4938
R16187 dvdd.n557 dvdd.n556 17.4938
R16188 dvdd.n561 dvdd.n560 17.4938
R16189 dvdd.n349 dvdd.n296 16.9359
R16190 dvdd.n360 dvdd.n359 16.9359
R16191 dvdd.n245 dvdd.n235 16.132
R16192 dvdd.n250 dvdd.n247 16.132
R16193 dvdd.n254 dvdd.n232 16.132
R16194 dvdd.n265 dvdd.n264 16.132
R16195 dvdd.n270 dvdd.n268 16.132
R16196 dvdd.n274 dvdd.n224 16.132
R16197 dvdd.n275 dvdd.n274 16.132
R16198 dvdd.n241 dvdd.n238 15.9567
R16199 dvdd.n105 dvdd.n95 15.914
R16200 dvdd.n110 dvdd.n107 15.914
R16201 dvdd.n114 dvdd.n92 15.914
R16202 dvdd.n125 dvdd.n124 15.914
R16203 dvdd.n130 dvdd.n128 15.914
R16204 dvdd.n134 dvdd.n84 15.914
R16205 dvdd.n135 dvdd.n134 15.914
R16206 dvdd.n162 dvdd.n152 15.914
R16207 dvdd.n167 dvdd.n164 15.914
R16208 dvdd.n171 dvdd.n149 15.914
R16209 dvdd.n182 dvdd.n181 15.914
R16210 dvdd.n187 dvdd.n185 15.914
R16211 dvdd.n191 dvdd.n141 15.914
R16212 dvdd.n192 dvdd.n191 15.914
R16213 dvdd.n347 dvdd.n299 15.7543
R16214 dvdd.n353 dvdd.n295 15.7543
R16215 dvdd.n101 dvdd.n98 15.741
R16216 dvdd.n158 dvdd.n155 15.741
R16217 dvdd.n263 dvdd.n262 15.606
R16218 dvdd.n335 dvdd.n304 15.5574
R16219 dvdd.n432 dvdd 15.5495
R16220 dvdd.n6 dvdd 15.5495
R16221 dvdd.n123 dvdd.n122 15.3951
R16222 dvdd.n180 dvdd.n179 15.3951
R16223 dvdd.n316 dvdd.n315 15.1636
R16224 dvdd.n340 dvdd.n300 15.1636
R16225 dvdd.n276 dvdd.n275 15.08
R16226 dvdd.n259 dvdd.n258 14.9046
R16227 dvdd.n119 dvdd.n118 14.8762
R16228 dvdd.n136 dvdd.n135 14.8762
R16229 dvdd.n176 dvdd.n175 14.8762
R16230 dvdd.n193 dvdd.n192 14.8762
R16231 dvdd.n258 dvdd.n257 14.2313
R16232 dvdd.n516 dvdd.n515 14.2313
R16233 dvdd.n513 dvdd.n509 14.2313
R16234 dvdd.n269 dvdd.n224 14.0279
R16235 dvdd.n262 dvdd.n229 13.8526
R16236 dvdd.n129 dvdd.n84 13.8383
R16237 dvdd.n186 dvdd.n141 13.8383
R16238 dvdd.n118 dvdd.n117 13.7042
R16239 dvdd.n175 dvdd.n174 13.7042
R16240 dvdd.n122 dvdd.n89 13.6654
R16241 dvdd.n179 dvdd.n146 13.6654
R16242 dvdd.n241 dvdd.n240 13.5019
R16243 dvdd.n265 dvdd.n225 13.5019
R16244 dvdd.n101 dvdd.n100 13.3194
R16245 dvdd.n125 dvdd.n85 13.3194
R16246 dvdd.n158 dvdd.n157 13.3194
R16247 dvdd.n182 dvdd.n142 13.3194
R16248 dvdd.n331 dvdd.n330 12.4067
R16249 dvdd.n321 dvdd.n320 12.0128
R16250 dvdd.n338 dvdd.n337 12.0128
R16251 dvdd.n337 dvdd.n336 11.2126
R16252 dvdd.n256 dvdd.n255 11.0471
R16253 dvdd.n116 dvdd.n115 10.8978
R16254 dvdd.n173 dvdd.n172 10.8978
R16255 dvdd.n246 dvdd.n245 10.6964
R16256 dvdd.n106 dvdd.n105 10.5519
R16257 dvdd.n163 dvdd.n162 10.5519
R16258 dvdd.n361 dvdd.n360 10.482
R16259 dvdd.n277 dvdd.n276 10.3526
R16260 dvdd.n137 dvdd.n136 10.3383
R16261 dvdd.n194 dvdd.n193 10.3383
R16262 dvdd.n434 dvdd.n433 10.0534
R16263 dvdd.n8 dvdd.n7 10.0534
R16264 dvdd.n471 dvdd.n362 9.76224
R16265 dvdd.n81 dvdd.n80 9.3005
R16266 dvdd.n242 dvdd.n241 9.3005
R16267 dvdd.n243 dvdd.n235 9.3005
R16268 dvdd.n245 dvdd.n244 9.3005
R16269 dvdd.n247 dvdd.n233 9.3005
R16270 dvdd.n251 dvdd.n250 9.3005
R16271 dvdd.n252 dvdd.n232 9.3005
R16272 dvdd.n254 dvdd.n253 9.3005
R16273 dvdd.n256 dvdd.n230 9.3005
R16274 dvdd.n260 dvdd.n259 9.3005
R16275 dvdd.n262 dvdd.n261 9.3005
R16276 dvdd.n264 dvdd.n226 9.3005
R16277 dvdd.n266 dvdd.n265 9.3005
R16278 dvdd.n268 dvdd.n267 9.3005
R16279 dvdd.n271 dvdd.n270 9.3005
R16280 dvdd.n272 dvdd.n224 9.3005
R16281 dvdd.n274 dvdd.n273 9.3005
R16282 dvdd.n275 dvdd.n222 9.3005
R16283 dvdd.n135 dvdd.n82 9.3005
R16284 dvdd.n134 dvdd.n133 9.3005
R16285 dvdd.n132 dvdd.n84 9.3005
R16286 dvdd.n131 dvdd.n130 9.3005
R16287 dvdd.n128 dvdd.n127 9.3005
R16288 dvdd.n126 dvdd.n125 9.3005
R16289 dvdd.n124 dvdd.n86 9.3005
R16290 dvdd.n122 dvdd.n121 9.3005
R16291 dvdd.n120 dvdd.n119 9.3005
R16292 dvdd.n116 dvdd.n90 9.3005
R16293 dvdd.n114 dvdd.n113 9.3005
R16294 dvdd.n112 dvdd.n92 9.3005
R16295 dvdd.n111 dvdd.n110 9.3005
R16296 dvdd.n107 dvdd.n93 9.3005
R16297 dvdd.n105 dvdd.n104 9.3005
R16298 dvdd.n103 dvdd.n95 9.3005
R16299 dvdd.n102 dvdd.n101 9.3005
R16300 dvdd.n192 dvdd.n139 9.3005
R16301 dvdd.n191 dvdd.n190 9.3005
R16302 dvdd.n189 dvdd.n141 9.3005
R16303 dvdd.n188 dvdd.n187 9.3005
R16304 dvdd.n185 dvdd.n184 9.3005
R16305 dvdd.n183 dvdd.n182 9.3005
R16306 dvdd.n181 dvdd.n143 9.3005
R16307 dvdd.n179 dvdd.n178 9.3005
R16308 dvdd.n177 dvdd.n176 9.3005
R16309 dvdd.n173 dvdd.n147 9.3005
R16310 dvdd.n171 dvdd.n170 9.3005
R16311 dvdd.n169 dvdd.n149 9.3005
R16312 dvdd.n168 dvdd.n167 9.3005
R16313 dvdd.n164 dvdd.n150 9.3005
R16314 dvdd.n162 dvdd.n161 9.3005
R16315 dvdd.n160 dvdd.n152 9.3005
R16316 dvdd.n159 dvdd.n158 9.3005
R16317 dvdd.n352 dvdd.n351 9.3005
R16318 dvdd.n359 dvdd.n293 9.3005
R16319 dvdd.n358 dvdd.n357 9.3005
R16320 dvdd.n356 dvdd.n295 9.3005
R16321 dvdd.n355 dvdd.n354 9.3005
R16322 dvdd.n350 dvdd.n349 9.3005
R16323 dvdd.n348 dvdd.n297 9.3005
R16324 dvdd.n347 dvdd.n346 9.3005
R16325 dvdd.n345 dvdd.n344 9.3005
R16326 dvdd.n343 dvdd.n342 9.3005
R16327 dvdd.n341 dvdd.n340 9.3005
R16328 dvdd.n339 dvdd.n301 9.3005
R16329 dvdd.n335 dvdd.n334 9.3005
R16330 dvdd.n333 dvdd.n332 9.3005
R16331 dvdd.n331 dvdd.n305 9.3005
R16332 dvdd.n329 dvdd.n328 9.3005
R16333 dvdd.n327 dvdd.n307 9.3005
R16334 dvdd.n326 dvdd.n325 9.3005
R16335 dvdd.n322 dvdd.n308 9.3005
R16336 dvdd.n320 dvdd.n319 9.3005
R16337 dvdd.n318 dvdd.n310 9.3005
R16338 dvdd.n317 dvdd.n316 9.3005
R16339 dvdd.n438 dvdd.n437 9.3005
R16340 dvdd.n442 dvdd.n441 9.3005
R16341 dvdd.n446 dvdd.n445 9.3005
R16342 dvdd.n450 dvdd.n449 9.3005
R16343 dvdd.n454 dvdd.n453 9.3005
R16344 dvdd.n458 dvdd.n457 9.3005
R16345 dvdd.n462 dvdd.n461 9.3005
R16346 dvdd.n466 dvdd.n465 9.3005
R16347 dvdd.n470 dvdd.n469 9.3005
R16348 dvdd.n560 dvdd.n559 9.3005
R16349 dvdd.n556 dvdd.n555 9.3005
R16350 dvdd.n552 dvdd.n551 9.3005
R16351 dvdd.n548 dvdd.n547 9.3005
R16352 dvdd.n544 dvdd.n543 9.3005
R16353 dvdd.n540 dvdd.n539 9.3005
R16354 dvdd.n536 dvdd.n535 9.3005
R16355 dvdd.n532 dvdd.n531 9.3005
R16356 dvdd.n528 dvdd.n527 9.3005
R16357 dvdd.n517 dvdd.n508 9.3005
R16358 dvdd.n324 dvdd.n307 9.25588
R16359 dvdd.n325 dvdd.n324 8.86204
R16360 dvdd.n249 dvdd.n232 8.2416
R16361 dvdd.n290 dvdd.n289 8.2025
R16362 dvdd.n487 dvdd.n475 8.19123
R16363 dvdd.n109 dvdd.n92 8.13023
R16364 dvdd.n166 dvdd.n149 8.13023
R16365 dvdd.n250 dvdd.n249 7.89091
R16366 dvdd.n110 dvdd.n109 7.78428
R16367 dvdd.n167 dvdd.n166 7.78428
R16368 dvdd.n138 dvdd 7.76009
R16369 dvdd.n520 dvdd.n487 6.79735
R16370 dvdd.n433 dvdd.n432 6.58874
R16371 dvdd.n7 dvdd.n6 6.58874
R16372 dvdd.n313 dvdd.n311 6.14225
R16373 dvdd.n322 dvdd.n321 6.10512
R16374 dvdd.n514 dvdd.t176 6.06249
R16375 dvdd.n218 dvdd.n199 5.96824
R16376 dvdd.t52 dvdd.n199 5.96824
R16377 dvdd.n214 dvdd.n213 5.96824
R16378 dvdd.t52 dvdd.n214 5.96824
R16379 dvdd.n521 dvdd.n474 5.9447
R16380 dvdd.n507 dvdd.n474 5.94023
R16381 dvdd.n238 dvdd.n236 5.87299
R16382 dvdd.n98 dvdd.n96 5.84114
R16383 dvdd.n155 dvdd.n153 5.84114
R16384 dvdd.n330 dvdd.n329 5.71127
R16385 dvdd.n337 dvdd.n335 5.51435
R16386 dvdd.n247 dvdd.n246 5.43612
R16387 dvdd.n107 dvdd.n106 5.36266
R16388 dvdd.n164 dvdd.n163 5.36266
R16389 dvdd.n362 dvdd 5.14764
R16390 dvdd.n195 dvdd 5.14243
R16391 dvdd.n138 dvdd 5.13722
R16392 dvdd.n255 dvdd.n254 5.08543
R16393 dvdd.n115 dvdd.n114 5.01672
R16394 dvdd.n172 dvdd.n171 5.01672
R16395 dvdd.n292 dvdd.n291 4.5005
R16396 dvdd.n79 dvdd.n78 4.32258
R16397 dvdd.n468 dvdd.n369 4.32258
R16398 dvdd.n464 dvdd.n376 4.32258
R16399 dvdd.n460 dvdd.n383 4.32258
R16400 dvdd.n456 dvdd.n390 4.32258
R16401 dvdd.n452 dvdd.n397 4.32258
R16402 dvdd.n448 dvdd.n404 4.32258
R16403 dvdd.n444 dvdd.n411 4.32258
R16404 dvdd.n440 dvdd.n418 4.32258
R16405 dvdd.n436 dvdd.n425 4.32258
R16406 dvdd.n529 dvdd.n70 4.32258
R16407 dvdd.n533 dvdd.n63 4.32258
R16408 dvdd.n537 dvdd.n56 4.32258
R16409 dvdd.n541 dvdd.n49 4.32258
R16410 dvdd.n545 dvdd.n42 4.32258
R16411 dvdd.n549 dvdd.n35 4.32258
R16412 dvdd.n553 dvdd.n28 4.32258
R16413 dvdd.n557 dvdd.n21 4.32258
R16414 dvdd.n561 dvdd.n14 4.32258
R16415 dvdd.n520 dvdd.n519 4.29291
R16416 dvdd.n508 dvdd.n507 4.26836
R16417 dvdd.n525 dvdd 4.0955
R16418 dvdd.n471 dvdd 3.73954
R16419 dvdd dvdd.n526 3.73954
R16420 dvdd.n512 dvdd.n511 3.36414
R16421 dvdd.n514 dvdd.n512 3.36414
R16422 dvdd.n518 dvdd.n510 3.36414
R16423 dvdd.n514 dvdd.n510 3.36414
R16424 dvdd.n220 dvdd.n219 3.36211
R16425 dvdd.n432 dvdd.n431 3.34378
R16426 dvdd.n6 dvdd.n5 3.34378
R16427 dvdd.n283 dvdd.n279 3.13609
R16428 dvdd.n284 dvdd.n283 3.13609
R16429 dvdd.n288 dvdd.n287 3.13609
R16430 dvdd.n287 dvdd.n286 3.13609
R16431 dvdd.n315 dvdd.n310 2.95435
R16432 dvdd.n343 dvdd.n300 2.95435
R16433 dvdd.n435 dvdd 2.9391
R16434 dvdd.n439 dvdd 2.9391
R16435 dvdd.n443 dvdd 2.9391
R16436 dvdd.n447 dvdd 2.9391
R16437 dvdd.n451 dvdd 2.9391
R16438 dvdd.n455 dvdd 2.9391
R16439 dvdd.n459 dvdd 2.9391
R16440 dvdd.n463 dvdd 2.9391
R16441 dvdd.n467 dvdd 2.9391
R16442 dvdd dvdd.n558 2.9391
R16443 dvdd dvdd.n554 2.9391
R16444 dvdd dvdd.n550 2.9391
R16445 dvdd dvdd.n546 2.9391
R16446 dvdd dvdd.n542 2.9391
R16447 dvdd dvdd.n538 2.9391
R16448 dvdd dvdd.n534 2.9391
R16449 dvdd dvdd.n530 2.9391
R16450 dvdd dvdd.n562 2.9369
R16451 dvdd.n203 dvdd.n197 2.90005
R16452 dvdd.n480 dvdd.n476 2.80353
R16453 dvdd.n481 dvdd.n480 2.80353
R16454 dvdd.n485 dvdd.n484 2.80353
R16455 dvdd.n484 dvdd.n483 2.80353
R16456 dvdd.n240 dvdd.n235 2.63064
R16457 dvdd.n268 dvdd.n225 2.63064
R16458 dvdd.n100 dvdd.n95 2.59509
R16459 dvdd.n128 dvdd.n85 2.59509
R16460 dvdd.n157 dvdd.n152 2.59509
R16461 dvdd.n185 dvdd.n142 2.59509
R16462 dvdd.n332 dvdd.n304 2.5605
R16463 dvdd.n221 dvdd.n220 2.52884
R16464 dvdd.n344 dvdd.n299 2.36358
R16465 dvdd.n354 dvdd.n353 2.36358
R16466 dvdd.n259 dvdd.n229 2.27995
R16467 dvdd.n119 dvdd.n89 2.24915
R16468 dvdd.n176 dvdd.n146 2.24915
R16469 dvdd.n270 dvdd.n269 2.10461
R16470 dvdd.n281 dvdd.n278 2.10277
R16471 dvdd.n285 dvdd.n281 2.10277
R16472 dvdd.n289 dvdd.n280 2.10277
R16473 dvdd.n282 dvdd.n280 2.10277
R16474 dvdd.n130 dvdd.n129 2.07618
R16475 dvdd.n187 dvdd.n186 2.07618
R16476 dvdd.n526 dvdd.n471 1.69386
R16477 dvdd.n292 dvdd.n221 1.26417
R16478 dvdd.n258 dvdd.n256 1.2279
R16479 dvdd.n352 dvdd.n296 1.18204
R16480 dvdd.n102 dvdd.n96 1.06234
R16481 dvdd.n159 dvdd.n153 1.06234
R16482 dvdd.n242 dvdd.n236 1.05227
R16483 dvdd.n118 dvdd.n116 1.03834
R16484 dvdd.n175 dvdd.n173 1.03834
R16485 dvdd.n317 dvdd.n311 0.968765
R16486 dvdd.n219 dvdd.n197 0.955857
R16487 dvdd.n526 dvdd.n525 0.951672
R16488 dvdd.n221 dvdd.n195 0.836438
R16489 dvdd.n195 dvdd.n138 0.808117
R16490 dvdd.n494 dvdd.n493 0.787085
R16491 dvdd.n204 dvdd.n203 0.705857
R16492 dvdd.n205 dvdd.n204 0.705857
R16493 dvdd.n211 dvdd.n210 0.705857
R16494 dvdd.n210 dvdd.n209 0.705857
R16495 dvdd.n209 dvdd.n196 0.705857
R16496 dvdd.n362 dvdd.n292 0.691906
R16497 dvdd.n291 dvdd 0.645031
R16498 dvdd.n291 dvdd.n290 0.633614
R16499 dvdd.n339 dvdd.n338 0.591269
R16500 dvdd.n212 dvdd.n205 0.529518
R16501 dvdd.n264 dvdd.n263 0.526527
R16502 dvdd.n124 dvdd.n123 0.519419
R16503 dvdd.n181 dvdd.n180 0.519419
R16504 dvdd.n290 dvdd.n278 0.517903
R16505 dvdd.n493 dvdd.n492 0.514219
R16506 dvdd.n506 dvdd.n505 0.492878
R16507 dvdd.n491 dvdd.n473 0.482207
R16508 dvdd.n502 dvdd.n494 0.482207
R16509 dvdd.n503 dvdd.n502 0.482207
R16510 dvdd.n504 dvdd.n503 0.482207
R16511 dvdd.n478 dvdd.n475 0.448442
R16512 dvdd.n479 dvdd.n478 0.448442
R16513 dvdd.n486 dvdd.n477 0.448442
R16514 dvdd.n482 dvdd.n477 0.448442
R16515 dvdd.n522 dvdd.n473 0.447146
R16516 dvdd.n507 dvdd.n506 0.419707
R16517 dvdd.n505 dvdd.n504 0.386171
R16518 dvdd.n522 dvdd.n521 0.372451
R16519 dvdd.n492 dvdd.n491 0.361781
R16520 dvdd.n220 dvdd.n196 0.346482
R16521 dvdd.n213 dvdd.n212 0.3105
R16522 dvdd.n219 dvdd.n218 0.3105
R16523 dvdd.n508 dvdd.n494 0.307565
R16524 dvdd.n519 dvdd.n508 0.272821
R16525 dvdd.n521 dvdd.n520 0.252732
R16526 dvdd.n506 dvdd.n497 0.206229
R16527 dvdd.n511 dvdd.n474 0.179346
R16528 dvdd.n519 dvdd.n518 0.179346
R16529 dvdd.n212 dvdd.n211 0.176839
R16530 dvdd.n504 dvdd.n499 0.152674
R16531 dvdd.n81 dvdd 0.121114
R16532 dvdd.n434 dvdd 0.121114
R16533 dvdd.n438 dvdd 0.121114
R16534 dvdd.n442 dvdd 0.121114
R16535 dvdd.n446 dvdd 0.121114
R16536 dvdd.n450 dvdd 0.121114
R16537 dvdd.n454 dvdd 0.121114
R16538 dvdd.n458 dvdd 0.121114
R16539 dvdd.n462 dvdd 0.121114
R16540 dvdd.n466 dvdd 0.121114
R16541 dvdd.n470 dvdd 0.121114
R16542 dvdd.n8 dvdd 0.121114
R16543 dvdd.n559 dvdd 0.121114
R16544 dvdd.n555 dvdd 0.121114
R16545 dvdd.n551 dvdd 0.121114
R16546 dvdd.n547 dvdd 0.121114
R16547 dvdd.n543 dvdd 0.121114
R16548 dvdd.n539 dvdd 0.121114
R16549 dvdd.n535 dvdd 0.121114
R16550 dvdd.n531 dvdd 0.121114
R16551 dvdd.n527 dvdd 0.121114
R16552 dvdd.n243 dvdd.n242 0.120292
R16553 dvdd.n244 dvdd.n243 0.120292
R16554 dvdd.n244 dvdd.n233 0.120292
R16555 dvdd.n251 dvdd.n233 0.120292
R16556 dvdd.n252 dvdd.n251 0.120292
R16557 dvdd.n253 dvdd.n252 0.120292
R16558 dvdd.n253 dvdd.n230 0.120292
R16559 dvdd.n260 dvdd.n230 0.120292
R16560 dvdd.n261 dvdd.n260 0.120292
R16561 dvdd.n261 dvdd.n226 0.120292
R16562 dvdd.n266 dvdd.n226 0.120292
R16563 dvdd.n267 dvdd.n266 0.120292
R16564 dvdd.n272 dvdd.n271 0.120292
R16565 dvdd.n273 dvdd.n272 0.120292
R16566 dvdd.n273 dvdd.n222 0.120292
R16567 dvdd.n277 dvdd.n222 0.120292
R16568 dvdd.n103 dvdd.n102 0.120292
R16569 dvdd.n104 dvdd.n103 0.120292
R16570 dvdd.n104 dvdd.n93 0.120292
R16571 dvdd.n111 dvdd.n93 0.120292
R16572 dvdd.n112 dvdd.n111 0.120292
R16573 dvdd.n113 dvdd.n112 0.120292
R16574 dvdd.n113 dvdd.n90 0.120292
R16575 dvdd.n120 dvdd.n90 0.120292
R16576 dvdd.n121 dvdd.n120 0.120292
R16577 dvdd.n121 dvdd.n86 0.120292
R16578 dvdd.n126 dvdd.n86 0.120292
R16579 dvdd.n127 dvdd.n126 0.120292
R16580 dvdd.n132 dvdd.n131 0.120292
R16581 dvdd.n133 dvdd.n132 0.120292
R16582 dvdd.n133 dvdd.n82 0.120292
R16583 dvdd.n137 dvdd.n82 0.120292
R16584 dvdd.n160 dvdd.n159 0.120292
R16585 dvdd.n161 dvdd.n160 0.120292
R16586 dvdd.n161 dvdd.n150 0.120292
R16587 dvdd.n168 dvdd.n150 0.120292
R16588 dvdd.n169 dvdd.n168 0.120292
R16589 dvdd.n170 dvdd.n169 0.120292
R16590 dvdd.n170 dvdd.n147 0.120292
R16591 dvdd.n177 dvdd.n147 0.120292
R16592 dvdd.n178 dvdd.n177 0.120292
R16593 dvdd.n178 dvdd.n143 0.120292
R16594 dvdd.n183 dvdd.n143 0.120292
R16595 dvdd.n184 dvdd.n183 0.120292
R16596 dvdd.n189 dvdd.n188 0.120292
R16597 dvdd.n190 dvdd.n189 0.120292
R16598 dvdd.n190 dvdd.n139 0.120292
R16599 dvdd.n194 dvdd.n139 0.120292
R16600 dvdd.n318 dvdd.n317 0.120292
R16601 dvdd.n319 dvdd.n318 0.120292
R16602 dvdd.n319 dvdd.n308 0.120292
R16603 dvdd.n326 dvdd.n308 0.120292
R16604 dvdd.n327 dvdd.n326 0.120292
R16605 dvdd.n328 dvdd.n327 0.120292
R16606 dvdd.n328 dvdd.n305 0.120292
R16607 dvdd.n333 dvdd.n305 0.120292
R16608 dvdd.n334 dvdd.n333 0.120292
R16609 dvdd.n334 dvdd.n301 0.120292
R16610 dvdd.n341 dvdd.n301 0.120292
R16611 dvdd.n342 dvdd.n341 0.120292
R16612 dvdd.n346 dvdd.n345 0.120292
R16613 dvdd.n346 dvdd.n297 0.120292
R16614 dvdd.n350 dvdd.n297 0.120292
R16615 dvdd.n351 dvdd.n350 0.120292
R16616 dvdd.n356 dvdd.n355 0.120292
R16617 dvdd.n357 dvdd.n356 0.120292
R16618 dvdd.n357 dvdd.n293 0.120292
R16619 dvdd.n361 dvdd.n293 0.120292
R16620 dvdd.n524 dvdd.n522 0.0789314
R16621 dvdd.n271 dvdd 0.0603958
R16622 dvdd.n131 dvdd 0.0603958
R16623 dvdd.n188 dvdd 0.0603958
R16624 dvdd.n345 dvdd 0.0603958
R16625 dvdd.n355 dvdd 0.0603958
R16626 dvdd dvdd.n81 0.0377807
R16627 dvdd dvdd.n434 0.0377807
R16628 dvdd.n435 dvdd 0.0377807
R16629 dvdd dvdd.n438 0.0377807
R16630 dvdd.n439 dvdd 0.0377807
R16631 dvdd dvdd.n442 0.0377807
R16632 dvdd.n443 dvdd 0.0377807
R16633 dvdd dvdd.n446 0.0377807
R16634 dvdd.n447 dvdd 0.0377807
R16635 dvdd dvdd.n450 0.0377807
R16636 dvdd.n451 dvdd 0.0377807
R16637 dvdd dvdd.n454 0.0377807
R16638 dvdd.n455 dvdd 0.0377807
R16639 dvdd dvdd.n458 0.0377807
R16640 dvdd.n459 dvdd 0.0377807
R16641 dvdd dvdd.n462 0.0377807
R16642 dvdd.n463 dvdd 0.0377807
R16643 dvdd dvdd.n466 0.0377807
R16644 dvdd.n467 dvdd 0.0377807
R16645 dvdd dvdd.n470 0.0377807
R16646 dvdd dvdd.n8 0.0377807
R16647 dvdd.n562 dvdd 0.0377807
R16648 dvdd.n559 dvdd 0.0377807
R16649 dvdd.n558 dvdd 0.0377807
R16650 dvdd.n555 dvdd 0.0377807
R16651 dvdd.n554 dvdd 0.0377807
R16652 dvdd.n551 dvdd 0.0377807
R16653 dvdd.n550 dvdd 0.0377807
R16654 dvdd.n547 dvdd 0.0377807
R16655 dvdd.n546 dvdd 0.0377807
R16656 dvdd.n543 dvdd 0.0377807
R16657 dvdd.n542 dvdd 0.0377807
R16658 dvdd.n539 dvdd 0.0377807
R16659 dvdd.n538 dvdd 0.0377807
R16660 dvdd.n535 dvdd 0.0377807
R16661 dvdd.n534 dvdd 0.0377807
R16662 dvdd.n531 dvdd 0.0377807
R16663 dvdd.n530 dvdd 0.0377807
R16664 dvdd.n527 dvdd 0.0377807
R16665 dvdd.n267 dvdd 0.0226354
R16666 dvdd dvdd.n277 0.0226354
R16667 dvdd.n127 dvdd 0.0226354
R16668 dvdd dvdd.n137 0.0226354
R16669 dvdd.n184 dvdd 0.0226354
R16670 dvdd dvdd.n194 0.0226354
R16671 dvdd.n342 dvdd 0.0226354
R16672 dvdd.n351 dvdd 0.0226354
R16673 dvdd dvdd.n361 0.0226354
R16674 osc_ck.n1 osc_ck.t5 236.361
R16675 osc_ck.n4 osc_ck.n2 214.567
R16676 osc_ck.n1 osc_ck.n0 207.792
R16677 osc_ck.n5 osc_ck.t3 88.3503
R16678 osc_ck.n4 osc_ck.n3 70.9231
R16679 osc_ck.n2 osc_ck.t7 29.5505
R16680 osc_ck.n2 osc_ck.t0 29.5505
R16681 osc_ck.n0 osc_ck.t4 28.5655
R16682 osc_ck.n0 osc_ck.t6 28.5655
R16683 osc_ck.n3 osc_ck.t1 18.0005
R16684 osc_ck.n3 osc_ck.t2 18.0005
R16685 osc_ck osc_ck.n5 9.94118
R16686 osc_ck.n5 osc_ck.n4 7.92796
R16687 osc_ck osc_ck.n1 3.48967
R16688 rc_osc_0.n.n4 rc_osc_0.n.t6 244.843
R16689 rc_osc_0.n.n2 rc_osc_0.n.t11 240.778
R16690 rc_osc_0.n.n3 rc_osc_0.n.t13 240.349
R16691 rc_osc_0.n.n2 rc_osc_0.n.t9 240.349
R16692 rc_osc_0.n.n10 rc_osc_0.n.n0 211.296
R16693 rc_osc_0.n.n11 rc_osc_0.n.n10 204.284
R16694 rc_osc_0.n.n7 rc_osc_0.n.t10 123.462
R16695 rc_osc_0.n.n5 rc_osc_0.n.t7 120.871
R16696 rc_osc_0.n.n6 rc_osc_0.n.t8 120.773
R16697 rc_osc_0.n.n5 rc_osc_0.n.t12 120.174
R16698 rc_osc_0.n.n9 rc_osc_0.n.n1 72.3553
R16699 rc_osc_0.n.n0 rc_osc_0.n.t1 28.5655
R16700 rc_osc_0.n.n0 rc_osc_0.n.t2 28.5655
R16701 rc_osc_0.n.n11 rc_osc_0.n.t3 28.5655
R16702 rc_osc_0.n.t5 rc_osc_0.n.n11 28.5655
R16703 rc_osc_0.n.n1 rc_osc_0.n.t4 17.4005
R16704 rc_osc_0.n.n1 rc_osc_0.n.t0 17.4005
R16705 rc_osc_0.n.n4 rc_osc_0.n.n3 9.0153
R16706 rc_osc_0.n.n7 rc_osc_0.n.n6 5.23012
R16707 rc_osc_0.n.n8 rc_osc_0.n.n7 3.78258
R16708 rc_osc_0.n.n9 rc_osc_0.n.n8 3.4105
R16709 rc_osc_0.n.n10 rc_osc_0.n.n9 1.35184
R16710 rc_osc_0.n.n3 rc_osc_0.n.n2 0.408448
R16711 rc_osc_0.n.n8 rc_osc_0.n.n4 0.147461
R16712 rc_osc_0.n.n6 rc_osc_0.n.n5 0.049413
R16713 pwup_filt.n2 pwup_filt.n0 243.458
R16714 pwup_filt.n2 pwup_filt.n1 205.059
R16715 pwup_filt.n4 pwup_filt.n3 205.059
R16716 pwup_filt.n6 pwup_filt.n5 205.059
R16717 pwup_filt.n8 pwup_filt.n7 205.059
R16718 pwup_filt.n10 pwup_filt.n9 205.059
R16719 pwup_filt.n12 pwup_filt.n11 205.059
R16720 pwup_filt.n14 pwup_filt.n13 205.059
R16721 pwup_filt.n18 pwup_filt.n16 133.534
R16722 pwup_filt.n18 pwup_filt.n17 99.1759
R16723 pwup_filt.n20 pwup_filt.n19 99.1759
R16724 pwup_filt.n22 pwup_filt.n21 99.1759
R16725 pwup_filt.n24 pwup_filt.n23 99.1759
R16726 pwup_filt.n26 pwup_filt.n25 99.1759
R16727 pwup_filt.n28 pwup_filt.n27 99.1759
R16728 pwup_filt pwup_filt.n29 97.4305
R16729 pwup_filt.n4 pwup_filt.n2 38.4005
R16730 pwup_filt.n6 pwup_filt.n4 38.4005
R16731 pwup_filt.n8 pwup_filt.n6 38.4005
R16732 pwup_filt.n10 pwup_filt.n8 38.4005
R16733 pwup_filt.n12 pwup_filt.n10 38.4005
R16734 pwup_filt.n14 pwup_filt.n12 38.4005
R16735 pwup_filt.n20 pwup_filt.n18 34.3584
R16736 pwup_filt.n22 pwup_filt.n20 34.3584
R16737 pwup_filt.n24 pwup_filt.n22 34.3584
R16738 pwup_filt.n26 pwup_filt.n24 34.3584
R16739 pwup_filt.n28 pwup_filt.n26 34.3584
R16740 pwup_filt.n30 pwup_filt.n28 34.3584
R16741 pwup_filt.n13 pwup_filt.t19 26.5955
R16742 pwup_filt.n13 pwup_filt.t25 26.5955
R16743 pwup_filt.n0 pwup_filt.t17 26.5955
R16744 pwup_filt.n0 pwup_filt.t24 26.5955
R16745 pwup_filt.n1 pwup_filt.t31 26.5955
R16746 pwup_filt.n1 pwup_filt.t27 26.5955
R16747 pwup_filt.n3 pwup_filt.t30 26.5955
R16748 pwup_filt.n3 pwup_filt.t22 26.5955
R16749 pwup_filt.n5 pwup_filt.t18 26.5955
R16750 pwup_filt.n5 pwup_filt.t21 26.5955
R16751 pwup_filt.n7 pwup_filt.t29 26.5955
R16752 pwup_filt.n7 pwup_filt.t23 26.5955
R16753 pwup_filt.n9 pwup_filt.t16 26.5955
R16754 pwup_filt.n9 pwup_filt.t28 26.5955
R16755 pwup_filt.n11 pwup_filt.t20 26.5955
R16756 pwup_filt.n11 pwup_filt.t26 26.5955
R16757 pwup_filt.n29 pwup_filt.t14 24.9236
R16758 pwup_filt.n29 pwup_filt.t4 24.9236
R16759 pwup_filt.n16 pwup_filt.t12 24.9236
R16760 pwup_filt.n16 pwup_filt.t3 24.9236
R16761 pwup_filt.n17 pwup_filt.t10 24.9236
R16762 pwup_filt.n17 pwup_filt.t6 24.9236
R16763 pwup_filt.n19 pwup_filt.t9 24.9236
R16764 pwup_filt.n19 pwup_filt.t1 24.9236
R16765 pwup_filt.n21 pwup_filt.t13 24.9236
R16766 pwup_filt.n21 pwup_filt.t0 24.9236
R16767 pwup_filt.n23 pwup_filt.t8 24.9236
R16768 pwup_filt.n23 pwup_filt.t2 24.9236
R16769 pwup_filt.n25 pwup_filt.t11 24.9236
R16770 pwup_filt.n25 pwup_filt.t7 24.9236
R16771 pwup_filt.n27 pwup_filt.t15 24.9236
R16772 pwup_filt.n27 pwup_filt.t5 24.9236
R16773 pwup_filt.n15 pwup_filt.n14 12.6066
R16774 pwup_filt pwup_filt.n30 11.4429
R16775 pwup_filt pwup_filt.n15 5.81868
R16776 pwup_filt.n15 pwup_filt 4.52868
R16777 pwup_filt.n30 pwup_filt 1.74595
R16778 rstring_mux_0.vtop.n4 rstring_mux_0.vtop.t0 87.3599
R16779 rstring_mux_0.vtop.n2 rstring_mux_0.vtop.n0 48.5415
R16780 rstring_mux_0.vtop.n13 rstring_mux_0.vtop.n12 48.4284
R16781 rstring_mux_0.vtop.n11 rstring_mux_0.vtop.n10 48.4284
R16782 rstring_mux_0.vtop.n9 rstring_mux_0.vtop.n8 48.4284
R16783 rstring_mux_0.vtop.n7 rstring_mux_0.vtop.n6 48.4284
R16784 rstring_mux_0.vtop.n2 rstring_mux_0.vtop.n1 48.4284
R16785 rstring_mux_0.vtop.n15 rstring_mux_0.vtop.n14 45.0184
R16786 rstring_mux_0.vtop.n4 rstring_mux_0.vtop.n3 45.0184
R16787 rstring_mux_0.vtop rstring_mux_0.vtop.t17 19.1879
R16788 rstring_mux_0.vtop.n14 rstring_mux_0.vtop.t4 5.5395
R16789 rstring_mux_0.vtop.n14 rstring_mux_0.vtop.t11 5.5395
R16790 rstring_mux_0.vtop.n12 rstring_mux_0.vtop.t5 5.5395
R16791 rstring_mux_0.vtop.n12 rstring_mux_0.vtop.t13 5.5395
R16792 rstring_mux_0.vtop.n10 rstring_mux_0.vtop.t7 5.5395
R16793 rstring_mux_0.vtop.n10 rstring_mux_0.vtop.t15 5.5395
R16794 rstring_mux_0.vtop.n8 rstring_mux_0.vtop.t2 5.5395
R16795 rstring_mux_0.vtop.n8 rstring_mux_0.vtop.t9 5.5395
R16796 rstring_mux_0.vtop.n6 rstring_mux_0.vtop.t3 5.5395
R16797 rstring_mux_0.vtop.n6 rstring_mux_0.vtop.t10 5.5395
R16798 rstring_mux_0.vtop.n3 rstring_mux_0.vtop.t14 5.5395
R16799 rstring_mux_0.vtop.n3 rstring_mux_0.vtop.t12 5.5395
R16800 rstring_mux_0.vtop.n1 rstring_mux_0.vtop.t16 5.5395
R16801 rstring_mux_0.vtop.n1 rstring_mux_0.vtop.t6 5.5395
R16802 rstring_mux_0.vtop.n0 rstring_mux_0.vtop.t1 5.5395
R16803 rstring_mux_0.vtop.n0 rstring_mux_0.vtop.t8 5.5395
R16804 rstring_mux_0.vtop.n15 rstring_mux_0.vtop.n13 3.5118
R16805 rstring_mux_0.vtop.n5 rstring_mux_0.vtop.n4 3.4105
R16806 rstring_mux_0.vtop rstring_mux_0.vtop.n15 0.829892
R16807 rstring_mux_0.vtop.n5 rstring_mux_0.vtop.n2 0.113554
R16808 rstring_mux_0.vtop.n7 rstring_mux_0.vtop.n5 0.113554
R16809 rstring_mux_0.vtop.n9 rstring_mux_0.vtop.n7 0.113554
R16810 rstring_mux_0.vtop.n11 rstring_mux_0.vtop.n9 0.113554
R16811 rstring_mux_0.vtop.n13 rstring_mux_0.vtop.n11 0.113554
R16812 otrip_decoded[0].n0 otrip_decoded[0].t1 186.374
R16813 otrip_decoded[0].n0 otrip_decoded[0].t0 170.308
R16814 otrip_decoded[0] otrip_decoded[0].n1 154.56
R16815 otrip_decoded[0].n2 otrip_decoded[0].n1 153.462
R16816 otrip_decoded[0].n1 otrip_decoded[0].n0 101.513
R16817 otrip_decoded[0].n3 otrip_decoded[0] 11.8005
R16818 otrip_decoded[0].n3 otrip_decoded[0].n2 4.96991
R16819 otrip_decoded[0].n2 otrip_decoded[0] 3.46403
R16820 otrip_decoded[0] otrip_decoded[0].n3 2.71109
R16821 vbg_1v2.n52 vbg_1v2.t32 384.709
R16822 vbg_1v2.n51 vbg_1v2.t32 384.709
R16823 vbg_1v2.n62 vbg_1v2.t13 384.226
R16824 vbg_1v2.t13 vbg_1v2.n47 384.226
R16825 vbg_1v2.n61 vbg_1v2.t41 384.226
R16826 vbg_1v2.t41 vbg_1v2.n60 384.226
R16827 vbg_1v2.t1 vbg_1v2.n48 384.226
R16828 vbg_1v2.n59 vbg_1v2.t1 384.226
R16829 vbg_1v2.t4 vbg_1v2.n57 384.226
R16830 vbg_1v2.n58 vbg_1v2.t4 384.226
R16831 vbg_1v2.n56 vbg_1v2.t7 384.226
R16832 vbg_1v2.t7 vbg_1v2.n49 384.226
R16833 vbg_1v2.n55 vbg_1v2.t16 384.226
R16834 vbg_1v2.t16 vbg_1v2.n54 384.226
R16835 vbg_1v2.t22 vbg_1v2.n50 384.226
R16836 vbg_1v2.n53 vbg_1v2.t22 384.226
R16837 vbg_1v2.t29 vbg_1v2.n51 384.226
R16838 vbg_1v2.n52 vbg_1v2.t29 384.226
R16839 vbg_1v2.t23 vbg_1v2.n63 384.226
R16840 vbg_1v2.n64 vbg_1v2.t23 384.226
R16841 vbg_1v2.n46 vbg_1v2.n45 48.1045
R16842 vbg_1v2 vbg_1v2.n14 22.5215
R16843 vbg_1v2.n44 vbg_1v2.t11 14.8978
R16844 vbg_1v2.n43 vbg_1v2.t11 14.8978
R16845 vbg_1v2.n40 vbg_1v2.t14 14.8978
R16846 vbg_1v2.n39 vbg_1v2.t14 14.8978
R16847 vbg_1v2.n36 vbg_1v2.t25 14.8978
R16848 vbg_1v2.n35 vbg_1v2.t25 14.8978
R16849 vbg_1v2.n32 vbg_1v2.t3 14.8978
R16850 vbg_1v2.n31 vbg_1v2.t3 14.8978
R16851 vbg_1v2.n28 vbg_1v2.t24 14.8978
R16852 vbg_1v2.n27 vbg_1v2.t24 14.8978
R16853 vbg_1v2.n24 vbg_1v2.t34 14.8978
R16854 vbg_1v2.n23 vbg_1v2.t34 14.8978
R16855 vbg_1v2.n20 vbg_1v2.t8 14.8978
R16856 vbg_1v2.n19 vbg_1v2.t8 14.8978
R16857 vbg_1v2.n16 vbg_1v2.t20 14.8978
R16858 vbg_1v2.t20 vbg_1v2.n15 14.8978
R16859 vbg_1v2.t28 vbg_1v2.n43 12.9902
R16860 vbg_1v2.n44 vbg_1v2.t28 12.9902
R16861 vbg_1v2.t30 vbg_1v2.n39 12.9902
R16862 vbg_1v2.n40 vbg_1v2.t30 12.9902
R16863 vbg_1v2.t40 vbg_1v2.n35 12.9902
R16864 vbg_1v2.n36 vbg_1v2.t40 12.9902
R16865 vbg_1v2.t19 vbg_1v2.n31 12.9902
R16866 vbg_1v2.n32 vbg_1v2.t19 12.9902
R16867 vbg_1v2.t39 vbg_1v2.n27 12.9902
R16868 vbg_1v2.n28 vbg_1v2.t39 12.9902
R16869 vbg_1v2.t6 vbg_1v2.n23 12.9902
R16870 vbg_1v2.n24 vbg_1v2.t6 12.9902
R16871 vbg_1v2.t27 vbg_1v2.n19 12.9902
R16872 vbg_1v2.n20 vbg_1v2.t27 12.9902
R16873 vbg_1v2.t33 vbg_1v2.n15 12.9902
R16874 vbg_1v2.n16 vbg_1v2.t33 12.9902
R16875 vbg_1v2.n7 vbg_1v2.t15 9.72783
R16876 vbg_1v2.n0 vbg_1v2.t0 9.65028
R16877 vbg_1v2.n14 vbg_1v2.n6 8.96563
R16878 vbg_1v2.n13 vbg_1v2.t31 8.73727
R16879 vbg_1v2.n12 vbg_1v2.t21 8.73727
R16880 vbg_1v2.n11 vbg_1v2.t9 8.73727
R16881 vbg_1v2.n10 vbg_1v2.t35 8.73727
R16882 vbg_1v2.n9 vbg_1v2.t10 8.73727
R16883 vbg_1v2.n8 vbg_1v2.t36 8.73727
R16884 vbg_1v2.n7 vbg_1v2.t26 8.73727
R16885 vbg_1v2.n6 vbg_1v2.t12 8.65985
R16886 vbg_1v2.n5 vbg_1v2.t2 8.65985
R16887 vbg_1v2.n4 vbg_1v2.t37 8.65985
R16888 vbg_1v2.n3 vbg_1v2.t17 8.65985
R16889 vbg_1v2.n2 vbg_1v2.t38 8.65985
R16890 vbg_1v2.n1 vbg_1v2.t18 8.65985
R16891 vbg_1v2.n0 vbg_1v2.t5 8.65985
R16892 vbg_1v2.n14 vbg_1v2.n13 5.98511
R16893 vbg_1v2.n17 vbg_1v2.n15 5.24569
R16894 vbg_1v2.n17 vbg_1v2.n16 4.5005
R16895 vbg_1v2.n19 vbg_1v2.n18 4.5005
R16896 vbg_1v2.n21 vbg_1v2.n20 4.5005
R16897 vbg_1v2.n23 vbg_1v2.n22 4.5005
R16898 vbg_1v2.n25 vbg_1v2.n24 4.5005
R16899 vbg_1v2.n27 vbg_1v2.n26 4.5005
R16900 vbg_1v2.n29 vbg_1v2.n28 4.5005
R16901 vbg_1v2.n31 vbg_1v2.n30 4.5005
R16902 vbg_1v2.n33 vbg_1v2.n32 4.5005
R16903 vbg_1v2.n35 vbg_1v2.n34 4.5005
R16904 vbg_1v2.n37 vbg_1v2.n36 4.5005
R16905 vbg_1v2.n39 vbg_1v2.n38 4.5005
R16906 vbg_1v2.n41 vbg_1v2.n40 4.5005
R16907 vbg_1v2.n43 vbg_1v2.n42 4.5005
R16908 vbg_1v2.n45 vbg_1v2.n44 4.5005
R16909 vbg_1v2.n63 vbg_1v2.n46 4.5005
R16910 vbg_1v2.n65 vbg_1v2.n64 4.5005
R16911 vbg_1v2.n65 vbg_1v2.n46 2.63992
R16912 vbg_1v2.n13 vbg_1v2.n12 0.99106
R16913 vbg_1v2.n12 vbg_1v2.n11 0.99106
R16914 vbg_1v2.n11 vbg_1v2.n10 0.99106
R16915 vbg_1v2.n10 vbg_1v2.n9 0.99106
R16916 vbg_1v2.n9 vbg_1v2.n8 0.99106
R16917 vbg_1v2.n8 vbg_1v2.n7 0.99106
R16918 vbg_1v2.n6 vbg_1v2.n5 0.99093
R16919 vbg_1v2.n5 vbg_1v2.n4 0.99093
R16920 vbg_1v2.n4 vbg_1v2.n3 0.99093
R16921 vbg_1v2.n3 vbg_1v2.n2 0.99093
R16922 vbg_1v2.n2 vbg_1v2.n1 0.99093
R16923 vbg_1v2.n1 vbg_1v2.n0 0.99093
R16924 vbg_1v2.n45 vbg_1v2.n42 0.745692
R16925 vbg_1v2.n41 vbg_1v2.n38 0.745692
R16926 vbg_1v2.n37 vbg_1v2.n34 0.745692
R16927 vbg_1v2.n33 vbg_1v2.n30 0.745692
R16928 vbg_1v2.n29 vbg_1v2.n26 0.745692
R16929 vbg_1v2.n25 vbg_1v2.n22 0.745692
R16930 vbg_1v2.n21 vbg_1v2.n18 0.745692
R16931 vbg_1v2.n53 vbg_1v2.n52 0.484196
R16932 vbg_1v2.n54 vbg_1v2.n53 0.484196
R16933 vbg_1v2.n54 vbg_1v2.n49 0.484196
R16934 vbg_1v2.n58 vbg_1v2.n49 0.484196
R16935 vbg_1v2.n59 vbg_1v2.n58 0.484196
R16936 vbg_1v2.n60 vbg_1v2.n59 0.484196
R16937 vbg_1v2.n60 vbg_1v2.n47 0.484196
R16938 vbg_1v2.n51 vbg_1v2.n50 0.484196
R16939 vbg_1v2.n55 vbg_1v2.n50 0.484196
R16940 vbg_1v2.n56 vbg_1v2.n55 0.484196
R16941 vbg_1v2.n57 vbg_1v2.n56 0.484196
R16942 vbg_1v2.n57 vbg_1v2.n48 0.484196
R16943 vbg_1v2.n61 vbg_1v2.n48 0.484196
R16944 vbg_1v2.n62 vbg_1v2.n61 0.484196
R16945 vbg_1v2.n64 vbg_1v2.n47 0.459739
R16946 vbg_1v2.n63 vbg_1v2.n62 0.459739
R16947 vbg_1v2.n42 vbg_1v2.n41 0.260115
R16948 vbg_1v2.n38 vbg_1v2.n37 0.260115
R16949 vbg_1v2.n34 vbg_1v2.n33 0.260115
R16950 vbg_1v2.n30 vbg_1v2.n29 0.260115
R16951 vbg_1v2.n26 vbg_1v2.n25 0.260115
R16952 vbg_1v2.n22 vbg_1v2.n21 0.260115
R16953 vbg_1v2.n18 vbg_1v2.n17 0.260115
R16954 vbg_1v2 vbg_1v2.n65 0.063
R16955 dcomp.n2 dcomp.n0 243.458
R16956 dcomp.n2 dcomp.n1 205.059
R16957 dcomp.n4 dcomp.n3 205.059
R16958 dcomp.n6 dcomp.n5 205.059
R16959 dcomp.n8 dcomp.n7 205.059
R16960 dcomp.n10 dcomp.n9 205.059
R16961 dcomp.n12 dcomp.n11 205.059
R16962 dcomp.n14 dcomp.n13 205.059
R16963 dcomp.n17 dcomp.n15 133.534
R16964 dcomp.n17 dcomp.n16 99.1759
R16965 dcomp.n19 dcomp.n18 99.1759
R16966 dcomp.n21 dcomp.n20 99.1759
R16967 dcomp.n23 dcomp.n22 99.1759
R16968 dcomp.n25 dcomp.n24 99.1759
R16969 dcomp.n27 dcomp.n26 99.1759
R16970 dcomp dcomp.n28 97.4305
R16971 dcomp.n4 dcomp.n2 38.4005
R16972 dcomp.n6 dcomp.n4 38.4005
R16973 dcomp.n8 dcomp.n6 38.4005
R16974 dcomp.n10 dcomp.n8 38.4005
R16975 dcomp.n12 dcomp.n10 38.4005
R16976 dcomp.n14 dcomp.n12 38.4005
R16977 dcomp.n19 dcomp.n17 34.3584
R16978 dcomp.n21 dcomp.n19 34.3584
R16979 dcomp.n23 dcomp.n21 34.3584
R16980 dcomp.n25 dcomp.n23 34.3584
R16981 dcomp.n27 dcomp.n25 34.3584
R16982 dcomp.n29 dcomp.n27 34.3584
R16983 dcomp.n13 dcomp.t26 26.5955
R16984 dcomp.n13 dcomp.t16 26.5955
R16985 dcomp.n0 dcomp.t24 26.5955
R16986 dcomp.n0 dcomp.t31 26.5955
R16987 dcomp.n1 dcomp.t22 26.5955
R16988 dcomp.n1 dcomp.t18 26.5955
R16989 dcomp.n3 dcomp.t21 26.5955
R16990 dcomp.n3 dcomp.t29 26.5955
R16991 dcomp.n5 dcomp.t25 26.5955
R16992 dcomp.n5 dcomp.t28 26.5955
R16993 dcomp.n7 dcomp.t20 26.5955
R16994 dcomp.n7 dcomp.t30 26.5955
R16995 dcomp.n9 dcomp.t23 26.5955
R16996 dcomp.n9 dcomp.t19 26.5955
R16997 dcomp.n11 dcomp.t27 26.5955
R16998 dcomp.n11 dcomp.t17 26.5955
R16999 dcomp.n28 dcomp.t4 24.9236
R17000 dcomp.n28 dcomp.t10 24.9236
R17001 dcomp.n15 dcomp.t2 24.9236
R17002 dcomp.n15 dcomp.t9 24.9236
R17003 dcomp.n16 dcomp.t0 24.9236
R17004 dcomp.n16 dcomp.t12 24.9236
R17005 dcomp.n18 dcomp.t15 24.9236
R17006 dcomp.n18 dcomp.t7 24.9236
R17007 dcomp.n20 dcomp.t3 24.9236
R17008 dcomp.n20 dcomp.t6 24.9236
R17009 dcomp.n22 dcomp.t14 24.9236
R17010 dcomp.n22 dcomp.t8 24.9236
R17011 dcomp.n24 dcomp.t1 24.9236
R17012 dcomp.n24 dcomp.t13 24.9236
R17013 dcomp.n26 dcomp.t5 24.9236
R17014 dcomp.n26 dcomp.t11 24.9236
R17015 dcomp dcomp.n14 18.4247
R17016 dcomp.n30 dcomp.n29 10.0853
R17017 dcomp.n30 dcomp 4.84706
R17018 dcomp.n29 dcomp 1.74595
R17019 dcomp dcomp.n30 1.35808
R17020 schmitt_trigger_0.in.n3 schmitt_trigger_0.in.t2 240.778
R17021 schmitt_trigger_0.in.n0 schmitt_trigger_0.in.t8 240.778
R17022 schmitt_trigger_0.in.n3 schmitt_trigger_0.in.t9 240.349
R17023 schmitt_trigger_0.in.n2 schmitt_trigger_0.in.t4 240.349
R17024 schmitt_trigger_0.in.n1 schmitt_trigger_0.in.t1 240.349
R17025 schmitt_trigger_0.in.n0 schmitt_trigger_0.in.t10 240.349
R17026 schmitt_trigger_0.in.n12 schmitt_trigger_0.in.t3 236.423
R17027 schmitt_trigger_0.in.n12 schmitt_trigger_0.in.t5 236.011
R17028 schmitt_trigger_0.in.n10 schmitt_trigger_0.in.n9 28.545
R17029 schmitt_trigger_0.in.n11 schmitt_trigger_0.in.n10 19.9248
R17030 schmitt_trigger_0.in.n10 schmitt_trigger_0.in.t0 5.93425
R17031 schmitt_trigger_0.in schmitt_trigger_0.in.n12 4.93075
R17032 schmitt_trigger_0.in.n11 schmitt_trigger_0.in.n4 4.72087
R17033 schmitt_trigger_0.in.n1 schmitt_trigger_0.in.n0 0.429848
R17034 schmitt_trigger_0.in.n2 schmitt_trigger_0.in.n1 0.429848
R17035 schmitt_trigger_0.in.n4 schmitt_trigger_0.in.n2 0.285826
R17036 schmitt_trigger_0.in schmitt_trigger_0.in.n11 0.216402
R17037 schmitt_trigger_0.in.n4 schmitt_trigger_0.in.n3 0.0956087
R17038 schmitt_trigger_0.in.n5 schmitt_trigger_0.in.t7 0.0791747
R17039 schmitt_trigger_0.in.n6 schmitt_trigger_0.in.n5 0.06865
R17040 schmitt_trigger_0.in.n7 schmitt_trigger_0.in.n6 0.06865
R17041 schmitt_trigger_0.in.n8 schmitt_trigger_0.in.n7 0.06865
R17042 schmitt_trigger_0.in.n9 schmitt_trigger_0.in.n8 0.06865
R17043 schmitt_trigger_0.in.n5 schmitt_trigger_0.in.t14 0.0110247
R17044 schmitt_trigger_0.in.n6 schmitt_trigger_0.in.t12 0.0110247
R17045 schmitt_trigger_0.in.n7 schmitt_trigger_0.in.t6 0.0110247
R17046 schmitt_trigger_0.in.n8 schmitt_trigger_0.in.t13 0.0110247
R17047 schmitt_trigger_0.in.n9 schmitt_trigger_0.in.t11 0.0110247
R17048 schmitt_trigger_0.m.n5 schmitt_trigger_0.m.t15 240.764
R17049 schmitt_trigger_0.m.n6 schmitt_trigger_0.m.t16 240.713
R17050 schmitt_trigger_0.m.n7 schmitt_trigger_0.m.t17 240.529
R17051 schmitt_trigger_0.m.n5 schmitt_trigger_0.m.t14 240.349
R17052 schmitt_trigger_0.m.n10 schmitt_trigger_0.m.n8 211.214
R17053 schmitt_trigger_0.m.n2 schmitt_trigger_0.m.n0 207.804
R17054 schmitt_trigger_0.m.n2 schmitt_trigger_0.m.n1 207.585
R17055 schmitt_trigger_0.m.n4 schmitt_trigger_0.m.n3 204.175
R17056 schmitt_trigger_0.m.n10 schmitt_trigger_0.m.n9 204.175
R17057 schmitt_trigger_0.m.n13 schmitt_trigger_0.m.n12 70.9014
R17058 schmitt_trigger_0.m.n15 schmitt_trigger_0.m.n14 70.9014
R17059 schmitt_trigger_0.m.n8 schmitt_trigger_0.m.t13 28.5655
R17060 schmitt_trigger_0.m.n8 schmitt_trigger_0.m.t2 28.5655
R17061 schmitt_trigger_0.m.n3 schmitt_trigger_0.m.t8 28.5655
R17062 schmitt_trigger_0.m.n3 schmitt_trigger_0.m.t11 28.5655
R17063 schmitt_trigger_0.m.n1 schmitt_trigger_0.m.t12 28.5655
R17064 schmitt_trigger_0.m.n1 schmitt_trigger_0.m.t10 28.5655
R17065 schmitt_trigger_0.m.n0 schmitt_trigger_0.m.t9 28.5655
R17066 schmitt_trigger_0.m.n0 schmitt_trigger_0.m.t7 28.5655
R17067 schmitt_trigger_0.m.n9 schmitt_trigger_0.m.t1 28.5655
R17068 schmitt_trigger_0.m.n9 schmitt_trigger_0.m.t0 28.5655
R17069 schmitt_trigger_0.m.n12 schmitt_trigger_0.m.t4 17.4005
R17070 schmitt_trigger_0.m.n12 schmitt_trigger_0.m.t3 17.4005
R17071 schmitt_trigger_0.m.n14 schmitt_trigger_0.m.t5 17.4005
R17072 schmitt_trigger_0.m.n14 schmitt_trigger_0.m.t6 17.4005
R17073 schmitt_trigger_0.m.n7 schmitt_trigger_0.m.n6 12.9318
R17074 schmitt_trigger_0.m.n11 schmitt_trigger_0.m.n10 8.3606
R17075 schmitt_trigger_0.m.n4 schmitt_trigger_0.m.n2 3.62811
R17076 schmitt_trigger_0.m schmitt_trigger_0.m.n4 0.819515
R17077 schmitt_trigger_0.m schmitt_trigger_0.m.n15 0.73133
R17078 schmitt_trigger_0.m.n15 schmitt_trigger_0.m.n13 0.688
R17079 schmitt_trigger_0.m.n11 schmitt_trigger_0.m.n7 0.358635
R17080 schmitt_trigger_0.m.n13 schmitt_trigger_0.m.n11 0.251558
R17081 schmitt_trigger_0.m.n6 schmitt_trigger_0.m.n5 0.0297969
R17082 ibias_gen_0.vn0.n9 ibias_gen_0.vn0.t19 50.4613
R17083 ibias_gen_0.vn0.n10 ibias_gen_0.vn0.t19 50.4344
R17084 ibias_gen_0.vn0.n1 ibias_gen_0.vn0.n7 49.6079
R17085 ibias_gen_0.vn0.n4 ibias_gen_0.vn0.t5 49.2687
R17086 ibias_gen_0.vn0.n1 ibias_gen_0.vn0.t5 49.1817
R17087 ibias_gen_0.vn0.t7 ibias_gen_0.vn0.n3 48.1029
R17088 ibias_gen_0.vn0.t20 ibias_gen_0.vn0.n9 48.1029
R17089 ibias_gen_0.vn0.n8 ibias_gen_0.vn0.t7 48.1029
R17090 ibias_gen_0.vn0.n10 ibias_gen_0.vn0.t20 48.1029
R17091 ibias_gen_0.vn0.n0 ibias_gen_0.vn0.t12 22.9447
R17092 ibias_gen_0.Mt4 ibias_gen_0.vn0.n2 21.105
R17093 ibias_gen_0.Mt4 ibias_gen_0.vn0.n15 19.6387
R17094 ibias_gen_0.Mt4 ibias_gen_0.vn0.n14 19.6387
R17095 ibias_gen_0.Mt4 ibias_gen_0.vn0.n13 19.6387
R17096 ibias_gen_0.vn0.n0 ibias_gen_0.vn0.n12 19.6387
R17097 ibias_gen_0.Mt4 ibias_gen_0.vn0.n16 19.6387
R17098 ibias_gen_0.vn0.n6 ibias_gen_0.vn0.n5 13.8791
R17099 ibias_gen_0.vn0.n9 ibias_gen_0.vn0.n8 13.7174
R17100 ibias_gen_0.vn0.n0 ibias_gen_0.vn0.n11 12.7887
R17101 ibias_gen_0.vn0.n11 ibias_gen_0.vn0.n3 7.26784
R17102 ibias_gen_0.vn0.n11 ibias_gen_0.vn0.n10 6.45004
R17103 ibias_gen_0.vn0.n7 ibias_gen_0.vn0.t1 5.5395
R17104 ibias_gen_0.vn0.n7 ibias_gen_0.vn0.t2 5.5395
R17105 ibias_gen_0.vn0.n15 ibias_gen_0.vn0.t11 3.3065
R17106 ibias_gen_0.vn0.n15 ibias_gen_0.vn0.t13 3.3065
R17107 ibias_gen_0.vn0.n14 ibias_gen_0.vn0.t14 3.3065
R17108 ibias_gen_0.vn0.n14 ibias_gen_0.vn0.t16 3.3065
R17109 ibias_gen_0.vn0.n13 ibias_gen_0.vn0.t17 3.3065
R17110 ibias_gen_0.vn0.n13 ibias_gen_0.vn0.t18 3.3065
R17111 ibias_gen_0.vn0.n12 ibias_gen_0.vn0.t9 3.3065
R17112 ibias_gen_0.vn0.n12 ibias_gen_0.vn0.t15 3.3065
R17113 ibias_gen_0.vn0.n5 ibias_gen_0.vn0.t8 3.3065
R17114 ibias_gen_0.vn0.n5 ibias_gen_0.vn0.t6 3.3065
R17115 ibias_gen_0.vn0.n2 ibias_gen_0.vn0.t4 3.3065
R17116 ibias_gen_0.vn0.n2 ibias_gen_0.vn0.t3 3.3065
R17117 ibias_gen_0.vn0.n16 ibias_gen_0.vn0.t0 3.3065
R17118 ibias_gen_0.vn0.n16 ibias_gen_0.vn0.t10 3.3065
R17119 ibias_gen_0.Mt4 ibias_gen_0.vn0.n0 2.11628
R17120 ibias_gen_0.vn0.n6 ibias_gen_0.vn0.n4 1.44615
R17121 ibias_gen_0.vn0.n8 ibias_gen_0.vn0.n1 1.30001
R17122 ibias_gen_0.vn0.n4 ibias_gen_0.vn0.n3 1.16626
R17123 ibias_gen_0.vn0.n1 ibias_gen_0.vn0.n6 1.15267
R17124 ibias_gen_0.vp0.n3 ibias_gen_0.vp0.n1 57.7416
R17125 ibias_gen_0.vp0.n8 ibias_gen_0.vp0.t13 50.9767
R17126 ibias_gen_0.vp0.t13 ibias_gen_0.vp0.n6 50.9767
R17127 ibias_gen_0.vp0.n7 ibias_gen_0.vp0.t6 49.8109
R17128 ibias_gen_0.vp0.n0 ibias_gen_0.vp0.t6 49.7239
R17129 ibias_gen_0.vp0.t8 ibias_gen_0.vp0.n9 48.6451
R17130 ibias_gen_0.vp0.t12 ibias_gen_0.vp0.n6 48.6451
R17131 ibias_gen_0.vp0.n10 ibias_gen_0.vp0.t8 48.6451
R17132 ibias_gen_0.vp0.n8 ibias_gen_0.vp0.t12 48.6451
R17133 ibias_gen_0.vp0.n5 ibias_gen_0.vp0.n4 42.4505
R17134 ibias_gen_0.vp0.n3 ibias_gen_0.vp0.n2 42.4505
R17135 ibias_gen_0.vp0.n14 ibias_gen_0.vp0.n13 18.2113
R17136 ibias_gen_0.vp0.n12 ibias_gen_0.vp0.n11 17.2812
R17137 ibias_gen_0.vp0.n10 ibias_gen_0.vp0.n6 13.7361
R17138 ibias_gen_0.vp0.n9 ibias_gen_0.vp0.n8 13.7361
R17139 ibias_gen_0.vp0.n13 ibias_gen_0.vp0.n12 13.3639
R17140 ibias_gen_0.vp0.n4 ibias_gen_0.vp0.t7 5.5395
R17141 ibias_gen_0.vp0.n4 ibias_gen_0.vp0.t9 5.5395
R17142 ibias_gen_0.vp0.n2 ibias_gen_0.vp0.t5 5.5395
R17143 ibias_gen_0.vp0.n2 ibias_gen_0.vp0.t1 5.5395
R17144 ibias_gen_0.vp0.n1 ibias_gen_0.vp0.t2 5.5395
R17145 ibias_gen_0.vp0.n1 ibias_gen_0.vp0.t4 5.5395
R17146 ibias_gen_0.vp0.n13 ibias_gen_0.vp0.n3 3.97054
R17147 ibias_gen_0.vp0.n12 ibias_gen_0.vp0.n0 3.77198
R17148 ibias_gen_0.vp0.n11 ibias_gen_0.vp0.t11 3.3065
R17149 ibias_gen_0.vp0.n11 ibias_gen_0.vp0.t10 3.3065
R17150 ibias_gen_0.vp0.n14 ibias_gen_0.vp0.t3 3.3065
R17151 ibias_gen_0.vp0.t0 ibias_gen_0.vp0.n14 3.3065
R17152 ibias_gen_0.vp0.n7 ibias_gen_0.vp0.n5 1.47061
R17153 ibias_gen_0.vp0.n0 ibias_gen_0.vp0.n10 1.3293
R17154 ibias_gen_0.vp0.n9 ibias_gen_0.vp0.n7 1.16626
R17155 ibias_gen_0.vp0.n0 ibias_gen_0.vp0.n5 1.13637
R17156 ibias_gen_0.vr.n2 ibias_gen_0.vr.n0 21.7373
R17157 ibias_gen_0.vr.n2 ibias_gen_0.vr.n1 20.4114
R17158 ibias_gen_0.vr.t2 ibias_gen_0.vr.n2 17.6029
R17159 ibias_gen_0.vr.n1 ibias_gen_0.vr.t0 3.3065
R17160 ibias_gen_0.vr.n1 ibias_gen_0.vr.t4 3.3065
R17161 ibias_gen_0.vr.n0 ibias_gen_0.vr.t3 3.3065
R17162 ibias_gen_0.vr.n0 ibias_gen_0.vr.t1 3.3065
R17163 por.n2 por.n0 243.458
R17164 por.n2 por.n1 205.059
R17165 por.n4 por.n3 205.059
R17166 por.n6 por.n5 205.059
R17167 por.n8 por.n7 205.059
R17168 por.n10 por.n9 205.059
R17169 por.n12 por.n11 205.059
R17170 por.n14 por.n13 205.059
R17171 por.n17 por.n15 133.534
R17172 por.n17 por.n16 99.1759
R17173 por.n19 por.n18 99.1759
R17174 por.n21 por.n20 99.1759
R17175 por.n23 por.n22 99.1759
R17176 por.n25 por.n24 99.1759
R17177 por.n27 por.n26 99.1759
R17178 por por.n28 97.4305
R17179 por.n4 por.n2 38.4005
R17180 por.n6 por.n4 38.4005
R17181 por.n8 por.n6 38.4005
R17182 por.n10 por.n8 38.4005
R17183 por.n12 por.n10 38.4005
R17184 por.n14 por.n12 38.4005
R17185 por.n19 por.n17 34.3584
R17186 por.n21 por.n19 34.3584
R17187 por.n23 por.n21 34.3584
R17188 por.n25 por.n23 34.3584
R17189 por.n27 por.n25 34.3584
R17190 por.n29 por.n27 34.3584
R17191 por.n13 por.t31 26.5955
R17192 por.n13 por.t21 26.5955
R17193 por.n0 por.t29 26.5955
R17194 por.n0 por.t20 26.5955
R17195 por.n1 por.t27 26.5955
R17196 por.n1 por.t23 26.5955
R17197 por.n3 por.t26 26.5955
R17198 por.n3 por.t18 26.5955
R17199 por.n5 por.t30 26.5955
R17200 por.n5 por.t17 26.5955
R17201 por.n7 por.t25 26.5955
R17202 por.n7 por.t19 26.5955
R17203 por.n9 por.t28 26.5955
R17204 por.n9 por.t24 26.5955
R17205 por.n11 por.t16 26.5955
R17206 por.n11 por.t22 26.5955
R17207 por.n28 por.t12 24.9236
R17208 por.n28 por.t2 24.9236
R17209 por.n15 por.t10 24.9236
R17210 por.n15 por.t1 24.9236
R17211 por.n16 por.t8 24.9236
R17212 por.n16 por.t4 24.9236
R17213 por.n18 por.t7 24.9236
R17214 por.n18 por.t15 24.9236
R17215 por.n20 por.t11 24.9236
R17216 por.n20 por.t14 24.9236
R17217 por.n22 por.t6 24.9236
R17218 por.n22 por.t0 24.9236
R17219 por.n24 por.t9 24.9236
R17220 por.n24 por.t5 24.9236
R17221 por.n26 por.t13 24.9236
R17222 por.n26 por.t3 24.9236
R17223 por por.n14 18.4247
R17224 por.n30 por.n29 10.0853
R17225 por.n30 por 4.84706
R17226 por.n29 por 1.74595
R17227 por por.n30 1.35808
R17228 porb_h.n2 porb_h.n1 157.593
R17229 porb_h.n43 porb_h.n42 157.591
R17230 porb_h.n38 porb_h.n37 157.591
R17231 porb_h.n32 porb_h.n31 157.591
R17232 porb_h.n26 porb_h.n25 157.591
R17233 porb_h.n20 porb_h.n19 157.591
R17234 porb_h.n14 porb_h.n13 157.591
R17235 porb_h.n8 porb_h.n7 157.591
R17236 porb_h.n43 porb_h.n41 136.965
R17237 porb_h.n38 porb_h.n36 136.965
R17238 porb_h.n32 porb_h.n30 136.965
R17239 porb_h.n26 porb_h.n24 136.965
R17240 porb_h.n20 porb_h.n18 136.965
R17241 porb_h.n14 porb_h.n12 136.965
R17242 porb_h.n8 porb_h.n6 136.965
R17243 porb_h.n2 porb_h.n0 136.965
R17244 porb_h.n41 porb_h.t7 21.2805
R17245 porb_h.n41 porb_h.t15 21.2805
R17246 porb_h.n36 porb_h.t11 21.2805
R17247 porb_h.n36 porb_h.t12 21.2805
R17248 porb_h.n30 porb_h.t13 21.2805
R17249 porb_h.n30 porb_h.t14 21.2805
R17250 porb_h.n24 porb_h.t3 21.2805
R17251 porb_h.n24 porb_h.t0 21.2805
R17252 porb_h.n18 porb_h.t5 21.2805
R17253 porb_h.n18 porb_h.t2 21.2805
R17254 porb_h.n12 porb_h.t8 21.2805
R17255 porb_h.n12 porb_h.t9 21.2805
R17256 porb_h.n6 porb_h.t4 21.2805
R17257 porb_h.n6 porb_h.t10 21.2805
R17258 porb_h.n0 porb_h.t1 21.2805
R17259 porb_h.n0 porb_h.t6 21.2805
R17260 porb_h.n42 porb_h.t18 17.8272
R17261 porb_h.n42 porb_h.t26 17.8272
R17262 porb_h.n37 porb_h.t22 17.8272
R17263 porb_h.n37 porb_h.t23 17.8272
R17264 porb_h.n31 porb_h.t24 17.8272
R17265 porb_h.n31 porb_h.t25 17.8272
R17266 porb_h.n25 porb_h.t30 17.8272
R17267 porb_h.n25 porb_h.t27 17.8272
R17268 porb_h.n19 porb_h.t16 17.8272
R17269 porb_h.n19 porb_h.t29 17.8272
R17270 porb_h.n13 porb_h.t19 17.8272
R17271 porb_h.n13 porb_h.t20 17.8272
R17272 porb_h.n7 porb_h.t31 17.8272
R17273 porb_h.n7 porb_h.t21 17.8272
R17274 porb_h.n1 porb_h.t28 17.8272
R17275 porb_h.n1 porb_h.t17 17.8272
R17276 porb_h.n44 porb_h.n43 10.1618
R17277 porb_h.n3 porb_h.n2 9.98018
R17278 porb_h.n39 porb_h.n38 9.98018
R17279 porb_h.n33 porb_h.n32 9.98018
R17280 porb_h.n27 porb_h.n26 9.98018
R17281 porb_h.n21 porb_h.n20 9.98018
R17282 porb_h.n15 porb_h.n14 9.98018
R17283 porb_h.n9 porb_h.n8 9.98018
R17284 porb_h.n40 porb_h 7.09609
R17285 porb_h.n34 porb_h 5.94903
R17286 porb_h.n35 porb_h 5.08746
R17287 porb_h.n28 porb_h 4.80197
R17288 porb_h.n29 porb_h 4.23963
R17289 porb_h porb_h.n45 3.88917
R17290 porb_h.n22 porb_h 3.65491
R17291 porb_h.n23 porb_h 3.3918
R17292 porb_h.n17 porb_h 2.54398
R17293 porb_h.n16 porb_h 2.50785
R17294 porb_h.n11 porb_h 1.69615
R17295 porb_h.n44 porb_h 1.37745
R17296 porb_h.n10 porb_h 1.36079
R17297 porb_h.n5 porb_h.n4 0.934324
R17298 porb_h.n11 porb_h.n10 0.934324
R17299 porb_h.n17 porb_h.n16 0.934324
R17300 porb_h.n23 porb_h.n22 0.934324
R17301 porb_h.n29 porb_h.n28 0.934324
R17302 porb_h.n35 porb_h.n34 0.934324
R17303 porb_h.n5 porb_h 0.848326
R17304 porb_h.n45 porb_h.n44 0.252453
R17305 porb_h.n45 porb_h.n40 0.224765
R17306 porb_h.n4 porb_h 0.213735
R17307 porb_h.n4 porb_h.n3 0.0793043
R17308 porb_h.n3 porb_h 0.0793043
R17309 porb_h.n10 porb_h.n9 0.0793043
R17310 porb_h.n9 porb_h.n5 0.0793043
R17311 porb_h.n16 porb_h.n15 0.0793043
R17312 porb_h.n15 porb_h.n11 0.0793043
R17313 porb_h.n22 porb_h.n21 0.0793043
R17314 porb_h.n21 porb_h.n17 0.0793043
R17315 porb_h.n28 porb_h.n27 0.0793043
R17316 porb_h.n27 porb_h.n23 0.0793043
R17317 porb_h.n34 porb_h.n33 0.0793043
R17318 porb_h.n33 porb_h.n29 0.0793043
R17319 porb_h.n40 porb_h.n39 0.0793043
R17320 porb_h.n39 porb_h.n35 0.0793043
R17321 ibias_gen_0.vp.n10 ibias_gen_0.vp.t4 56.5501
R17322 ibias_gen_0.vp.n4 ibias_gen_0.vp.t11 50.9767
R17323 ibias_gen_0.vp.n5 ibias_gen_0.vp.t11 50.9767
R17324 ibias_gen_0.vp.t9 ibias_gen_0.vp.n6 50.9767
R17325 ibias_gen_0.vp.t8 ibias_gen_0.vp.n4 48.6451
R17326 ibias_gen_0.vp.n7 ibias_gen_0.vp.t9 48.6451
R17327 ibias_gen_0.vp.n6 ibias_gen_0.vp.t7 48.6451
R17328 ibias_gen_0.vp.n5 ibias_gen_0.vp.t8 48.6451
R17329 ibias_gen_0.vp.t7 ibias_gen_0.vp.n3 48.6451
R17330 ibias_gen_0.vp.n0 ibias_gen_0.vp.n11 42.5266
R17331 ibias_gen_0.vp.n0 ibias_gen_0.vp.n2 42.4505
R17332 ibias_gen_0.vp.n9 ibias_gen_0.vp.n8 26.1532
R17333 ibias_gen_0.vp.n8 ibias_gen_0.vp.t12 25.4891
R17334 ibias_gen_0.vp.n8 ibias_gen_0.vp.t10 24.3233
R17335 ibias_gen_0.vp.n13 ibias_gen_0.vp.n12 15.1165
R17336 ibias_gen_0.vp.n12 ibias_gen_0.vp.n1 14.8365
R17337 ibias_gen_0.vp.n10 ibias_gen_0.vp.n9 8.08875
R17338 ibias_gen_0.vp.n12 ibias_gen_0.vp.n0 7.57893
R17339 ibias_gen_0.vp.n0 ibias_gen_0.vp.n10 6.28836
R17340 ibias_gen_0.vp.n2 ibias_gen_0.vp.t2 5.5395
R17341 ibias_gen_0.vp.t1 ibias_gen_0.vp.n2 5.5395
R17342 ibias_gen_0.vp.n11 ibias_gen_0.vp.t1 5.5395
R17343 ibias_gen_0.vp.n11 ibias_gen_0.vp.t6 5.5395
R17344 ibias_gen_0.vp.n1 ibias_gen_0.vp.t5 3.3065
R17345 ibias_gen_0.vp.t0 ibias_gen_0.vp.n1 3.3065
R17346 ibias_gen_0.vp.t0 ibias_gen_0.vp.n13 3.3065
R17347 ibias_gen_0.vp.n13 ibias_gen_0.vp.t3 3.3065
R17348 ibias_gen_0.vp.n9 ibias_gen_0.vp.n7 2.37524
R17349 ibias_gen_0.vp.n6 ibias_gen_0.vp.n5 2.33202
R17350 ibias_gen_0.vp.n4 ibias_gen_0.vp.n3 2.33202
R17351 ibias_gen_0.vp.n7 ibias_gen_0.vp.n3 2.33126
R17352 itest itest.n0 45.907
R17353 itest.n0 itest.t0 5.5395
R17354 itest.n0 itest.t1 5.5395
R17355 rstring_mux_0.vtrip7.n5 rstring_mux_0.vtrip7.n3 50.7022
R17356 rstring_mux_0.vtrip7.n2 rstring_mux_0.vtrip7.n0 50.7022
R17357 rstring_mux_0.vtrip7.n6 rstring_mux_0.vtrip7.n5 15.3935
R17358 rstring_mux_0.vtrip7.n5 rstring_mux_0.vtrip7.n4 13.8791
R17359 rstring_mux_0.vtrip7.n2 rstring_mux_0.vtrip7.n1 13.8791
R17360 rstring_mux_0.vtrip7.t0 rstring_mux_0.vtrip7.n7 10.5857
R17361 rstring_mux_0.vtrip7.n7 rstring_mux_0.vtrip7.t7 10.5847
R17362 rstring_mux_0.vtrip7.n3 rstring_mux_0.vtrip7.t9 5.5395
R17363 rstring_mux_0.vtrip7.n3 rstring_mux_0.vtrip7.t8 5.5395
R17364 rstring_mux_0.vtrip7.n0 rstring_mux_0.vtrip7.t1 5.5395
R17365 rstring_mux_0.vtrip7.n0 rstring_mux_0.vtrip7.t2 5.5395
R17366 rstring_mux_0.vtrip7.n6 rstring_mux_0.vtrip7.n2 5.2741
R17367 rstring_mux_0.vtrip7.n4 rstring_mux_0.vtrip7.t5 3.3065
R17368 rstring_mux_0.vtrip7.n4 rstring_mux_0.vtrip7.t6 3.3065
R17369 rstring_mux_0.vtrip7.n1 rstring_mux_0.vtrip7.t3 3.3065
R17370 rstring_mux_0.vtrip7.n1 rstring_mux_0.vtrip7.t4 3.3065
R17371 rstring_mux_0.vtrip7.n7 rstring_mux_0.vtrip7.n6 2.48711
R17372 rstring_mux_0.vtrip2.n5 rstring_mux_0.vtrip2.n3 50.7022
R17373 rstring_mux_0.vtrip2.n2 rstring_mux_0.vtrip2.n0 50.7022
R17374 rstring_mux_0.vtrip2.n7 rstring_mux_0.vtrip2.n6 23.8383
R17375 rstring_mux_0.vtrip2.n6 rstring_mux_0.vtrip2.n5 14.3726
R17376 rstring_mux_0.vtrip2.n5 rstring_mux_0.vtrip2.n4 13.8791
R17377 rstring_mux_0.vtrip2.n2 rstring_mux_0.vtrip2.n1 13.8791
R17378 rstring_mux_0.vtrip2 rstring_mux_0.vtrip2.t3 10.5739
R17379 rstring_mux_0.vtrip2.n3 rstring_mux_0.vtrip2.t2 5.5395
R17380 rstring_mux_0.vtrip2.n3 rstring_mux_0.vtrip2.t1 5.5395
R17381 rstring_mux_0.vtrip2.n0 rstring_mux_0.vtrip2.t8 5.5395
R17382 rstring_mux_0.vtrip2.n0 rstring_mux_0.vtrip2.t9 5.5395
R17383 rstring_mux_0.vtrip2.n6 rstring_mux_0.vtrip2.n2 4.21994
R17384 rstring_mux_0.vtrip2.n4 rstring_mux_0.vtrip2.t6 3.3065
R17385 rstring_mux_0.vtrip2.n4 rstring_mux_0.vtrip2.t7 3.3065
R17386 rstring_mux_0.vtrip2.n1 rstring_mux_0.vtrip2.t5 3.3065
R17387 rstring_mux_0.vtrip2.n1 rstring_mux_0.vtrip2.t4 3.3065
R17388 rstring_mux_0.vtrip2.n7 rstring_mux_0.vtrip2.t0 0.826075
R17389 rstring_mux_0.vtrip2 rstring_mux_0.vtrip2.n7 0.0563195
R17390 ibias_gen_0.vp1.n5 ibias_gen_0.vp1.n4 53.0003
R17391 ibias_gen_0.vp1.t13 ibias_gen_0.vp1.n3 49.8109
R17392 ibias_gen_0.vp1.n3 ibias_gen_0.vp1.t11 49.8109
R17393 ibias_gen_0.vp1.t11 ibias_gen_0.vp1.n0 49.7878
R17394 ibias_gen_0.vp1.n0 ibias_gen_0.vp1.t13 49.6053
R17395 ibias_gen_0.vp1 ibias_gen_0.vp1.n6 45.7548
R17396 ibias_gen_0.vp1.n2 ibias_gen_0.vp1.n1 42.4505
R17397 ibias_gen_0.vp1.n9 ibias_gen_0.vp1.n7 18.5825
R17398 ibias_gen_0.vp1.n15 ibias_gen_0.vp1.n14 17.1535
R17399 ibias_gen_0.vp1.n11 ibias_gen_0.vp1.n10 16.3247
R17400 ibias_gen_0.vp1.n9 ibias_gen_0.vp1.n8 16.3247
R17401 ibias_gen_0.vp1.n13 ibias_gen_0.vp1.n12 15.5548
R17402 ibias_gen_0.vp1.n15 ibias_gen_0.vp1.n13 11.684
R17403 ibias_gen_0.vp1.n6 ibias_gen_0.vp1.t9 5.5395
R17404 ibias_gen_0.vp1.n6 ibias_gen_0.vp1.t10 5.5395
R17405 ibias_gen_0.vp1.n4 ibias_gen_0.vp1.t15 5.5395
R17406 ibias_gen_0.vp1.n4 ibias_gen_0.vp1.t17 5.5395
R17407 ibias_gen_0.vp1.n1 ibias_gen_0.vp1.t12 5.5395
R17408 ibias_gen_0.vp1.n1 ibias_gen_0.vp1.t14 5.5395
R17409 ibias_gen_0.vp1.n5 ibias_gen_0.vp1.n0 4.85318
R17410 ibias_gen_0.vp1.n11 ibias_gen_0.vp1.n9 4.51612
R17411 ibias_gen_0.vp1.n12 ibias_gen_0.vp1.t5 3.3065
R17412 ibias_gen_0.vp1.n12 ibias_gen_0.vp1.t0 3.3065
R17413 ibias_gen_0.vp1.n10 ibias_gen_0.vp1.t7 3.3065
R17414 ibias_gen_0.vp1.n10 ibias_gen_0.vp1.t4 3.3065
R17415 ibias_gen_0.vp1.n8 ibias_gen_0.vp1.t3 3.3065
R17416 ibias_gen_0.vp1.n8 ibias_gen_0.vp1.t6 3.3065
R17417 ibias_gen_0.vp1.n7 ibias_gen_0.vp1.t1 3.3065
R17418 ibias_gen_0.vp1.n7 ibias_gen_0.vp1.t2 3.3065
R17419 ibias_gen_0.vp1.n14 ibias_gen_0.vp1.t8 3.3065
R17420 ibias_gen_0.vp1.n14 ibias_gen_0.vp1.t16 3.3065
R17421 ibias_gen_0.vp1.n13 ibias_gen_0.vp1.n11 2.27562
R17422 ibias_gen_0.vp1 ibias_gen_0.vp1.n15 1.87819
R17423 ibias_gen_0.vp1.n2 ibias_gen_0.vp1.n0 1.48628
R17424 ibias_gen_0.vp1.n3 ibias_gen_0.vp1.n2 1.47061
R17425 ibias_gen_0.vp1 ibias_gen_0.vp1.n5 1.36236
R17426 ibias_gen_0.vn1.n0 ibias_gen_0.vn1.n1 47.4959
R17427 ibias_gen_0.vn1.n3 ibias_gen_0.vn1.t14 27.5855
R17428 ibias_gen_0.vn1.n2 ibias_gen_0.vn1.t10 27.5855
R17429 ibias_gen_0.vn1.n6 ibias_gen_0.vn1.t16 27.5855
R17430 ibias_gen_0.vn1.n5 ibias_gen_0.vn1.t12 27.5855
R17431 ibias_gen_0.vn1.n10 ibias_gen_0.vn1.t2 26.004
R17432 ibias_gen_0.vn1.n0 ibias_gen_0.vn1.n13 24.5059
R17433 ibias_gen_0.vn1.n3 ibias_gen_0.vn1.t17 24.3247
R17434 ibias_gen_0.vn1.n2 ibias_gen_0.vn1.t15 24.3247
R17435 ibias_gen_0.vn1.n6 ibias_gen_0.vn1.t13 24.3247
R17436 ibias_gen_0.vn1.n5 ibias_gen_0.vn1.t11 24.3247
R17437 ibias_gen_0.vn1.n9 ibias_gen_0.vn1.t0 24.3247
R17438 ibias_gen_0.vn1.n14 ibias_gen_0.vn1.n0 17.1535
R17439 ibias_gen_0.vn1.n12 ibias_gen_0.vn1.n11 13.8791
R17440 ibias_gen_0.vn1.n0 ibias_gen_0.vn1.n12 12.7397
R17441 ibias_gen_0.vn1.n1 ibias_gen_0.vn1.t7 5.5395
R17442 ibias_gen_0.vn1.n1 ibias_gen_0.vn1.t5 5.5395
R17443 ibias_gen_0.vn1.n4 ibias_gen_0.vn1.n2 4.66645
R17444 ibias_gen_0.vn1.n7 ibias_gen_0.vn1.n5 4.66645
R17445 ibias_gen_0.vn1.n13 ibias_gen_0.vn1.t8 3.3065
R17446 ibias_gen_0.vn1.n13 ibias_gen_0.vn1.t6 3.3065
R17447 ibias_gen_0.vn1.n11 ibias_gen_0.vn1.t1 3.3065
R17448 ibias_gen_0.vn1.n11 ibias_gen_0.vn1.t3 3.3065
R17449 ibias_gen_0.vn1.n14 ibias_gen_0.vn1.t9 3.3065
R17450 ibias_gen_0.vn1.t4 ibias_gen_0.vn1.n14 3.3065
R17451 ibias_gen_0.vn1.n8 ibias_gen_0.vn1.n4 2.41645
R17452 ibias_gen_0.vn1.n8 ibias_gen_0.vn1.n7 2.41645
R17453 ibias_gen_0.vn1.n4 ibias_gen_0.vn1.n3 2.2505
R17454 ibias_gen_0.vn1.n7 ibias_gen_0.vn1.n6 2.2505
R17455 ibias_gen_0.vn1.n9 ibias_gen_0.vn1.n8 2.2505
R17456 ibias_gen_0.vn1.n10 ibias_gen_0.vn1.n9 1.58202
R17457 ibias_gen_0.vn1.n12 ibias_gen_0.vn1.n10 1.37822
R17458 por_unbuf.n15 por_unbuf.t7 212.081
R17459 por_unbuf.n17 por_unbuf.t3 212.081
R17460 por_unbuf.n14 por_unbuf.t12 212.081
R17461 por_unbuf.n22 por_unbuf.t2 212.081
R17462 por_unbuf.n2 por_unbuf.t9 212.081
R17463 por_unbuf.n1 por_unbuf.t6 212.081
R17464 por_unbuf.n6 por_unbuf.t14 212.081
R17465 por_unbuf.n8 por_unbuf.t4 212.081
R17466 por_unbuf.n23 por_unbuf.n22 188.516
R17467 por_unbuf.n9 por_unbuf.n8 188.516
R17468 por_unbuf.n10 por_unbuf.t5 186.374
R17469 por_unbuf.n10 por_unbuf.t15 170.308
R17470 por_unbuf.n11 por_unbuf 155.511
R17471 por_unbuf.n16 por_unbuf 154.304
R17472 por_unbuf por_unbuf.n3 154.304
R17473 por_unbuf.n12 por_unbuf.n11 153.462
R17474 por_unbuf.n21 por_unbuf.n20 152
R17475 por_unbuf.n19 por_unbuf.n18 152
R17476 por_unbuf.n7 por_unbuf.n0 152
R17477 por_unbuf.n5 por_unbuf.n4 152
R17478 por_unbuf.n15 por_unbuf.t16 139.78
R17479 por_unbuf.n17 por_unbuf.t11 139.78
R17480 por_unbuf.n14 por_unbuf.t0 139.78
R17481 por_unbuf.n22 por_unbuf.t8 139.78
R17482 por_unbuf.n2 por_unbuf.t17 139.78
R17483 por_unbuf.n1 por_unbuf.t13 139.78
R17484 por_unbuf.n6 por_unbuf.t1 139.78
R17485 por_unbuf.n8 por_unbuf.t10 139.78
R17486 por_unbuf.n11 por_unbuf.n10 101.513
R17487 por_unbuf.n16 por_unbuf.n15 30.6732
R17488 por_unbuf.n17 por_unbuf.n16 30.6732
R17489 por_unbuf.n18 por_unbuf.n17 30.6732
R17490 por_unbuf.n18 por_unbuf.n14 30.6732
R17491 por_unbuf.n21 por_unbuf.n14 30.6732
R17492 por_unbuf.n22 por_unbuf.n21 30.6732
R17493 por_unbuf.n3 por_unbuf.n2 30.6732
R17494 por_unbuf.n3 por_unbuf.n1 30.6732
R17495 por_unbuf.n5 por_unbuf.n1 30.6732
R17496 por_unbuf.n6 por_unbuf.n5 30.6732
R17497 por_unbuf.n7 por_unbuf.n6 30.6732
R17498 por_unbuf.n8 por_unbuf.n7 30.6732
R17499 por_unbuf.n26 por_unbuf.n13 25.3344
R17500 por_unbuf.n27 por_unbuf.n26 20.7505
R17501 por_unbuf.n19 por_unbuf 19.2005
R17502 por_unbuf.n4 por_unbuf 19.2005
R17503 por_unbuf.n20 por_unbuf 17.1525
R17504 por_unbuf por_unbuf.n0 17.1525
R17505 por_unbuf.n26 por_unbuf.n25 14.6677
R17506 por_unbuf por_unbuf.n27 12.5445
R17507 por_unbuf.n24 por_unbuf.n23 10.4965
R17508 por_unbuf.n25 por_unbuf.n24 6.90245
R17509 por_unbuf.n24 por_unbuf 6.6565
R17510 por_unbuf.n20 por_unbuf 6.4005
R17511 por_unbuf.n23 por_unbuf 6.4005
R17512 por_unbuf por_unbuf.n0 6.4005
R17513 por_unbuf.n9 por_unbuf 6.4005
R17514 por_unbuf.n13 por_unbuf.n12 5.9876
R17515 por_unbuf.n12 por_unbuf 4.74889
R17516 por_unbuf.n27 por_unbuf.n9 4.6085
R17517 por_unbuf.n13 por_unbuf 4.54244
R17518 por_unbuf por_unbuf.n19 4.3525
R17519 por_unbuf.n4 por_unbuf 4.3525
R17520 por_unbuf.n25 por_unbuf 0.172375
R17521 osc_ena.n1 osc_ena.t3 413.582
R17522 osc_ena.n0 osc_ena.t0 348.789
R17523 osc_ena.n1 osc_ena.t1 227.718
R17524 osc_ena.n0 osc_ena.t2 224.327
R17525 osc_ena.n2 osc_ena.n0 13.8663
R17526 osc_ena.n2 osc_ena.n1 4.5005
R17527 osc_ena osc_ena.n2 0.0755
R17528 rstring_mux_0.vtrip3.n5 rstring_mux_0.vtrip3.n3 50.7022
R17529 rstring_mux_0.vtrip3.n2 rstring_mux_0.vtrip3.n0 50.7022
R17530 rstring_mux_0.vtrip3.n6 rstring_mux_0.vtrip3.n5 14.2209
R17531 rstring_mux_0.vtrip3.n5 rstring_mux_0.vtrip3.n4 13.8791
R17532 rstring_mux_0.vtrip3.n2 rstring_mux_0.vtrip3.n1 13.8791
R17533 rstring_mux_0.vtrip3.t0 rstring_mux_0.vtrip3.n7 10.5857
R17534 rstring_mux_0.vtrip3.n7 rstring_mux_0.vtrip3.t5 10.5847
R17535 rstring_mux_0.vtrip3.n6 rstring_mux_0.vtrip3.n2 5.7125
R17536 rstring_mux_0.vtrip3.n3 rstring_mux_0.vtrip3.t8 5.5395
R17537 rstring_mux_0.vtrip3.n3 rstring_mux_0.vtrip3.t9 5.5395
R17538 rstring_mux_0.vtrip3.n0 rstring_mux_0.vtrip3.t3 5.5395
R17539 rstring_mux_0.vtrip3.n0 rstring_mux_0.vtrip3.t4 5.5395
R17540 rstring_mux_0.vtrip3.n4 rstring_mux_0.vtrip3.t2 3.3065
R17541 rstring_mux_0.vtrip3.n4 rstring_mux_0.vtrip3.t1 3.3065
R17542 rstring_mux_0.vtrip3.n1 rstring_mux_0.vtrip3.t6 3.3065
R17543 rstring_mux_0.vtrip3.n1 rstring_mux_0.vtrip3.t7 3.3065
R17544 rstring_mux_0.vtrip3.n7 rstring_mux_0.vtrip3.n6 3.16869
R17545 ibias_gen_0.vstart.n0 ibias_gen_0.vstart.t0 56.685
R17546 ibias_gen_0.vstart.n5 ibias_gen_0.vstart.n3 20.328
R17547 ibias_gen_0.vstart.n0 ibias_gen_0.vstart.n1 20.2356
R17548 ibias_gen_0.vstart.n5 ibias_gen_0.vstart.n4 20.069
R17549 ibias_gen_0.vstart.n0 ibias_gen_0.vstart.n2 20.069
R17550 ibias_gen_0.vstart.n7 ibias_gen_0.vstart.n6 20.069
R17551 ibias_gen_0.vstart.n4 ibias_gen_0.vstart.t10 3.3065
R17552 ibias_gen_0.vstart.n4 ibias_gen_0.vstart.t1 3.3065
R17553 ibias_gen_0.vstart.n3 ibias_gen_0.vstart.t7 3.3065
R17554 ibias_gen_0.vstart.n3 ibias_gen_0.vstart.t4 3.3065
R17555 ibias_gen_0.vstart.n2 ibias_gen_0.vstart.t5 3.3065
R17556 ibias_gen_0.vstart.n2 ibias_gen_0.vstart.t6 3.3065
R17557 ibias_gen_0.vstart.n1 ibias_gen_0.vstart.t2 3.3065
R17558 ibias_gen_0.vstart.n1 ibias_gen_0.vstart.t3 3.3065
R17559 ibias_gen_0.vstart.n7 ibias_gen_0.vstart.t8 3.3065
R17560 ibias_gen_0.vstart.t9 ibias_gen_0.vstart.n7 3.3065
R17561 ibias_gen_0.vstart.n6 ibias_gen_0.vstart.n0 0.280933
R17562 ibias_gen_0.vstart.n6 ibias_gen_0.vstart.n5 0.2449
R17563 schmitt_trigger_0.out.n8 schmitt_trigger_0.out.t12 248.236
R17564 schmitt_trigger_0.out.n6 schmitt_trigger_0.out.t11 240.778
R17565 schmitt_trigger_0.out.n7 schmitt_trigger_0.out.t4 240.613
R17566 schmitt_trigger_0.out.n6 schmitt_trigger_0.out.t5 240.349
R17567 schmitt_trigger_0.out.n5 schmitt_trigger_0.out.t2 236.369
R17568 schmitt_trigger_0.out.n0 schmitt_trigger_0.out.t8 212.081
R17569 schmitt_trigger_0.out.n2 schmitt_trigger_0.out.t7 212.081
R17570 schmitt_trigger_0.out.n15 schmitt_trigger_0.out.t13 212.081
R17571 schmitt_trigger_0.out.n3 schmitt_trigger_0.out.t6 212.081
R17572 schmitt_trigger_0.out.n5 schmitt_trigger_0.out.n4 207.585
R17573 schmitt_trigger_0.out.n12 schmitt_trigger_0.out.n3 188.516
R17574 sky130_fd_sc_hd__inv_4_0.A schmitt_trigger_0.out.n1 154.304
R17575 schmitt_trigger_0.out.n14 schmitt_trigger_0.out.n13 152
R17576 schmitt_trigger_0.out.n17 schmitt_trigger_0.out.n16 152
R17577 schmitt_trigger_0.out.n0 schmitt_trigger_0.out.t14 139.78
R17578 schmitt_trigger_0.out.n2 schmitt_trigger_0.out.t10 139.78
R17579 schmitt_trigger_0.out.n15 schmitt_trigger_0.out.t15 139.78
R17580 schmitt_trigger_0.out.n3 schmitt_trigger_0.out.t9 139.78
R17581 schmitt_trigger_0.out.n10 schmitt_trigger_0.out.t0 91.727
R17582 schmitt_trigger_0.out.n1 schmitt_trigger_0.out.n0 30.6732
R17583 schmitt_trigger_0.out.n2 schmitt_trigger_0.out.n1 30.6732
R17584 schmitt_trigger_0.out.n16 schmitt_trigger_0.out.n2 30.6732
R17585 schmitt_trigger_0.out.n16 schmitt_trigger_0.out.n15 30.6732
R17586 schmitt_trigger_0.out.n15 schmitt_trigger_0.out.n14 30.6732
R17587 schmitt_trigger_0.out.n14 schmitt_trigger_0.out.n3 30.6732
R17588 schmitt_trigger_0.out.n4 schmitt_trigger_0.out.t3 28.5655
R17589 schmitt_trigger_0.out.n4 schmitt_trigger_0.out.t1 28.5655
R17590 schmitt_trigger_0.out.n11 schmitt_trigger_0.out.n10 20.1312
R17591 sky130_fd_sc_hd__inv_4_0.A schmitt_trigger_0.out.n17 19.2005
R17592 sky130_fd_sc_hd__inv_4_0.A schmitt_trigger_0.out.n12 17.1525
R17593 schmitt_trigger_0.out.n11 sky130_fd_sc_hd__inv_4_0.A 12.8005
R17594 schmitt_trigger_0.out.n9 schmitt_trigger_0.out.n5 8.66251
R17595 schmitt_trigger_0.out.n13 sky130_fd_sc_hd__inv_4_0.A 6.4005
R17596 schmitt_trigger_0.out.n12 sky130_fd_sc_hd__inv_4_0.A 6.4005
R17597 schmitt_trigger_0.out.n8 schmitt_trigger_0.out.n7 4.94425
R17598 schmitt_trigger_0.out.n17 sky130_fd_sc_hd__inv_4_0.A 4.3525
R17599 schmitt_trigger_0.out.n13 schmitt_trigger_0.out.n11 4.3525
R17600 schmitt_trigger_0.out.n9 schmitt_trigger_0.out.n8 4.05633
R17601 schmitt_trigger_0.out.n10 schmitt_trigger_0.out.n9 0.230017
R17602 schmitt_trigger_0.out.n7 schmitt_trigger_0.out.n6 0.117348
R17603 otrip_decoded[6].n0 otrip_decoded[6].t0 186.374
R17604 otrip_decoded[6].n0 otrip_decoded[6].t1 170.308
R17605 otrip_decoded[6] otrip_decoded[6].n1 154.56
R17606 otrip_decoded[6].n2 otrip_decoded[6].n1 153.462
R17607 otrip_decoded[6].n1 otrip_decoded[6].n0 101.513
R17608 otrip_decoded[6].n3 otrip_decoded[6] 11.8005
R17609 otrip_decoded[6].n3 otrip_decoded[6].n2 4.96991
R17610 otrip_decoded[6].n2 otrip_decoded[6] 3.46403
R17611 otrip_decoded[6] otrip_decoded[6].n3 2.71109
R17612 rstring_mux_0.vtrip5.n5 rstring_mux_0.vtrip5.n3 50.7022
R17613 rstring_mux_0.vtrip5.n2 rstring_mux_0.vtrip5.n0 50.7022
R17614 rstring_mux_0.vtrip5.n6 rstring_mux_0.vtrip5.n2 14.7069
R17615 rstring_mux_0.vtrip5.n5 rstring_mux_0.vtrip5.n4 13.8791
R17616 rstring_mux_0.vtrip5.n2 rstring_mux_0.vtrip5.n1 13.8791
R17617 rstring_mux_0.vtrip5.t0 rstring_mux_0.vtrip5.n7 10.5857
R17618 rstring_mux_0.vtrip5.n7 rstring_mux_0.vtrip5.t9 10.5847
R17619 rstring_mux_0.vtrip5.n3 rstring_mux_0.vtrip5.t1 5.5395
R17620 rstring_mux_0.vtrip5.n3 rstring_mux_0.vtrip5.t2 5.5395
R17621 rstring_mux_0.vtrip5.n0 rstring_mux_0.vtrip5.t6 5.5395
R17622 rstring_mux_0.vtrip5.n0 rstring_mux_0.vtrip5.t5 5.5395
R17623 rstring_mux_0.vtrip5.n7 rstring_mux_0.vtrip5.n6 5.07153
R17624 rstring_mux_0.vtrip5.n6 rstring_mux_0.vtrip5.n5 3.33746
R17625 rstring_mux_0.vtrip5.n4 rstring_mux_0.vtrip5.t7 3.3065
R17626 rstring_mux_0.vtrip5.n4 rstring_mux_0.vtrip5.t8 3.3065
R17627 rstring_mux_0.vtrip5.n1 rstring_mux_0.vtrip5.t4 3.3065
R17628 rstring_mux_0.vtrip5.n1 rstring_mux_0.vtrip5.t3 3.3065
R17629 otrip_decoded[4].n0 otrip_decoded[4].t0 186.374
R17630 otrip_decoded[4].n0 otrip_decoded[4].t1 170.308
R17631 otrip_decoded[4] otrip_decoded[4].n1 154.56
R17632 otrip_decoded[4].n2 otrip_decoded[4].n1 153.462
R17633 otrip_decoded[4].n1 otrip_decoded[4].n0 101.513
R17634 otrip_decoded[4].n3 otrip_decoded[4] 11.8005
R17635 otrip_decoded[4].n3 otrip_decoded[4].n2 4.96991
R17636 otrip_decoded[4].n2 otrip_decoded[4] 3.46403
R17637 otrip_decoded[4] otrip_decoded[4].n3 2.71109
R17638 rstring_mux_0.vtrip1.n5 rstring_mux_0.vtrip1.n3 50.7022
R17639 rstring_mux_0.vtrip1.n2 rstring_mux_0.vtrip1.n0 50.7022
R17640 rstring_mux_0.vtrip1.n6 rstring_mux_0.vtrip1.n5 14.0767
R17641 rstring_mux_0.vtrip1.n5 rstring_mux_0.vtrip1.n4 13.8791
R17642 rstring_mux_0.vtrip1.n2 rstring_mux_0.vtrip1.n1 13.8791
R17643 rstring_mux_0.vtrip1.t2 rstring_mux_0.vtrip1.n7 10.5857
R17644 rstring_mux_0.vtrip1.n7 rstring_mux_0.vtrip1.t3 10.5847
R17645 rstring_mux_0.vtrip1.n7 rstring_mux_0.vtrip1.n6 5.61984
R17646 rstring_mux_0.vtrip1.n3 rstring_mux_0.vtrip1.t5 5.5395
R17647 rstring_mux_0.vtrip1.n3 rstring_mux_0.vtrip1.t4 5.5395
R17648 rstring_mux_0.vtrip1.n0 rstring_mux_0.vtrip1.t7 5.5395
R17649 rstring_mux_0.vtrip1.n0 rstring_mux_0.vtrip1.t6 5.5395
R17650 rstring_mux_0.vtrip1.n6 rstring_mux_0.vtrip1.n2 3.9186
R17651 rstring_mux_0.vtrip1.n4 rstring_mux_0.vtrip1.t0 3.3065
R17652 rstring_mux_0.vtrip1.n4 rstring_mux_0.vtrip1.t1 3.3065
R17653 rstring_mux_0.vtrip1.n1 rstring_mux_0.vtrip1.t9 3.3065
R17654 rstring_mux_0.vtrip1.n1 rstring_mux_0.vtrip1.t8 3.3065
R17655 otrip_decoded[2].n0 otrip_decoded[2].t0 186.374
R17656 otrip_decoded[2].n0 otrip_decoded[2].t1 170.308
R17657 otrip_decoded[2] otrip_decoded[2].n1 154.56
R17658 otrip_decoded[2].n2 otrip_decoded[2].n1 153.462
R17659 otrip_decoded[2].n1 otrip_decoded[2].n0 101.513
R17660 otrip_decoded[2].n3 otrip_decoded[2] 11.8005
R17661 otrip_decoded[2].n3 otrip_decoded[2].n2 4.96991
R17662 otrip_decoded[2].n2 otrip_decoded[2] 3.46403
R17663 otrip_decoded[2] otrip_decoded[2].n3 2.71109
R17664 rstring_mux_0.vtrip6.n5 rstring_mux_0.vtrip6.n3 50.7022
R17665 rstring_mux_0.vtrip6.n2 rstring_mux_0.vtrip6.n0 50.7022
R17666 rstring_mux_0.vtrip6.n7 rstring_mux_0.vtrip6.n6 21.6754
R17667 rstring_mux_0.vtrip6.n6 rstring_mux_0.vtrip6.n5 14.944
R17668 rstring_mux_0.vtrip6.n5 rstring_mux_0.vtrip6.n4 13.8791
R17669 rstring_mux_0.vtrip6.n2 rstring_mux_0.vtrip6.n1 13.8791
R17670 rstring_mux_0.vtrip6.n7 rstring_mux_0.vtrip6.t9 10.6303
R17671 rstring_mux_0.vtrip6.n3 rstring_mux_0.vtrip6.t2 5.5395
R17672 rstring_mux_0.vtrip6.n3 rstring_mux_0.vtrip6.t1 5.5395
R17673 rstring_mux_0.vtrip6.n0 rstring_mux_0.vtrip6.t6 5.5395
R17674 rstring_mux_0.vtrip6.n0 rstring_mux_0.vtrip6.t5 5.5395
R17675 rstring_mux_0.vtrip6.n6 rstring_mux_0.vtrip6.n2 5.01904
R17676 rstring_mux_0.vtrip6.n4 rstring_mux_0.vtrip6.t4 3.3065
R17677 rstring_mux_0.vtrip6.n4 rstring_mux_0.vtrip6.t3 3.3065
R17678 rstring_mux_0.vtrip6.n1 rstring_mux_0.vtrip6.t8 3.3065
R17679 rstring_mux_0.vtrip6.n1 rstring_mux_0.vtrip6.t7 3.3065
R17680 rstring_mux_0.vtrip6 rstring_mux_0.vtrip6.t0 0.769662
R17681 rstring_mux_0.vtrip6 rstring_mux_0.vtrip6.n7 0.0563195
R17682 ibias_gen_0.ve.t1 ibias_gen_0.ve.n0 31121.7
R17683 ibias_gen_0.ve.n1 ibias_gen_0.ve.t1 146.25
R17684 ibias_gen_0.ve.n5 ibias_gen_0.ve.n4 62.2607
R17685 ibias_gen_0.ve.n4 ibias_gen_0.ve.n3 21.4545
R17686 ibias_gen_0.ve.n4 ibias_gen_0.ve.n2 20.7025
R17687 ibias_gen_0.ve.n5 ibias_gen_0.ve.n1 8.57525
R17688 sky130_fd_pr__rf_pnp_05v5_W0p68L0p68_0.Emitter ibias_gen_0.ve.n5 6.71196
R17689 ibias_gen_0.ve.n3 ibias_gen_0.ve.t4 3.3065
R17690 ibias_gen_0.ve.n3 ibias_gen_0.ve.t0 3.3065
R17691 ibias_gen_0.ve.n2 ibias_gen_0.ve.t2 3.3065
R17692 ibias_gen_0.ve.n2 ibias_gen_0.ve.t3 3.3065
R17693 sky130_fd_pr__rf_pnp_05v5_W0p68L0p68_0.Emitter ibias_gen_0.ve.n1 1.86379
R17694 rstring_mux_0.vtrip0.n5 rstring_mux_0.vtrip0.n3 50.7022
R17695 rstring_mux_0.vtrip0.n2 rstring_mux_0.vtrip0.n0 50.7022
R17696 rstring_mux_0.vtrip0.n7 rstring_mux_0.vtrip0.n6 25.1771
R17697 rstring_mux_0.vtrip0.n5 rstring_mux_0.vtrip0.n4 13.8791
R17698 rstring_mux_0.vtrip0.n2 rstring_mux_0.vtrip0.n1 13.8791
R17699 rstring_mux_0.vtrip0.n6 rstring_mux_0.vtrip0.n5 13.7519
R17700 rstring_mux_0.vtrip0.n7 rstring_mux_0.vtrip0.t3 10.6303
R17701 rstring_mux_0.vtrip0.n3 rstring_mux_0.vtrip0.t7 5.5395
R17702 rstring_mux_0.vtrip0.n3 rstring_mux_0.vtrip0.t6 5.5395
R17703 rstring_mux_0.vtrip0.n0 rstring_mux_0.vtrip0.t0 5.5395
R17704 rstring_mux_0.vtrip0.n0 rstring_mux_0.vtrip0.t1 5.5395
R17705 rstring_mux_0.vtrip0.n6 rstring_mux_0.vtrip0.n2 3.60196
R17706 rstring_mux_0.vtrip0.n4 rstring_mux_0.vtrip0.t8 3.3065
R17707 rstring_mux_0.vtrip0.n4 rstring_mux_0.vtrip0.t9 3.3065
R17708 rstring_mux_0.vtrip0.n1 rstring_mux_0.vtrip0.t5 3.3065
R17709 rstring_mux_0.vtrip0.n1 rstring_mux_0.vtrip0.t4 3.3065
R17710 rstring_mux_0.vtrip0 rstring_mux_0.vtrip0.t2 0.769662
R17711 rstring_mux_0.vtrip0 rstring_mux_0.vtrip0.n7 0.0563195
R17712 isrc_sel.n0 isrc_sel.t1 186.374
R17713 isrc_sel.n0 isrc_sel.t0 170.308
R17714 isrc_sel isrc_sel.n1 154.56
R17715 isrc_sel.n2 isrc_sel.n1 153.462
R17716 isrc_sel.n1 isrc_sel.n0 101.513
R17717 isrc_sel.n3 isrc_sel 11.8005
R17718 isrc_sel.n3 isrc_sel.n2 4.96991
R17719 isrc_sel.n2 isrc_sel 3.46403
R17720 isrc_sel isrc_sel.n3 2.71109
R17721 force_pdnb.n0 force_pdnb.t1 186.374
R17722 force_pdnb.n0 force_pdnb.t0 170.308
R17723 force_pdnb force_pdnb.n1 154.56
R17724 force_pdnb.n2 force_pdnb.n1 153.462
R17725 force_pdnb.n1 force_pdnb.n0 101.513
R17726 force_pdnb.n3 force_pdnb 11.8005
R17727 force_pdnb.n3 force_pdnb.n2 4.96991
R17728 force_pdnb.n2 force_pdnb 3.46403
R17729 force_pdnb force_pdnb.n3 2.71109
R17730 otrip_decoded[7].n0 otrip_decoded[7].t1 186.374
R17731 otrip_decoded[7].n0 otrip_decoded[7].t0 170.308
R17732 otrip_decoded[7] otrip_decoded[7].n1 154.56
R17733 otrip_decoded[7].n2 otrip_decoded[7].n1 153.462
R17734 otrip_decoded[7].n1 otrip_decoded[7].n0 101.513
R17735 otrip_decoded[7].n3 otrip_decoded[7] 11.8005
R17736 otrip_decoded[7].n3 otrip_decoded[7].n2 4.96991
R17737 otrip_decoded[7].n2 otrip_decoded[7] 3.46403
R17738 otrip_decoded[7] otrip_decoded[7].n3 2.71109
R17739 otrip_decoded[5].n0 otrip_decoded[5].t1 186.374
R17740 otrip_decoded[5].n0 otrip_decoded[5].t0 170.308
R17741 otrip_decoded[5] otrip_decoded[5].n1 154.56
R17742 otrip_decoded[5].n2 otrip_decoded[5].n1 153.462
R17743 otrip_decoded[5].n1 otrip_decoded[5].n0 101.513
R17744 otrip_decoded[5].n3 otrip_decoded[5] 11.8005
R17745 otrip_decoded[5].n3 otrip_decoded[5].n2 4.96991
R17746 otrip_decoded[5].n2 otrip_decoded[5] 3.46403
R17747 otrip_decoded[5] otrip_decoded[5].n3 2.71109
R17748 otrip_decoded[3].n0 otrip_decoded[3].t1 186.374
R17749 otrip_decoded[3].n0 otrip_decoded[3].t0 170.308
R17750 otrip_decoded[3] otrip_decoded[3].n1 154.56
R17751 otrip_decoded[3].n2 otrip_decoded[3].n1 153.462
R17752 otrip_decoded[3].n1 otrip_decoded[3].n0 101.513
R17753 otrip_decoded[3].n3 otrip_decoded[3] 11.8005
R17754 otrip_decoded[3].n3 otrip_decoded[3].n2 4.96991
R17755 otrip_decoded[3].n2 otrip_decoded[3] 3.46403
R17756 otrip_decoded[3] otrip_decoded[3].n3 2.71109
R17757 otrip_decoded[1].n0 otrip_decoded[1].t1 186.374
R17758 otrip_decoded[1].n0 otrip_decoded[1].t0 170.308
R17759 otrip_decoded[1] otrip_decoded[1].n1 154.56
R17760 otrip_decoded[1].n2 otrip_decoded[1].n1 153.462
R17761 otrip_decoded[1].n1 otrip_decoded[1].n0 101.513
R17762 otrip_decoded[1].n3 otrip_decoded[1] 11.8005
R17763 otrip_decoded[1].n3 otrip_decoded[1].n2 4.96991
R17764 otrip_decoded[1].n2 otrip_decoded[1] 3.46403
R17765 otrip_decoded[1] otrip_decoded[1].n3 2.71109
C0 schmitt_trigger_0.m dvdd 2.68752f
C1 rc_osc_0.m osc_ck 1.09227f
C2 comparator_0.vnn avdd 37.3292f
C3 rc_osc_0.m dvdd 2.38628f
C4 vl dvdd 1.78644f
C5 sky130_fd_sc_hd__inv_4_1.Y porb 1.48088f
C6 rstring_mux_0.otrip_decoded_avdd[3] avss 1.341f
C7 comparator_1.vt avss 29.094501f
C8 rstring_mux_0.vtrip6 vin 2.08469f
C9 comparator_0.n1 avss 3.03066f
C10 rstring_mux_0.ena ibias_gen_0.ena_b 1.24167f
C11 dvdd osc_ck 1.35201f
C12 comparator_1.n1 dcomp3v3 1.70353f
C13 vl avdd 2.83098f
C14 rstring_mux_0.otrip_decoded_avdd[6] avdd 1.62903f
C15 rstring_mux_0.ena_b avdd 6.38079f
C16 rstring_mux_0.vtrip_decoded_avdd[7] rstring_mux_0.vtrip_decoded_avdd[6] 3.06282f
C17 ibias_gen_0.isrc_sel avss 3.29158f
C18 avdd vbg_1v2 6.81536f
C19 avdd dvdd 46.8833f
C20 ibias_gen_0.vp1 avdd 6.59272f
C21 comparator_1.vm avss 10.3557f
C22 dvdd dcomp 1.54533f
C23 ibias_gen_0.ibias0 vbg_1v2 2.28759f
C24 comparator_1.vpp avss 1.79171f
C25 rstring_mux_0.otrip_decoded_avdd[0] avss 1.64125f
C26 rstring_mux_0.ena ibias_gen_0.isrc_sel_b 1.98919f
C27 rstring_mux_0.otrip_decoded_avdd[4] avdd 1.52975f
C28 rc_osc_0.vr dvdd 1.51499f
C29 rstring_mux_0.vtrip_decoded_avdd[5] rstring_mux_0.vtrip_decoded_avdd[6] 1.33995f
C30 ibias_gen_0.ibias0 avdd 2.5318f
C31 comparator_0.vt comparator_0.vnn 4.29222f
C32 comparator_0.vn comparator_0.n0 1.99139f
C33 comparator_0.n0 avdd 1.07016f
C34 comparator_1.n1 avss 3.02944f
C35 rstring_mux_0.otrip_decoded_avdd[2] avdd 1.52848f
C36 avss vin 13.112f
C37 rstring_mux_0.vtrip_decoded_avdd[5] rstring_mux_0.vtrip_decoded_avdd[4] 2.29102f
C38 sky130_fd_sc_hvl__inv_1_0.A avss 2.32435f
C39 rstring_mux_0.vtrip_decoded_avdd[6] avss 1.44633f
C40 ibias_gen_0.ena_b avdd 2.96986f
C41 comparator_0.vt vbg_1v2 24.362598f
C42 rstring_mux_0.ena rstring_mux_0.vtrip_decoded_avdd[7] 1.91505f
C43 rstring_mux_0.ena comparator_0.ibias 2.32983f
C44 sky130_fd_sc_hd__inv_4_0.Y pwup_filt 1.46398f
C45 comparator_0.vt avdd 0.142093p
C46 rstring_mux_0.vtrip_decoded_avdd[3] rstring_mux_0.vtrip_decoded_avdd[4] 1.04751f
C47 rstring_mux_0.vtrip_decoded_avdd[4] avss 1.50015f
C48 ibias_gen_0.isrc_sel_b avdd 3.36468f
C49 comparator_1.vnn vbg_1v2 3.55942f
C50 rstring_mux_0.otrip_decoded_avdd[1] avdd 1.73972f
C51 dcomp3v3uv dvdd 1.09406f
C52 rstring_mux_0.vtrip_decoded_avdd[3] rstring_mux_0.vtrip_decoded_avdd[2] 1.78143f
C53 dcomp3v3 vl 10.054f
C54 rstring_mux_0.vtrip_decoded_avdd[2] avss 1.41004f
C55 comparator_1.vnn avdd 37.3119f
C56 comparator_1.vnn ibias_gen_0.ibias0 1.84751f
C57 sky130_fd_sc_hd__inv_4_4.Y dvdd 1.32154f
C58 dcomp3v3uv avdd 5.82321f
C59 rstring_mux_0.ena avss 18.5982f
C60 dcomp3v3 dvdd 1.10728f
C61 sky130_fd_sc_hvl__inv_16_0.A porb_h 2.44559f
C62 ibias_gen_0.ena_b ibias_gen_0.isrc_sel_b 3.0701f
C63 comparator_1.vt comparator_1.vpp 2.58192f
C64 rstring_mux_0.vtrip_decoded_avdd[7] avdd 1.81913f
C65 rstring_mux_0.ena schmitt_trigger_0.in 1.1842f
C66 rstring_mux_0.vtrip_decoded_avdd[0] avss 1.37856f
C67 avss porb_h 1.14661f
C68 dcomp3v3 avdd 6.72641f
C69 sky130_fd_sc_hvl__inv_4_0.A avdd 1.01652f
C70 comparator_0.ibias avdd 7.48432f
C71 comparator_0.vnn avss 3.71294f
C72 dvdd porb 1.54357f
C73 comparator_1.vn comparator_1.n0 1.97873f
C74 sky130_fd_sc_hd__inv_4_3.Y dvdd 1.31104f
C75 comparator_0.vpp comparator_0.vnn 8.55337f
C76 rstring_mux_0.vtrip_decoded_avdd[5] avdd 2.25645f
C77 rstring_mux_0.vtrip_decoded_avdd[1] rstring_mux_0.vtrip_decoded_avdd[0] 1.27051f
C78 comparator_1.vt vin 24.7245f
C79 vl avss 1.65817f
C80 rstring_mux_0.otrip_decoded_avdd[6] avss 1.36421f
C81 rstring_mux_0.ena_b avss 1.61845f
C82 sky130_fd_sc_hvl__lsbufhv2lv_1_1.X dvdd 1.00946f
C83 sky130_fd_sc_hd__inv_4_3.Y dcomp 1.48254f
C84 avss vbg_1v2 12.430799f
C85 sky130_fd_sc_hvl__lsbufhv2lv_1_1.X avdd 3.01571f
C86 avss dvdd 2.39761f
C87 comparator_0.vn avss 8.98359f
C88 sky130_fd_sc_hvl__inv_16_0.A avdd 3.72269f
C89 ibias_gen_0.vp1 avss 2.02475f
C90 dvdd por 1.54891f
C91 rstring_mux_0.vtrip_decoded_avdd[3] avdd 1.87754f
C92 comparator_0.vpp vbg_1v2 2.95415f
C93 avdd avss 2.43719p
C94 schmitt_trigger_0.in dvdd 2.4917f
C95 rstring_mux_0.otrip_decoded_avdd[4] avss 1.34995f
C96 rstring_mux_0.vtrip0 avss 2.36542f
C97 comparator_1.vpp vin 3.00612f
C98 ibias_gen_0.ibias0 avss 1.14374f
C99 schmitt_trigger_0.in avdd 4.44429f
C100 comparator_0.vpp avdd 37.286697f
C101 comparator_0.n0 avss 4.20459f
C102 rstring_mux_0.vtrip_decoded_avdd[1] avdd 1.96911f
C103 rstring_mux_0.otrip_decoded_avdd[7] rstring_mux_0.otrip_decoded_avdd[6] 1.12965f
C104 rstring_mux_0.otrip_decoded_avdd[2] avss 1.41238f
C105 rstring_mux_0.ena_b rstring_mux_0.vtop 2.52783f
C106 comparator_0.ena_b comparator_0.vn 1.12681f
C107 ibias_gen_0.ena_b avss 2.71238f
C108 rstring_mux_0.vtrip2 avss 2.19733f
C109 sky130_fd_sc_hd__inv_4_0.Y dvdd 1.35239f
C110 comparator_0.ena_b avdd 1.01938f
C111 comparator_1.vn avss 8.76998f
C112 rstring_mux_0.otrip_decoded_avdd[7] avdd 1.82047f
C113 comparator_0.vt avss 29.296902f
C114 rstring_mux_0.ena ibias_gen_0.isrc_sel 1.49913f
C115 rstring_mux_0.vtop avdd 10.640901f
C116 comparator_0.vt comparator_0.vpp 2.58192f
C117 ibias_gen_0.isrc_sel_b avss 2.66768f
C118 comparator_0.vn comparator_0.vm 4.66142f
C119 rstring_mux_0.vtrip4 avss 2.05606f
C120 rstring_mux_0.otrip_decoded_avdd[1] avss 1.63066f
C121 rstring_mux_0.otrip_decoded_avdd[5] avdd 1.82417f
C122 rstring_mux_0.otrip_decoded_avdd[5] rstring_mux_0.otrip_decoded_avdd[4] 1.15427f
C123 dvdd por_unbuf 1.64561f
C124 comparator_1.n0 avss 3.94624f
C125 dcomp3v3uv sky130_fd_sc_hvl__lsbufhv2lv_1_1.X 2.56892f
C126 comparator_1.vnn avss 3.08013f
C127 dcomp3v3uv avss 7.27403f
C128 comparator_1.vt vbg_1v2 25.626f
C129 comparator_0.vm comparator_0.n0 2.61558f
C130 rstring_mux_0.otrip_decoded_avdd[3] avdd 1.72135f
C131 rstring_mux_0.ena vin 2.34886f
C132 rstring_mux_0.vtrip6 avss 2.27146f
C133 comparator_1.ena_b comparator_1.vn 1.12092f
C134 comparator_1.vt avdd 0.141755p
C135 rstring_mux_0.vtrip_decoded_avdd[7] avss 1.38048f
C136 comparator_0.n1 avdd 2.68846f
C137 dcomp3v3 avss 3.78844f
C138 sky130_fd_sc_hd__inv_4_4.Y por 1.48254f
C139 comparator_0.ibias avss 5.42518f
C140 sky130_fd_sc_hd__inv_4_1.Y dvdd 1.26215f
C141 ibias_gen_0.isrc_sel avdd 10.48f
C142 comparator_1.vpp vbg_1v2 2.54472f
C143 dvdd pwup_filt 1.55425f
C144 rstring_mux_0.otrip_decoded_avdd[3] rstring_mux_0.otrip_decoded_avdd[2] 1.42613f
C145 rstring_mux_0.vtrip_decoded_avdd[5] avss 1.50537f
C146 comparator_1.vpp avdd 37.1895f
C147 rstring_mux_0.otrip_decoded_avdd[0] avdd 1.34894f
C148 comparator_1.vpp ibias_gen_0.ibias0 1.31426f
C149 sky130_fd_sc_hvl__inv_16_0.A avss 4.17343f
C150 vbg_1v2 vin 7.66271f
C151 ibias_gen_0.ena_b ibias_gen_0.isrc_sel 1.07804f
C152 rstring_mux_0.vtrip_decoded_avdd[3] avss 1.48249f
C153 rc_osc_0.in rc_osc_0.m 1.10731f
C154 comparator_1.n1 avdd 2.69603f
C155 avdd vin 7.70762f
C156 rstring_mux_0.vtrip_decoded_avdd[6] avdd 1.9364f
C157 rc_osc_0.in osc_ck 1.05774f
C158 rstring_mux_0.vtrip0 vin 2.24047f
C159 schmitt_trigger_0.in avss 8.85536f
C160 comparator_0.vpp avss 2.41468f
C161 comparator_1.vn comparator_1.vm 4.6608f
C162 rc_osc_0.in dvdd 5.2937f
C163 rstring_mux_0.vtrip_decoded_avdd[1] avss 1.39274f
C164 ibias_gen_0.isrc_sel ibias_gen_0.isrc_sel_b 1.79811f
C165 comparator_1.vt comparator_1.vnn 4.17609f
C166 rstring_mux_0.vtrip_decoded_avdd[4] avdd 1.61396f
C167 dcomp3v3uv comparator_0.n1 1.71428f
C168 rstring_mux_0.vtrip2 vin 2.09579f
C169 comparator_0.ena_b avss 2.38822f
C170 comparator_1.vm comparator_1.n0 2.59034f
C171 rstring_mux_0.otrip_decoded_avdd[7] avss 1.37218f
C172 rstring_mux_0.otrip_decoded_avdd[1] rstring_mux_0.otrip_decoded_avdd[0] 3.24722f
C173 comparator_1.vt dcomp3v3 2.36366f
C174 rstring_mux_0.vtop avss 3.67651f
C175 comparator_1.ena_b avss 1.77799f
C176 rstring_mux_0.vtrip_decoded_avdd[2] avdd 1.66091f
C177 comparator_1.vpp comparator_1.vnn 8.65712f
C178 dcomp3v3 ibias_gen_0.isrc_sel 10.963901f
C179 rstring_mux_0.ena avdd 16.1312f
C180 rstring_mux_0.vtrip4 vin 2.26482f
C181 rstring_mux_0.otrip_decoded_avdd[5] avss 1.34873f
C182 comparator_0.vm avss 10.3984f
C183 rstring_mux_0.ena ibias_gen_0.ibias0 1.70445f
C184 rstring_mux_0.vtrip_decoded_avdd[0] avdd 1.59456f
C185 avdd porb_h 3.53805f
C186 rstring_mux_0.otrip_decoded_avdd[3] sky130_fd_sc_hvl__lsbufhv2lv_1_1.X 1.37931f
C187 osc_ck dvss 3.25723f
C188 osc_ena dvss 2.21578f
C189 porb dvss 1.2588f
C190 pwup_filt dvss 1.31705f
C191 dcomp dvss 1.25321f
C192 por dvss 1.2619f
C193 por_unbuf dvss 5.05078f
C194 vin dvss 24.4908f
C195 vbg_1v2 dvss 47.514263f
C196 porb_h dvss -3.025187f
C197 dvdd dvss 0.988996p
C198 avss dvss 0.214264p
C199 avdd dvss 3.614321p
C200 a_12321_n25357# dvss 1.27808f
C201 a_n10279_n24979# dvss 1.13069f
C202 a_n10279_n24223# dvss 1.13821f
C203 a_n10279_n23467# dvss 1.31493f
C204 a_n10279_n22711# dvss 1.20647f
C205 a_12321_n22333# dvss 1.27347f
C206 rc_osc_0.vr dvss 4.10332f
C207 rc_osc_0.m dvss 3.35349f
C208 rc_osc_0.in dvss 0.439703p
C209 rc_osc_0.ena_b dvss 1.39535f
C210 a_n8941_n11914# dvss 1.04349f
C211 comparator_0.n1 dvss 1.57269f
C212 comparator_0.vm dvss 4.68965f
C213 comparator_0.vn dvss 5.29407f
C214 comparator_0.vnn dvss 44.4245f
C215 comparator_0.vpp dvss 38.2361f
C216 rstring_mux_0.vtrip6 dvss 6.108224f
C217 rstring_mux_0.vtrip4 dvss 6.24356f
C218 rstring_mux_0.vtrip2 dvss 6.0667f
C219 rstring_mux_0.vtrip0 dvss 6.512494f
C220 rstring_mux_0.vtop dvss 16.18401f
C221 rstring_mux_0.ena_b dvss 2.14258f
C222 sky130_fd_sc_hvl__lsbufhv2lv_1_1.X dvss 3.25948f
C223 a_9145_n3946# dvss 1.70782f
C224 a_7033_n3946# dvss 1.72434f
C225 a_4921_n3946# dvss 1.72666f
C226 a_2809_n3946# dvss 1.72672f
C227 a_697_n3946# dvss 1.72474f
C228 a_n1415_n3946# dvss 1.71031f
C229 a_n3527_n3946# dvss 1.70837f
C230 a_n5639_n3946# dvss 1.70837f
C231 a_n7751_n3946# dvss 1.70982f
C232 a_10873_n3956# dvss 1.0124f
C233 dcomp3v3uv dvss 7.64891f
C234 a_10514_n2760# dvss 1.27441f
C235 rstring_mux_0.vtrip_decoded_avdd[6] dvss 1.45969f
C236 rstring_mux_0.vtrip_decoded_avdd[4] dvss 1.44257f
C237 rstring_mux_0.vtrip_decoded_avdd[2] dvss 1.71779f
C238 rstring_mux_0.vtrip_decoded_avdd[0] dvss 1.50396f
C239 rstring_mux_0.otrip_decoded_avdd[6] dvss 1.25109f
C240 rstring_mux_0.otrip_decoded_avdd[4] dvss 1.06381f
C241 rstring_mux_0.otrip_decoded_avdd[2] dvss 1.43078f
C242 rstring_mux_0.otrip_decoded_avdd[0] dvss 1.07955f
C243 a_8877_n2876# dvss 1.52129f
C244 a_8777_n2964# dvss 1.97869f
C245 a_6765_n2876# dvss 1.52795f
C246 a_6665_n2964# dvss 2.199f
C247 a_4653_n2876# dvss 1.52792f
C248 a_4553_n2964# dvss 2.19988f
C249 a_2541_n2876# dvss 1.52796f
C250 a_2441_n2964# dvss 2.19989f
C251 a_429_n2876# dvss 1.52795f
C252 a_329_n2964# dvss 2.19989f
C253 a_n1683_n2876# dvss 1.52227f
C254 a_n1783_n2964# dvss 1.97975f
C255 a_n3795_n2876# dvss 1.52226f
C256 a_n3895_n2964# dvss 1.97975f
C257 a_n5907_n2876# dvss 1.52226f
C258 a_n6007_n2964# dvss 1.97975f
C259 a_n8019_n2876# dvss 1.53095f
C260 a_n8119_n2964# dvss 2.03637f
C261 a_9145_n2212# dvss 1.69093f
C262 a_7033_n2212# dvss 1.7079f
C263 a_4921_n2212# dvss 1.70983f
C264 a_2809_n2212# dvss 1.70983f
C265 a_697_n2212# dvss 1.70983f
C266 a_n1415_n2212# dvss 1.69341f
C267 a_n3527_n2212# dvss 1.69148f
C268 a_n5639_n2212# dvss 1.69215f
C269 a_n7751_n2212# dvss 1.69294f
C270 a_10874_n2222# dvss 1.00525f
C271 a_10515_n1026# dvss 1.27471f
C272 rstring_mux_0.vtrip_decoded_avdd[7] dvss 2.19603f
C273 rstring_mux_0.vtrip_decoded_avdd[5] dvss 2.01311f
C274 rstring_mux_0.vtrip_decoded_avdd[3] dvss 2.08084f
C275 rstring_mux_0.vtrip_decoded_avdd[1] dvss 2.16902f
C276 rstring_mux_0.otrip_decoded_avdd[7] dvss 1.93903f
C277 rstring_mux_0.otrip_decoded_avdd[5] dvss 1.92238f
C278 rstring_mux_0.otrip_decoded_avdd[3] dvss 1.59657f
C279 rstring_mux_0.otrip_decoded_avdd[1] dvss 1.7578f
C280 a_8877_n1142# dvss 1.52856f
C281 a_8777_n1230# dvss 1.97228f
C282 a_6765_n1142# dvss 1.53263f
C283 a_6665_n1230# dvss 2.18683f
C284 a_4653_n1142# dvss 1.53264f
C285 a_4553_n1230# dvss 2.18683f
C286 a_2541_n1142# dvss 1.53264f
C287 a_2441_n1230# dvss 2.18683f
C288 a_429_n1142# dvss 1.53264f
C289 a_329_n1230# dvss 2.18683f
C290 a_n1683_n1142# dvss 1.52954f
C291 a_n1783_n1230# dvss 1.96643f
C292 a_n3795_n1142# dvss 1.52683f
C293 a_n3895_n1230# dvss 1.96734f
C294 a_n5907_n1142# dvss 1.53695f
C295 a_n6007_n1230# dvss 1.97338f
C296 a_n8019_n1142# dvss 1.53771f
C297 a_n8119_n1230# dvss 2.02842f
C298 sky130_fd_sc_hd__inv_4_1.Y dvss 2.05067f
C299 sky130_fd_sc_hd__inv_4_0.Y dvss 1.95044f
C300 schmitt_trigger_0.m dvss 2.262503f
C301 sky130_fd_sc_hd__inv_4_3.Y dvss 1.97752f
C302 sky130_fd_sc_hd__inv_4_4.Y dvss 1.98989f
C303 ibias_gen_0.isrc_sel_b dvss 1.33811f
C304 ibias_gen_0.isrc_sel dvss 5.25818f
C305 ibias_gen_0.ena_b dvss 1.24326f
C306 a_n3510_6789# dvss 1.69444f
C307 a_n3778_7859# dvss 1.54444f
C308 a_n3878_7771# dvss 2.03411f
C309 comparator_0.ibias dvss 2.76603f
C310 ibias_gen_0.vp1 dvss 4.798203f
C311 schmitt_trigger_0.in dvss 0.409533p
C312 vl dvss 7.07645f
C313 dcomp3v3 dvss 1.23522f
C314 comparator_1.n1 dvss 1.34067f
C315 comparator_1.vm dvss 4.47408f
C316 comparator_1.vn dvss 4.961259f
C317 rstring_mux_0.ena dvss 8.83325f
C318 sky130_fd_sc_hvl__inv_16_0.A dvss 1.75005f
C319 sky130_fd_sc_hvl__inv_1_0.A dvss 3.80079f
C320 comparator_1.vnn dvss 30.1825f
C321 comparator_1.vpp dvss 29.323698f
C322 comparator_0.vt dvss 11.7607f
C323 comparator_1.vt dvss 4.36096f
C324 rstring_mux_0.vtrip0.n5 dvss 1.22742f
C325 rstring_mux_0.vtrip0.n6 dvss 2.02058f
C326 rstring_mux_0.vtrip0.n7 dvss 2.41105f
C327 ibias_gen_0.ve.n0 dvss -12.6698f
C328 ibias_gen_0.ve.t1 dvss 12.8312f
C329 ibias_gen_0.ve.n4 dvss 10.320901f
C330 ibias_gen_0.ve.n5 dvss 11.6084f
C331 rstring_mux_0.vtrip6.n5 dvss 1.249f
C332 rstring_mux_0.vtrip6.n6 dvss 1.9489f
C333 rstring_mux_0.vtrip6.n7 dvss 2.19091f
C334 rstring_mux_0.vtrip1.n5 dvss 1.52407f
C335 rstring_mux_0.vtrip1.n6 dvss 1.30427f
C336 rstring_mux_0.vtrip1.n7 dvss 3.51872f
C337 rstring_mux_0.vtrip5.n2 dvss 1.20735f
C338 rstring_mux_0.vtrip5.n7 dvss 2.7123f
C339 ibias_gen_0.vstart.n0 dvss 1.41043f
C340 rstring_mux_0.vtrip3.n5 dvss 1.08769f
C341 rstring_mux_0.vtrip3.n7 dvss 2.47396f
C342 ibias_gen_0.vn1.t0 dvss 2.11164f
C343 ibias_gen_0.vn1.t15 dvss 2.11164f
C344 ibias_gen_0.vn1.t10 dvss 2.19722f
C345 ibias_gen_0.vn1.n2 dvss 1.40052f
C346 ibias_gen_0.vn1.t17 dvss 2.11164f
C347 ibias_gen_0.vn1.t14 dvss 2.19722f
C348 ibias_gen_0.vn1.n3 dvss 1.3685f
C349 ibias_gen_0.vn1.t11 dvss 2.11164f
C350 ibias_gen_0.vn1.t12 dvss 2.19722f
C351 ibias_gen_0.vn1.n5 dvss 1.40052f
C352 ibias_gen_0.vn1.t13 dvss 2.11164f
C353 ibias_gen_0.vn1.t16 dvss 2.19722f
C354 ibias_gen_0.vn1.n6 dvss 1.3685f
C355 ibias_gen_0.vn1.t2 dvss 2.15704f
C356 ibias_gen_0.vp1.n0 dvss 2.2551f
C357 ibias_gen_0.vp1.t11 dvss 2.72493f
C358 ibias_gen_0.vp1.n3 dvss 2.14115f
C359 ibias_gen_0.vp1.t13 dvss 2.72114f
C360 rstring_mux_0.vtrip2.n5 dvss 1.50485f
C361 rstring_mux_0.vtrip2.n6 dvss 2.43692f
C362 rstring_mux_0.vtrip2.n7 dvss 2.0739f
C363 rstring_mux_0.vtrip7.n5 dvss 1.19247f
C364 rstring_mux_0.vtrip7.n7 dvss 2.50533f
C365 ibias_gen_0.vp.t11 dvss 1.71268f
C366 ibias_gen_0.vp.n4 dvss 1.29098f
C367 ibias_gen_0.vp.t8 dvss 1.65245f
C368 ibias_gen_0.vp.n5 dvss 1.29098f
C369 ibias_gen_0.vp.t7 dvss 1.65245f
C370 ibias_gen_0.vp.n6 dvss 1.29098f
C371 ibias_gen_0.vp.t9 dvss 1.68256f
C372 ibias_gen_0.vp.t10 dvss 2.31092f
C373 ibias_gen_0.vp.t12 dvss 2.34104f
C374 ibias_gen_0.vp.n9 dvss 1.1851f
C375 ibias_gen_0.vr.n2 dvss 1.54735f
C376 ibias_gen_0.vp0.t6 dvss 1.72871f
C377 ibias_gen_0.vp0.n6 dvss 1.47471f
C378 ibias_gen_0.vp0.t13 dvss 1.76142f
C379 ibias_gen_0.vp0.t12 dvss 1.69947f
C380 ibias_gen_0.vp0.n8 dvss 1.47471f
C381 ibias_gen_0.vp0.t8 dvss 1.69947f
C382 ibias_gen_0.vp0.n13 dvss 1.07524f
C383 ibias_gen_0.Mt4 dvss 1.25878f
C384 ibias_gen_0.vn0.n1 dvss 1.39652f
C385 ibias_gen_0.vn0.t19 dvss 2.24075f
C386 ibias_gen_0.vn0.t5 dvss 2.19836f
C387 ibias_gen_0.vn0.t7 dvss 2.16084f
C388 ibias_gen_0.vn0.n8 dvss 1.01955f
C389 ibias_gen_0.vn0.n9 dvss 1.87632f
C390 ibias_gen_0.vn0.t20 dvss 2.16084f
C391 ibias_gen_0.vn0.n10 dvss 1.71213f
C392 schmitt_trigger_0.in.t7 dvss 2.42609f
C393 schmitt_trigger_0.in.t14 dvss 1.30645f
C394 schmitt_trigger_0.in.n5 dvss 1.47048f
C395 schmitt_trigger_0.in.t12 dvss 1.30645f
C396 schmitt_trigger_0.in.n6 dvss 1.29757f
C397 schmitt_trigger_0.in.t6 dvss 1.30645f
C398 schmitt_trigger_0.in.n7 dvss 1.29757f
C399 schmitt_trigger_0.in.t13 dvss 1.30645f
C400 schmitt_trigger_0.in.n8 dvss 1.29757f
C401 schmitt_trigger_0.in.t11 dvss 1.30645f
C402 schmitt_trigger_0.in.n9 dvss 1.38463f
C403 vbg_1v2.t0 dvss 1.85934f
C404 vbg_1v2.t5 dvss 1.77938f
C405 vbg_1v2.n0 dvss 1.48175f
C406 vbg_1v2.t18 dvss 1.77938f
C407 vbg_1v2.t38 dvss 1.77938f
C408 vbg_1v2.t17 dvss 1.77938f
C409 vbg_1v2.t37 dvss 1.77938f
C410 vbg_1v2.t2 dvss 1.77938f
C411 vbg_1v2.t12 dvss 1.77938f
C412 vbg_1v2.t15 dvss 1.87524f
C413 vbg_1v2.t26 dvss 1.79416f
C414 vbg_1v2.n7 dvss 1.51506f
C415 vbg_1v2.t36 dvss 1.79416f
C416 vbg_1v2.t10 dvss 1.79416f
C417 vbg_1v2.t35 dvss 1.79416f
C418 vbg_1v2.t9 dvss 1.79416f
C419 vbg_1v2.t21 dvss 1.79416f
C420 vbg_1v2.t31 dvss 1.79416f
C421 vbg_1v2.n14 dvss 1.48593f
C422 vbg_1v2.n15 dvss 1.03806f
C423 vbg_1v2.t20 dvss 1.66117f
C424 vbg_1v2.t33 dvss 1.52003f
C425 vbg_1v2.n16 dvss 1.03384f
C426 vbg_1v2.t8 dvss 1.66117f
C427 vbg_1v2.n19 dvss 1.03384f
C428 vbg_1v2.t27 dvss 1.52003f
C429 vbg_1v2.n20 dvss 1.03384f
C430 vbg_1v2.t34 dvss 1.66117f
C431 vbg_1v2.n23 dvss 1.03384f
C432 vbg_1v2.t6 dvss 1.52003f
C433 vbg_1v2.n24 dvss 1.03384f
C434 vbg_1v2.t24 dvss 1.66117f
C435 vbg_1v2.n27 dvss 1.03384f
C436 vbg_1v2.t39 dvss 1.52003f
C437 vbg_1v2.n28 dvss 1.03384f
C438 vbg_1v2.t3 dvss 1.66117f
C439 vbg_1v2.n31 dvss 1.03384f
C440 vbg_1v2.t19 dvss 1.52003f
C441 vbg_1v2.n32 dvss 1.03384f
C442 vbg_1v2.t25 dvss 1.66117f
C443 vbg_1v2.n35 dvss 1.03384f
C444 vbg_1v2.t40 dvss 1.52003f
C445 vbg_1v2.n36 dvss 1.03384f
C446 vbg_1v2.t14 dvss 1.66117f
C447 vbg_1v2.n39 dvss 1.03384f
C448 vbg_1v2.t30 dvss 1.52003f
C449 vbg_1v2.n40 dvss 1.03384f
C450 vbg_1v2.t11 dvss 1.66117f
C451 vbg_1v2.n43 dvss 1.03384f
C452 vbg_1v2.t28 dvss 1.52003f
C453 vbg_1v2.n44 dvss 1.03384f
C454 vbg_1v2.n45 dvss 1.29901f
C455 vbg_1v2.n46 dvss 1.64068f
C456 rstring_mux_0.vtop.n2 dvss 1.02937f
C457 rstring_mux_0.vtop.t17 dvss 2.67225f
C458 dvdd.n282 dvss 1.35829f
C459 dvdd.n284 dvss 1.37226f
C460 dvdd.n285 dvss 1.35801f
C461 dvdd.n286 dvss 1.37198f
C462 dvdd.n475 dvss 2.0428f
C463 dvdd.n477 dvss 1.1648f
C464 dvdd.n478 dvss 1.1648f
C465 dvdd.n479 dvss 4.44184f
C466 dvdd.n480 dvss 1.16863f
C467 dvdd.n481 dvss 4.50046f
C468 dvdd.n482 dvss 4.44184f
C469 dvdd.n483 dvss 4.50046f
C470 dvdd.n484 dvss 1.16863f
C471 dvdd.n486 dvss 2.5207f
C472 dvdd.n520 dvss 1.06744f
C473 dvdd.n525 dvss 2.07496f
C474 avdd.t163 dvss 1.7701f
C475 avdd.t6 dvss 1.23737f
C476 avdd.n7 dvss 1.51706f
C477 avdd.n22 dvss 1.0555f
C478 avdd.t10 dvss 1.95275f
C479 avdd.t159 dvss 1.30536f
C480 avdd.t438 dvss 1.95275f
C481 avdd.t151 dvss 1.30536f
C482 avdd.t14 dvss 1.95275f
C483 avdd.t492 dvss 1.30536f
C484 avdd.t147 dvss 1.95275f
C485 avdd.t149 dvss 1.30536f
C486 avdd.t442 dvss 1.95275f
C487 avdd.t422 dvss 1.30536f
C488 avdd.t107 dvss 1.95275f
C489 avdd.t99 dvss 1.30536f
C490 avdd.t207 dvss 1.95275f
C491 avdd.t103 dvss 1.30536f
C492 avdd.t101 dvss 1.95275f
C493 avdd.t123 dvss 1.30536f
C494 avdd.t42 dvss 1.37501f
C495 avdd.n111 dvss 1.209f
C496 avdd.t211 dvss 1.2819f
C497 avdd.n159 dvss 1.37272f
C498 avdd.n162 dvss 1.16441f
C499 avdd.n187 dvss 1.37272f
C500 avdd.n190 dvss 1.16441f
C501 avdd.n215 dvss 1.37272f
C502 avdd.n218 dvss 1.16441f
C503 avdd.n243 dvss 1.37272f
C504 avdd.n246 dvss 1.16441f
C505 avdd.n271 dvss 1.37272f
C506 avdd.n274 dvss 1.16441f
C507 avdd.n299 dvss 1.37272f
C508 avdd.n302 dvss 1.16441f
C509 avdd.n327 dvss 1.37272f
C510 avdd.n330 dvss 1.16441f
C511 avdd.n355 dvss 1.37272f
C512 avdd.n358 dvss 1.16441f
C513 avdd.n370 dvss 7.35223f
C514 avdd.t498 dvss 1.95275f
C515 avdd.t588 dvss 1.30536f
C516 avdd.t2 dvss 1.95275f
C517 avdd.t91 dvss 1.30536f
C518 avdd.t155 dvss 1.95275f
C519 avdd.t173 dvss 1.30536f
C520 avdd.t127 dvss 1.95275f
C521 avdd.t142 dvss 1.30536f
C522 avdd.t396 dvss 1.95275f
C523 avdd.t34 dvss 1.30536f
C524 avdd.t576 dvss 1.95275f
C525 avdd.t619 dvss 1.30536f
C526 avdd.t452 dvss 1.95275f
C527 avdd.t36 dvss 1.30536f
C528 avdd.t38 dvss 1.95275f
C529 avdd.t586 dvss 1.30536f
C530 avdd.t45 dvss 1.37471f
C531 avdd.n448 dvss 1.209f
C532 avdd.t131 dvss 1.2819f
C533 avdd.n496 dvss 1.37272f
C534 avdd.n499 dvss 1.16441f
C535 avdd.n524 dvss 1.37272f
C536 avdd.n527 dvss 1.16441f
C537 avdd.n552 dvss 1.37272f
C538 avdd.n555 dvss 1.16441f
C539 avdd.n580 dvss 1.37272f
C540 avdd.n583 dvss 1.16441f
C541 avdd.n608 dvss 1.37272f
C542 avdd.n611 dvss 1.16441f
C543 avdd.n636 dvss 1.37272f
C544 avdd.n639 dvss 1.16441f
C545 avdd.n664 dvss 1.37272f
C546 avdd.n667 dvss 1.16441f
C547 avdd.n692 dvss 1.37272f
C548 avdd.n695 dvss 1.16441f
C549 avdd.n707 dvss 4.01271f
C550 avdd.n708 dvss 5.91925f
C551 avdd.n709 dvss 5.175931f
C552 avdd.n723 dvss 1.07024f
C553 avdd.n725 dvss 1.0502f
C554 avdd.n727 dvss 2.0713f
C555 avdd.n728 dvss 2.0713f
C556 avdd.n730 dvss 1.05069f
C557 avdd.n967 dvss 1.01886f
C558 avdd.n984 dvss 2.45955f
C559 avdd.n985 dvss 9.45219f
C560 avdd.n987 dvss 2.68905f
C561 avdd.t220 dvss 2.83122f
C562 avdd.n988 dvss 1.37069f
C563 avdd.n992 dvss 1.32443f
C564 avdd.n993 dvss 1.40599f
C565 avdd.n994 dvss 2.23246f
C566 avdd.t221 dvss 47.8713f
C567 avdd.n996 dvss 2.67548f
C568 avdd.n997 dvss 2.46292f
C569 avdd.n998 dvss 1.52014f
C570 avdd.n999 dvss 1.44595f
C571 avdd.t167 dvss 1.31907f
C572 avdd.t141 dvss 1.82555f
C573 avdd.n1005 dvss 1.61596f
C574 avdd.t169 dvss 1.50199f
C575 avdd.t165 dvss 1.65232f
C576 avdd.n1007 dvss 1.42336f
C577 avdd.n1012 dvss 2.11868f
C578 avdd.n1013 dvss 1.52014f
C579 avdd.t186 dvss 45.4238f
C580 avdd.t177 dvss 60.565098f
C581 avdd.t179 dvss 45.4238f
C582 avdd.n1014 dvss 1.40599f
C583 avdd.n1018 dvss 1.90355f
C584 avdd.n1019 dvss 1.76059f
C585 avdd.n1046 dvss 2.54367f
C586 avdd.n1050 dvss 4.16674f
C587 avdd.n1051 dvss 4.1662f
C588 avdd.n1052 dvss 15.7194f
C589 avdd.n1053 dvss 1.01273f
C590 avdd.n1056 dvss 1.77866f
C591 avdd.n1058 dvss 1.51886f
C592 avdd.n1064 dvss 2.80462f
C593 avdd.n1065 dvss 3.09468f
C594 avdd.n1066 dvss 2.79818f
C595 avdd.t53 dvss 1.14721f
C596 avdd.n1071 dvss 1.51918f
C597 avdd.t418 dvss 1.14721f
C598 avdd.n1072 dvss 1.51918f
C599 avdd.n1097 dvss 3.57199f
C600 avdd.n1098 dvss 2.68905f
C601 avdd.t281 dvss 2.81462f
C602 avdd.t376 dvss 2.81531f
C603 avdd.t249 dvss 2.81531f
C604 avdd.n1104 dvss 1.38758f
C605 avdd.t385 dvss 2.81531f
C606 avdd.n1107 dvss 1.38758f
C607 avdd.t239 dvss 2.81531f
C608 avdd.n1112 dvss 1.38758f
C609 avdd.t369 dvss 2.81531f
C610 avdd.n1115 dvss 1.38758f
C611 avdd.n1118 dvss 1.38758f
C612 avdd.t365 dvss 2.81531f
C613 avdd.n1121 dvss 1.38758f
C614 avdd.t363 dvss 2.81531f
C615 avdd.n1126 dvss 1.38758f
C616 avdd.t349 dvss 2.81462f
C617 avdd.n1129 dvss 1.38262f
C618 avdd.n1132 dvss 1.38262f
C619 avdd.t283 dvss 2.81462f
C620 avdd.n1135 dvss 1.38262f
C621 avdd.t276 dvss 2.81462f
C622 avdd.n1140 dvss 1.38262f
C623 avdd.n1142 dvss 1.98405f
C624 avdd.n1157 dvss 2.19884f
C625 avdd.t182 dvss 60.565098f
C626 avdd.t240 dvss 47.8713f
C627 avdd.n1160 dvss 1.40416f
C628 avdd.n1161 dvss 19.3239f
C629 avdd.n1162 dvss 1.17692f
C630 avdd.t267 dvss 2.83122f
C631 avdd.n1168 dvss 1.37069f
C632 avdd.n1171 dvss 2.02177f
C633 avdd.n1172 dvss 2.47268f
C634 avdd.n1173 dvss 1.94224f
C635 avdd.n1176 dvss 4.18315f
C636 avdd.n1177 dvss 15.9837f
C637 avdd.n1178 dvss 15.717299f
C638 avdd.n1179 dvss 15.9837f
C639 avdd.n1180 dvss 4.18315f
C640 avdd.n1183 dvss 1.94224f
C641 avdd.n1184 dvss 1.74935f
C642 avdd.n1185 dvss 1.93268f
C643 avdd.n1187 dvss 1.14544f
C644 avdd.n1188 dvss 1.90907f
C645 avdd.n1194 dvss 2.13204f
C646 avdd.n1195 dvss 30.2826f
C647 avdd.n1196 dvss 2.13204f
C648 avdd.n1197 dvss 1.24982f
C649 avdd.n1200 dvss 1.40416f
C650 avdd.n1201 dvss 19.3239f
C651 avdd.n1202 dvss 1.17692f
C652 avdd.t387 dvss 2.81531f
C653 avdd.n1207 dvss 1.38758f
C654 avdd.t334 dvss 2.81531f
C655 avdd.n1209 dvss 1.38758f
C656 avdd.t382 dvss 2.81531f
C657 avdd.n1211 dvss 1.38758f
C658 avdd.t321 dvss 2.81531f
C659 avdd.n1213 dvss 1.38758f
C660 avdd.t326 dvss 2.81531f
C661 avdd.n1215 dvss 1.38758f
C662 avdd.t311 dvss 2.81531f
C663 avdd.n1217 dvss 1.38758f
C664 avdd.t308 dvss 2.81531f
C665 avdd.n1219 dvss 1.38758f
C666 avdd.t288 dvss 2.81462f
C667 avdd.n1221 dvss 1.38262f
C668 avdd.t251 dvss 2.81462f
C669 avdd.n1223 dvss 1.38262f
C670 avdd.t254 dvss 2.81462f
C671 avdd.n1225 dvss 1.38262f
C672 avdd.t244 dvss 2.81462f
C673 avdd.n1227 dvss 1.38262f
C674 avdd.n1229 dvss 1.30446f
C675 avdd.n1231 dvss 1.03155f
C676 avdd.n1233 dvss 2.68905f
C677 avdd.t271 dvss 2.83122f
C678 avdd.n1234 dvss 1.37069f
C679 avdd.n1238 dvss 1.32443f
C680 avdd.n1239 dvss 1.40599f
C681 avdd.n1240 dvss 2.23246f
C682 avdd.t230 dvss 47.8713f
C683 avdd.n1242 dvss 2.67548f
C684 avdd.n1243 dvss 2.46292f
C685 avdd.n1244 dvss 1.52014f
C686 avdd.n1245 dvss 1.44595f
C687 avdd.t525 dvss 1.31907f
C688 avdd.t446 dvss 1.82555f
C689 avdd.n1251 dvss 1.61596f
C690 avdd.t519 dvss 1.50199f
C691 avdd.t527 dvss 1.65232f
C692 avdd.n1253 dvss 1.42336f
C693 avdd.n1258 dvss 2.11868f
C694 avdd.n1259 dvss 1.52014f
C695 avdd.t73 dvss 45.4238f
C696 avdd.t63 dvss 60.565098f
C697 avdd.t65 dvss 45.4238f
C698 avdd.n1260 dvss 1.40599f
C699 avdd.n1264 dvss 1.90355f
C700 avdd.n1265 dvss 1.76059f
C701 avdd.n1292 dvss 2.54367f
C702 avdd.n1296 dvss 4.16674f
C703 avdd.n1297 dvss 4.1662f
C704 avdd.n1298 dvss 15.7194f
C705 avdd.n1299 dvss 1.01273f
C706 avdd.n1302 dvss 1.77866f
C707 avdd.n1304 dvss 1.51886f
C708 avdd.n1310 dvss 2.80462f
C709 avdd.n1311 dvss 3.09468f
C710 avdd.n1312 dvss 2.79818f
C711 avdd.t24 dvss 1.14721f
C712 avdd.n1317 dvss 1.51918f
C713 avdd.t582 dvss 1.14721f
C714 avdd.n1318 dvss 1.51918f
C715 avdd.n1497 dvss 1.96012f
C716 avdd.n1518 dvss 3.57199f
C717 avdd.n1519 dvss 2.68905f
C718 avdd.t351 dvss 2.81462f
C719 avdd.t265 dvss 2.81531f
C720 avdd.t263 dvss 2.81531f
C721 avdd.n1525 dvss 1.38758f
C722 avdd.t294 dvss 2.81531f
C723 avdd.n1528 dvss 1.38758f
C724 avdd.t301 dvss 2.81531f
C725 avdd.n1533 dvss 1.38758f
C726 avdd.t319 dvss 2.81531f
C727 avdd.n1536 dvss 1.38758f
C728 avdd.n1539 dvss 1.38758f
C729 avdd.t324 dvss 2.81531f
C730 avdd.n1542 dvss 1.38758f
C731 avdd.t269 dvss 2.81531f
C732 avdd.n1547 dvss 1.38758f
C733 avdd.t343 dvss 2.81462f
C734 avdd.n1550 dvss 1.38262f
C735 avdd.n1553 dvss 1.38262f
C736 avdd.t345 dvss 2.81462f
C737 avdd.n1556 dvss 1.38262f
C738 avdd.t361 dvss 2.81462f
C739 avdd.n1561 dvss 1.38262f
C740 avdd.n1563 dvss 1.29008f
C741 avdd.n1564 dvss 5.64129f
C742 avdd.n1579 dvss 2.19884f
C743 avdd.t80 dvss 60.565098f
C744 avdd.t234 dvss 47.8713f
C745 avdd.n1582 dvss 1.40416f
C746 avdd.n1583 dvss 19.3239f
C747 avdd.n1584 dvss 1.17692f
C748 avdd.t233 dvss 2.83122f
C749 avdd.n1590 dvss 1.37069f
C750 avdd.n1593 dvss 2.02177f
C751 avdd.n1594 dvss 2.47268f
C752 avdd.n1595 dvss 1.94224f
C753 avdd.n1598 dvss 4.18315f
C754 avdd.n1599 dvss 15.9837f
C755 avdd.n1600 dvss 15.717299f
C756 avdd.n1601 dvss 15.9837f
C757 avdd.n1602 dvss 4.18315f
C758 avdd.n1605 dvss 1.94224f
C759 avdd.n1606 dvss 1.74935f
C760 avdd.n1607 dvss 1.93268f
C761 avdd.n1609 dvss 1.14544f
C762 avdd.n1610 dvss 1.90907f
C763 avdd.n1616 dvss 2.13204f
C764 avdd.n1617 dvss 30.2826f
C765 avdd.n1618 dvss 2.13204f
C766 avdd.n1619 dvss 1.24982f
C767 avdd.n1622 dvss 1.40416f
C768 avdd.n1623 dvss 19.3239f
C769 avdd.n1624 dvss 1.17692f
C770 avdd.t298 dvss 2.81531f
C771 avdd.n1629 dvss 1.38758f
C772 avdd.t353 dvss 2.81531f
C773 avdd.n1631 dvss 1.38758f
C774 avdd.t356 dvss 2.81531f
C775 avdd.n1633 dvss 1.38758f
C776 avdd.t371 dvss 2.81531f
C777 avdd.n1635 dvss 1.38758f
C778 avdd.t229 dvss 2.81531f
C779 avdd.n1637 dvss 1.38758f
C780 avdd.t278 dvss 2.81531f
C781 avdd.n1639 dvss 1.38758f
C782 avdd.t236 dvss 2.81531f
C783 avdd.n1641 dvss 1.38758f
C784 avdd.t285 dvss 2.81462f
C785 avdd.n1643 dvss 1.38262f
C786 avdd.t305 dvss 2.81462f
C787 avdd.n1645 dvss 1.38262f
C788 avdd.t291 dvss 2.81462f
C789 avdd.n1647 dvss 1.38262f
C790 avdd.t314 dvss 2.81462f
C791 avdd.n1649 dvss 1.38262f
C792 avdd.n1651 dvss 1.30446f
C793 avdd.n1653 dvss 1.03155f
C794 avdd.n1655 dvss 3.15606f
C795 avdd.n1656 dvss 5.12462f
C796 avdd.n1657 dvss 2.93435f
C797 avdd.n1658 dvss 1.89729f
C798 avdd.n1659 dvss 12.8817f
C799 avdd.n1660 dvss 9.06993f
C800 avdd.n1661 dvss 49.4963f
C801 avdd.n1662 dvss 42.2644f
C802 avdd.n1663 dvss 4.32748f
C803 avdd.n1664 dvss 4.62882f
C804 avdd.n1665 dvss 1.04951f
C805 avdd.n1666 dvss 6.41647f
C806 avdd.n1667 dvss 2.2627f
C807 avdd.n1668 dvss 8.686629f
C808 avdd.n1669 dvss 14.2293f
C809 avdd.n1670 dvss 3.65641f
C810 avdd.n1672 dvss 1.72911f
C811 avdd.n1673 dvss 7.02872f
C812 avdd.n1674 dvss 1.41053f
C813 avdd.n1675 dvss 7.84867f
C814 avdd.n1676 dvss 2.20022f
C815 avdd.n1677 dvss 2.2013f
C816 avdd.n1678 dvss 26.9724f
C817 avdd.n1679 dvss 7.04023f
C818 avdd.n1680 dvss 1.03048f
C819 avdd.n1681 dvss 1.03497f
C820 avdd.n1682 dvss 3.67326f
C821 avdd.n1683 dvss 3.63832f
C822 avdd.n1684 dvss 1.73296f
C823 avdd.n1686 dvss 5.18296f
C824 avdd.n1687 dvss 20.367401f
C825 avdd.n1688 dvss 33.481102f
C826 avdd.n1689 dvss 41.3242f
C827 avdd.n1690 dvss 9.97857f
C828 avdd.n1691 dvss 2.26189f
C829 avdd.n1692 dvss 2.62828f
C830 avdd.n1693 dvss 10.6368f
C831 avdd.n1694 dvss 9.92241f
C832 avdd.n1695 dvss 5.22348f
C833 avdd.n1696 dvss 2.40308f
C834 avdd.n1697 dvss 1.59228f
C835 avdd.n1698 dvss 5.74641f
C836 avdd.n1699 dvss 6.63089f
C837 avdd.n1700 dvss 1.05252f
C838 avdd.n1701 dvss 2.00936f
C839 avdd.n1702 dvss 5.18797f
C840 avdd.n1703 dvss 26.8078f
C841 avdd.n1704 dvss 34.7635f
C842 avdd.n1705 dvss 57.0747f
C843 avdd.n1706 dvss 14.862299f
C844 avdd.n1707 dvss 1.4718f
C845 avdd.n1708 dvss 2.30536f
C846 avdd.n1709 dvss 6.41203f
C847 avdd.n1710 dvss 3.70548f
C848 avdd.n1711 dvss 30.2797f
C849 avdd.n1712 dvss 70.8322f
C850 avdd.n1713 dvss 8.8336f
C851 avdd.n1714 dvss 1.92239f
C852 avdd.n1717 dvss 1.46895f
C853 avdd.n1718 dvss 1.37249f
C854 avdd.t488 dvss 4.57304f
C855 avdd.t97 dvss 2.28652f
C856 avdd.t434 dvss 5.88329f
C857 avdd.t228 dvss 4.57304f
C858 avdd.t491 dvss 4.57304f
C859 avdd.t505 dvss 3.08295f
C860 avdd.t95 dvss 2.86457f
C861 avdd.n1728 dvss 6.7311f
C862 avdd.t529 dvss 8.95339f
C863 avdd.t430 dvss 5.88329f
C864 avdd.t521 dvss 7.47614f
C865 avdd.n1730 dvss 1.51399f
C866 avdd.n1731 dvss 1.08238f
C867 avdd.n1735 dvss 1.05547f
C868 avdd.n1738 dvss 1.02013f
C869 avdd.n1740 dvss 1.39737f
C870 avdd.n1742 dvss 1.22482f
C871 avdd.t317 dvss 1.4131f
C872 avdd.n1746 dvss 2.94725f
C873 avdd.t534 dvss 3.1481f
C874 avdd.t489 dvss 8.22119f
C875 avdd.t523 dvss 8.68363f
C876 avdd.t225 dvss 4.66296f
C877 avdd.n1749 dvss 5.24101f
C878 avdd.t517 dvss 5.36946f
C879 avdd.n1750 dvss 3.20394f
C880 avdd.n1751 dvss 3.20394f
C881 avdd.n1752 dvss 1.87957f
C882 avdd.n1753 dvss 1.85982f
C883 avdd.n1754 dvss 1.80118f
C884 avdd.t533 dvss 3.49401f
C885 avdd.t338 dvss 4.57304f
C886 avdd.t531 dvss 4.57304f
C887 avdd.t506 dvss 5.15109f
C888 avdd.n1755 dvss 2.95449f
C889 avdd.t428 dvss 6.56091f
C890 avdd.t424 dvss 9.543679f
C891 avdd.t426 dvss 7.38165f
C892 avdd.n1756 dvss 4.9211f
C893 avdd.t432 dvss 7.38165f
C894 avdd.t330 dvss 9.8422f
C895 avdd.t400 dvss 9.8422f
C896 avdd.t402 dvss 9.8422f
C897 avdd.t341 dvss 9.8422f
C898 avdd.t404 dvss 9.8422f
C899 avdd.t406 dvss 9.8422f
C900 avdd.t258 dvss 8.27857f
C901 avdd.n1757 dvss 7.414411f
C902 avdd.n1760 dvss 2.91391f
C903 avdd.t329 dvss 4.41001f
C904 avdd.n1761 dvss 1.62921f
C905 avdd.n1762 dvss 1.80249f
C906 avdd.t257 dvss 4.51891f
C907 avdd.n1764 dvss 4.00524f
C908 avdd.n1767 dvss 1.47868f
C909 avdd.n1768 dvss 1.47868f
C910 avdd.t340 dvss 4.51079f
C911 avdd.n1771 dvss 3.97651f
C912 avdd.n1772 dvss 1.41766f
C913 avdd.n1775 dvss 1.47921f
C914 avdd.n1776 dvss 1.01812f
C915 avdd.n1778 dvss 1.79057f
C916 avdd.n1779 dvss 1.60607f
C917 avdd.n1780 dvss 1.77806f
C918 avdd.n1782 dvss 1.40626f
C919 avdd.n1784 dvss 1.9356f
C920 avdd.n1786 dvss 1.9356f
C921 avdd.n1787 dvss 1.47868f
C922 avdd.t224 dvss 4.51891f
C923 avdd.n1789 dvss 4.00524f
C924 avdd.n1791 dvss 3.29609f
C925 avdd.n1794 dvss 3.2239f
C926 avdd.n1795 dvss 3.28672f
C927 avdd.t318 dvss 2.71656f
C928 avdd.t515 dvss 9.428679f
C929 avdd.t348 dvss 3.36555f
C930 avdd.n1813 dvss 1.51296f
C931 avdd.n1814 dvss 2.19544f
C932 avdd.n1815 dvss 14.582801f
C933 avdd.n1816 dvss 30.6303f
C934 avdd.n1817 dvss 19.9303f
C935 avdd.n1835 dvss 1.02497f
C936 avdd.n1836 dvss 1.00624f
C937 avdd.n1842 dvss 3.0341f
C938 avdd.t454 dvss 2.36338f
C939 avdd.t468 dvss 1.95219f
C940 avdd.t484 dvss 1.95219f
C941 avdd.t464 dvss 1.95219f
C942 avdd.t480 dvss 1.95219f
C943 avdd.t476 dvss 1.95219f
C944 avdd.t458 dvss 1.95219f
C945 avdd.t472 dvss 1.46414f
C946 avdd.t456 dvss 1.46414f
C947 avdd.t470 dvss 1.95219f
C948 avdd.t466 dvss 1.95219f
C949 avdd.t482 dvss 1.95219f
C950 avdd.t462 dvss 1.95219f
C951 avdd.t478 dvss 1.95219f
C952 avdd.t460 dvss 1.95219f
C953 avdd.t474 dvss 2.36338f
C954 avdd.n1844 dvss 3.0341f
C955 avdd.n1847 dvss 1.07158f
C956 avdd.n1848 dvss 1.00518f
C957 avdd.n1850 dvss 1.36396f
C958 avdd.n1851 dvss 1.1527f
C959 avdd.n1852 dvss 1.08071f
C960 avdd.n1853 dvss 1.79526f
C961 avdd.n1854 dvss 1.07713f
C962 avdd.n1857 dvss 4.1896f
C963 avdd.t416 dvss 2.36338f
C964 avdd.t415 dvss 1.95219f
C965 avdd.t304 dvss 1.95219f
C966 avdd.t94 dvss 1.95219f
C967 avdd.t93 dvss 1.95219f
C968 avdd.t243 dvss 1.95219f
C969 avdd.t579 dvss 1.95219f
C970 avdd.t578 dvss 1.95219f
C971 avdd.t333 dvss 1.95219f
C972 avdd.t497 dvss 1.95219f
C973 avdd.t496 dvss 1.95219f
C974 avdd.t275 dvss 1.95219f
C975 avdd.t444 dvss 1.95219f
C976 avdd.t445 dvss 1.95219f
C977 avdd.t375 dvss 1.95219f
C978 avdd.t138 dvss 1.95219f
C979 avdd.t137 dvss 1.95219f
C980 avdd.t262 dvss 1.95219f
C981 avdd.t176 dvss 1.95219f
C982 avdd.t175 dvss 1.95219f
C983 avdd.t393 dvss 1.95219f
C984 avdd.t508 dvss 1.95219f
C985 avdd.t507 dvss 1.95219f
C986 avdd.t381 dvss 1.95219f
C987 avdd.t4 dvss 1.95219f
C988 avdd.t5 dvss 1.95219f
C989 avdd.t368 dvss 1.95219f
C990 avdd.t451 dvss 1.95219f
C991 avdd.t450 dvss 1.95219f
C992 avdd.t379 dvss 1.95219f
C993 avdd.t157 dvss 1.95219f
C994 avdd.t158 dvss 1.95219f
C995 avdd.t297 dvss 1.95219f
C996 avdd.t109 dvss 1.95219f
C997 avdd.t110 dvss 1.95219f
C998 avdd.t391 dvss 1.95219f
C999 avdd.t171 dvss 1.95219f
C1000 avdd.t172 dvss 1.95219f
C1001 avdd.t395 dvss 1.95219f
C1002 avdd.t627 dvss 1.95219f
C1003 avdd.t628 dvss 1.95219f
C1004 avdd.t360 dvss 1.95219f
C1005 avdd.t414 dvss 1.95219f
C1006 avdd.t413 dvss 1.95219f
C1007 avdd.t248 dvss 1.95219f
C1008 avdd.t139 dvss 1.95219f
C1009 avdd.t140 dvss 2.36338f
C1010 avdd.n1858 dvss 4.1896f
C1011 avdd.n1862 dvss 1.28347f
C1012 rstring_mux_0.vtrip4.n2 dvss 1.18871f
C1013 rstring_mux_0.vtrip4.n6 dvss 1.88678f
C1014 rstring_mux_0.vtrip4.n7 dvss 1.68899f
C1015 comparator_0.vinn.t56 dvss 2.07495f
C1016 comparator_0.vinn.t53 dvss 1.98572f
C1017 comparator_0.vinn.n38 dvss 1.65357f
C1018 comparator_0.vinn.t61 dvss 1.98572f
C1019 comparator_0.vinn.t58 dvss 1.98572f
C1020 comparator_0.vinn.t49 dvss 1.98572f
C1021 comparator_0.vinn.t59 dvss 1.98572f
C1022 comparator_0.vinn.t55 dvss 1.98572f
C1023 comparator_0.vinn.t54 dvss 1.98572f
C1024 comparator_0.vinn.n44 dvss 1.03295f
C1025 comparator_0.vinn.t50 dvss 2.0927f
C1026 comparator_0.vinn.t62 dvss 2.00221f
C1027 comparator_0.vinn.n45 dvss 1.69074f
C1028 comparator_0.vinn.t57 dvss 2.00221f
C1029 comparator_0.vinn.t51 dvss 2.00221f
C1030 comparator_0.vinn.t60 dvss 2.00221f
C1031 comparator_0.vinn.t52 dvss 2.00221f
C1032 comparator_0.vinn.t48 dvss 2.00221f
C1033 comparator_0.vinn.t63 dvss 2.00221f
C1034 comparator_0.vinn.n52 dvss 3.5161f
C1035 comparator_0.vinn.n53 dvss 3.47781f
C1036 avss.n7 dvss 2.7103f
C1037 avss.t235 dvss 7.03977f
C1038 avss.n8 dvss 7.86722f
C1039 avss.t4 dvss 6.74374f
C1040 avss.t242 dvss 6.74374f
C1041 avss.t114 dvss 9.30791f
C1042 avss.t334 dvss 9.692531f
C1043 avss.t259 dvss 11.7439f
C1044 avss.t318 dvss 9.692531f
C1045 avss.t70 dvss 5.87193f
C1046 avss.n18 dvss 9.692531f
C1047 avss.t264 dvss 5.87193f
C1048 avss.t316 dvss 9.692531f
C1049 avss.t321 dvss 9.66689f
C1050 avss.t120 dvss 3.53854f
C1051 avss.t303 dvss 8.23096f
C1052 avss.t8 dvss 9.30791f
C1053 avss.t277 dvss 5.58987f
C1054 avss.n26 dvss 2.06484f
C1055 avss.n27 dvss 1.04658f
C1056 avss.t145 dvss 4.16769f
C1057 avss.n28 dvss 1.57338f
C1058 avss.n33 dvss 1.27709f
C1059 avss.n34 dvss 1.27709f
C1060 avss.t166 dvss 4.16769f
C1061 avss.n36 dvss 1.57338f
C1062 avss.t180 dvss 4.16769f
C1063 avss.n41 dvss 1.57338f
C1064 avss.t332 dvss 2.10261f
C1065 avss.t328 dvss 9.692531f
C1066 avss.t276 dvss 6.61553f
C1067 avss.t221 dvss 7.58992f
C1068 avss.n46 dvss 6.61553f
C1069 avss.n47 dvss 1.11125f
C1070 avss.n48 dvss 1.11125f
C1071 avss.n49 dvss 8.43383f
C1072 avss.t305 dvss 4.94883f
C1073 avss.n50 dvss 1.75517f
C1074 avss.n51 dvss 1.75517f
C1075 avss.n52 dvss 1.75517f
C1076 avss.n53 dvss 2.78756f
C1077 avss.n54 dvss 1.75702f
C1078 avss.t403 dvss 1.3887f
C1079 avss.t261 dvss 7.43774f
C1080 avss.n66 dvss 1.75702f
C1081 avss.n67 dvss 55.223396f
C1082 avss.t402 dvss 9.77267f
C1083 avss.t106 dvss 11.6901f
C1084 avss.t270 dvss 11.6901f
C1085 avss.t9 dvss 11.6901f
C1086 avss.t132 dvss 11.5818f
C1087 avss.t237 dvss 11.6901f
C1088 avss.t257 dvss 11.6901f
C1089 avss.t260 dvss 11.6901f
C1090 avss.t41 dvss 11.6901f
C1091 avss.t404 dvss 11.6901f
C1092 avss.t241 dvss 11.6901f
C1093 avss.t322 dvss 11.6901f
C1094 avss.t387 dvss 11.6901f
C1095 avss.t62 dvss 11.6901f
C1096 avss.t407 dvss 5.95329f
C1097 avss.n68 dvss 68.496895f
C1098 avss.n69 dvss 40.796898f
C1099 avss.n308 dvss 13.6537f
C1100 avss.n321 dvss 6.87897f
C1101 avss.t20 dvss 10.0988f
C1102 avss.t249 dvss 10.0988f
C1103 avss.t11 dvss 10.0988f
C1104 avss.t240 dvss 10.0988f
C1105 avss.t105 dvss 10.0988f
C1106 avss.t320 dvss 10.0988f
C1107 avss.t5 dvss 10.0988f
C1108 avss.t115 dvss 10.6197f
C1109 avss.n322 dvss 5.77505f
C1110 avss.t116 dvss 5.22652f
C1111 avss.n341 dvss 5.84504f
C1112 avss.t238 dvss 3.44827f
C1113 avss.t313 dvss 5.535779f
C1114 avss.t314 dvss 3.06169f
C1115 avss.t250 dvss 2.75243f
C1116 avss.t188 dvss 5.1956f
C1117 avss.t298 dvss 3.40188f
C1118 avss.t251 dvss 2.75243f
C1119 avss.t299 dvss 4.85541f
C1120 avss.t157 dvss 3.74207f
C1121 avss.t275 dvss 2.75243f
C1122 avss.t338 dvss 2.92252f
C1123 avss.n342 dvss 2.75243f
C1124 avss.t339 dvss 2.92252f
C1125 avss.t236 dvss 2.75243f
C1126 avss.t197 dvss 4.17503f
C1127 avss.t255 dvss 4.42244f
C1128 avss.t42 dvss 2.75243f
C1129 avss.t252 dvss 3.83484f
C1130 avss.t143 dvss 4.76263f
C1131 avss.t243 dvss 2.75243f
C1132 avss.t76 dvss 3.49466f
C1133 avss.t77 dvss 5.10282f
C1134 avss.t2 dvss 2.75243f
C1135 avss.t161 dvss 3.15447f
C1136 avss.t398 dvss 5.443009f
C1137 avss.t113 dvss 2.75243f
C1138 avss.t395 dvss 2.81428f
C1139 avss.t152 dvss 5.50486f
C1140 avss.t308 dvss 3.03076f
C1141 avss.t405 dvss 2.75243f
C1142 avss.t309 dvss 5.22652f
C1143 avss.t139 dvss 3.37095f
C1144 avss.t1 dvss 2.75243f
C1145 avss.t102 dvss 4.88633f
C1146 avss.t99 dvss 3.71114f
C1147 avss.t269 dvss 2.75243f
C1148 avss.t159 dvss 4.54615f
C1149 avss.t375 dvss 4.05133f
C1150 avss.t97 dvss 2.75243f
C1151 avss.t374 dvss 4.20596f
C1152 avss.t184 dvss 4.39152f
C1153 avss.t13 dvss 2.75243f
C1154 avss.t19 dvss 3.86577f
C1155 avss.t16 dvss 4.7317f
C1156 avss.t386 dvss 2.75243f
C1157 avss.t208 dvss 3.52558f
C1158 avss.t381 dvss 5.07189f
C1159 avss.t262 dvss 2.75243f
C1160 avss.t380 dvss 3.1854f
C1161 avss.t212 dvss 5.41208f
C1162 avss.t63 dvss 2.75243f
C1163 avss.t72 dvss 2.84521f
C1164 avss.t75 dvss 5.50486f
C1165 avss.t206 dvss 2.99984f
C1166 avss.t7 dvss 2.75243f
C1167 avss.t24 dvss 5.25745f
C1168 avss.t21 dvss 3.34003f
C1169 avss.t61 dvss 2.75243f
C1170 avss.t216 dvss 4.91726f
C1171 avss.t247 dvss 3.68021f
C1172 avss.t66 dvss 2.75243f
C1173 avss.t248 dvss 4.57707f
C1174 avss.t210 dvss 4.0204f
C1175 avss.t258 dvss 2.75243f
C1176 avss.t93 dvss 4.23688f
C1177 avss.t94 dvss 4.36059f
C1178 avss.t244 dvss 2.75243f
C1179 avss.t150 dvss 3.8967f
C1180 avss.t266 dvss 4.700779f
C1181 avss.t233 dvss 2.75243f
C1182 avss.t265 dvss 4.25235f
C1183 avss.n343 dvss 5.04096f
C1184 avss.n348 dvss 1.10722f
C1185 avss.n349 dvss 3.14083f
C1186 avss.n351 dvss 1.43901f
C1187 avss.n352 dvss 1.283f
C1188 avss.n353 dvss 1.0984f
C1189 avss.n355 dvss 3.90688f
C1190 avss.t146 dvss 0.151748p
C1191 avss.t0 dvss 16.6336f
C1192 avss.n362 dvss 3.35439f
C1193 avss.n363 dvss 30.591002f
C1194 avss.t231 dvss 1.09033f
C1195 avss.t273 dvss 5.6687f
C1196 avss.t141 dvss 5.15396f
C1197 avss.n368 dvss 1.93072f
C1198 avss.n369 dvss 11.9005f
C1199 avss.n370 dvss 37.942303f
C1200 avss.n376 dvss 1.12284f
C1201 avss.t111 dvss 1.15849f
C1202 avss.t48 dvss 3.68438f
C1203 avss.n378 dvss 3.38361f
C1204 avss.n398 dvss 2.19837f
C1205 avss.t176 dvss 1.13638f
C1206 avss.n439 dvss 2.10206f
C1207 avss.n443 dvss 2.11702f
C1208 avss.n444 dvss 2.10206f
C1209 avss.n445 dvss 2.11702f
C1210 avss.t169 dvss 1.1846f
C1211 avss.n473 dvss 1.5803f
C1212 avss.n507 dvss 1.47018f
C1213 avss.n514 dvss 1.44335f
C1214 avss.n530 dvss 1.52582f
C1215 avss.n537 dvss 3.80011f
C1216 avss.n538 dvss 14.4679f
C1217 avss.t426 dvss 1.76078f
C1218 avss.n539 dvss 1.7372f
C1219 avss.t192 dvss 1.13638f
C1220 avss.n548 dvss 1.18285f
C1221 avss.t325 dvss 2.17246f
C1222 avss.n562 dvss 2.90041f
C1223 avss.t384 dvss 1.24373f
C1224 avss.n563 dvss 9.61362f
C1225 avss.n564 dvss 47.927197f
C1226 avss.n565 dvss 1.57146f
C1227 avss.n570 dvss 1.08013f
C1228 avss.n575 dvss 1.10033f
C1229 avss.n578 dvss 1.52524f
C1230 avss.t15 dvss 1.47902f
C1231 avss.t3 dvss 1.47902f
C1232 avss.t98 dvss 1.47902f
C1233 avss.t360 dvss 1.15548f
C1234 avss.t342 dvss 1.47902f
C1235 avss.t370 dvss 1.47902f
C1236 avss.t364 dvss 1.47902f
C1237 avss.t71 dvss 4.60652f
C1238 avss.n633 dvss 2.17231f
C1239 avss.n642 dvss 2.54206f
C1240 avss.t356 dvss 1.47902f
C1241 avss.n643 dvss 1.89499f
C1242 avss.n644 dvss 2.21852f
C1243 avss.n645 dvss 1.98743f
C1244 avss.n656 dvss 1.52524f
C1245 avss.n657 dvss 2.35718f
C1246 avss.t366 dvss 1.47902f
C1247 avss.n658 dvss 2.4034f
C1248 avss.t368 dvss 1.47902f
C1249 avss.n659 dvss 1.2017f
C1250 avss.t310 dvss 1.47902f
C1251 avss.n660 dvss 1.2017f
C1252 avss.n676 dvss 1.71011f
C1253 avss.n677 dvss 1.98743f
C1254 avss.n678 dvss 1.61767f
C1255 avss.n679 dvss 2.26474f
C1256 avss.n697 dvss 2.4034f
C1257 avss.t352 dvss 1.47902f
C1258 avss.t10 dvss 1.47902f
C1259 avss.t346 dvss 1.24792f
C1260 avss.n699 dvss 1.57145f
C1261 avss.n702 dvss 1.66389f
C1262 avss.t358 dvss 1.47902f
C1263 avss.n703 dvss 1.80255f
C1264 avss.n704 dvss 1.52524f
C1265 avss.n717 dvss 2.07987f
C1266 avss.n718 dvss 1.80255f
C1267 avss.t350 dvss 1.47902f
C1268 avss.t362 dvss 1.47902f
C1269 avss.n720 dvss 2.4034f
C1270 avss.n731 dvss 1.94121f
C1271 avss.t344 dvss 1.47902f
C1272 avss.n732 dvss 2.26474f
C1273 avss.n733 dvss 1.47902f
C1274 avss.t354 dvss 1.47902f
C1275 avss.n734 dvss 1.61767f
C1276 avss.n745 dvss 2.71153f
C1277 avss.t80 dvss 1.47902f
C1278 avss.n746 dvss 1.58686f
C1279 avss.t82 dvss 1.47902f
C1280 avss.n748 dvss 2.29556f
C1281 avss.n761 dvss 1.69471f
C1282 avss.t84 dvss 1.47902f
C1283 avss.n762 dvss 2.4034f
C1284 avss.t86 dvss 1.47902f
C1285 avss.t234 dvss 1.47902f
C1286 avss.n763 dvss 1.72552f
C1287 avss.n774 dvss 2.85019f
C1288 avss.t388 dvss 1.38658f
C1289 avss.n794 dvss 1.01948f
C1290 avss.t171 dvss 7.18523f
C1291 avss.t170 dvss 1.13638f
C1292 avss.t178 dvss 1.13638f
C1293 avss.t434 dvss 1.76078f
C1294 avss.t410 dvss 1.76078f
C1295 avss.t423 dvss 1.76078f
C1296 avss.t444 dvss 1.76078f
C1297 avss.t421 dvss 1.76078f
C1298 avss.t428 dvss 1.76078f
C1299 avss.t440 dvss 1.76078f
C1300 avss.t282 dvss 9.0905f
C1301 avss.t280 dvss 6.81788f
C1302 avss.t193 dvss 7.18523f
C1303 avss.t284 dvss 9.0905f
C1304 avss.t278 dvss 6.81788f
C1305 avss.n826 dvss 4.54525f
C1306 avss.n829 dvss 3.02453f
C1307 avss.n836 dvss 1.57202f
C1308 avss.n842 dvss 2.81938f
C1309 avss.t302 dvss 7.16399f
C1310 avss.t104 dvss 11.6473f
C1311 avss.t409 dvss 11.6473f
C1312 avss.t401 dvss 11.6473f
C1313 avss.t60 dvss 11.6473f
C1314 avss.t6 dvss 7.93431f
C1315 avss.t65 dvss 9.73687f
C1316 avss.t103 dvss 11.6473f
C1317 avss.t256 dvss 11.6473f
C1318 avss.t69 dvss 9.53658f
C1319 avss.n843 dvss 35.0856f
C1320 avss.t327 dvss 2.07038f
C1321 avss.n844 dvss 33.2797f
C1322 avss.n845 dvss 19.873098f
C1323 avss.n846 dvss 15.552501f
C1324 avss.t67 dvss 23.9649f
C1325 avss.t200 dvss 1.84674f
C1326 avss.n853 dvss 1.63541f
C1327 avss.t144 dvss 2.36498f
C1328 avss.n855 dvss 1.88667f
C1329 avss.t164 dvss 1.84674f
C1330 avss.n856 dvss 1.63541f
C1331 avss.t131 dvss 4.98317f
C1332 avss.t130 dvss 6.11728f
C1333 avss.t129 dvss 6.11728f
C1334 avss.t128 dvss 51.730602f
C1335 avss.n867 dvss 1.0955f
C1336 avss.n872 dvss 22.547098f
C1337 avss.n873 dvss 17.083199f
C1338 avss.n881 dvss 24.1913f
C1339 avss.n882 dvss 31.336498f
C1340 avss.n883 dvss 16.0328f
C1341 avss.n884 dvss 1.39611f
C1342 avss.t290 dvss 2.19799f
C1343 avss.t286 dvss 1.23457f
C1344 avss.n885 dvss 1.13568f
C1345 avss.n893 dvss 2.19837f
C1346 avss.n898 dvss 1.26555f
C1347 avss.t202 dvss 1.13638f
C1348 avss.t430 dvss 1.74842f
C1349 avss.t417 dvss 1.74842f
C1350 avss.t411 dvss 1.74842f
C1351 avss.t436 dvss 1.74842f
C1352 avss.t412 dvss 1.74842f
C1353 avss.t437 dvss 1.74842f
C1354 avss.t419 dvss 1.74842f
C1355 avss.t415 dvss 1.74842f
C1356 avss.n913 dvss 4.01308f
C1357 avss.n914 dvss 11.1563f
C1358 avss.n915 dvss 12.5098f
C1359 avss.n920 dvss 4.50696f
C1360 avss.n921 dvss 6.85339f
C1361 avss.t153 dvss 1.13638f
C1362 avss.n934 dvss 1.26555f
C1363 avss.t217 dvss 1.13638f
C1364 avss.t435 dvss 1.74842f
C1365 avss.t438 dvss 1.74842f
C1366 avss.t442 dvss 1.74842f
C1367 avss.t424 dvss 1.74842f
C1368 avss.t441 dvss 1.74842f
C1369 avss.t414 dvss 1.74842f
C1370 avss.t432 dvss 1.74842f
C1371 avss.t439 dvss 1.74842f
C1372 avss.n949 dvss 6.94092f
C1373 avss.t427 dvss 1.76078f
C1374 avss.n950 dvss 1.7372f
C1375 avss.t420 dvss 1.76078f
C1376 avss.t443 dvss 1.76078f
C1377 avss.t431 dvss 1.76078f
C1378 avss.t413 dvss 1.76078f
C1379 avss.t433 dvss 1.76078f
C1380 avss.t425 dvss 1.76078f
C1381 avss.t422 dvss 1.76078f
C1382 avss.t133 dvss 1.13638f
C1383 avss.n969 dvss 1.18285f
C1384 avss.t109 dvss 2.60214f
C1385 avss.t271 dvss 3.80237f
C1386 avss.n979 dvss 3.17247f
C1387 avss.t46 dvss 2.75009f
C1388 avss.t88 dvss 3.17247f
C1389 avss.t50 dvss 4.31247f
C1390 avss.t58 dvss 4.36165f
C1391 avss.n981 dvss 1.58624f
C1392 avss.n990 dvss 3.9745f
C1393 avss.n996 dvss 4.418241f
C1394 avss.n997 dvss 35.3597f
C1395 avss.n998 dvss 39.5265f
C1396 avss.n1004 dvss 7.85272f
C1397 avss.n1005 dvss 4.8794f
C1398 avss.n1007 dvss 1.53339f
C1399 avss.n1008 dvss 1.5511f
C1400 avss.n1009 dvss 2.8965f
C1401 avss.n1010 dvss 2.88997f
C1402 avss.n1011 dvss 1.75517f
C1403 avss.n1012 dvss 1.75702f
C1404 avss.n1013 dvss 1.75702f
C1405 avss.n1014 dvss 1.69234f
C1406 avss.t117 dvss -1.14726f
C1407 avss.t214 dvss 5.20525f
C1408 avss.t323 dvss 4.56421f
C1409 avss.t337 dvss 6.79503f
C1410 avss.t186 dvss 7.46171f
C1411 avss.t43 dvss 4.56421f
C1412 avss.t336 dvss 6.23091f
C1413 avss.t324 dvss 4.69241f
C1414 avss.n1016 dvss 1.11045f
C1415 avss.n1017 dvss 3.46162f
C1416 avss.n1018 dvss 1.11045f
C1417 avss.n1022 dvss 1.27709f
C1418 avss.n1023 dvss 1.27709f
C1419 avss.t198 dvss 4.16769f
C1420 avss.n1025 dvss 1.57338f
C1421 avss.t162 dvss 4.16769f
C1422 avss.n1030 dvss 1.57338f
C1423 avss.n1032 dvss 1.27709f
C1424 avss.n1034 dvss 1.27709f
C1425 avss.t189 dvss 4.16769f
C1426 avss.n1035 dvss 1.57338f
C1427 avss.n1041 dvss 1.04658f
C1428 avss.n1042 dvss 1.04658f
C1429 avss.t225 dvss 4.16769f
C1430 avss.n1044 dvss 1.57338f
C1431 avss.n1047 dvss 1.27709f
C1432 avss.n1048 dvss 1.27709f
C1433 avss.t135 dvss 4.16769f
C1434 avss.n1050 dvss 1.57338f
C1435 avss.t228 dvss 4.16769f
C1436 avss.n1055 dvss 1.57338f
C1437 avss.n1057 dvss 1.27709f
C1438 avss.n1059 dvss 1.27709f
C1439 avss.t222 dvss 4.16769f
C1440 avss.n1060 dvss 1.57338f
C1441 avss.n1066 dvss 1.06639f
C1442 avss.n1067 dvss 1.10583f
C1443 avss.n1074 dvss 6.53861f
C1444 avss.n1075 dvss 7.43607f
C1445 avss.n1088 dvss 2.2821f
C1446 avss.t136 dvss 6.17963f
C1447 avss.n1089 dvss 7.41043f
C1448 avss.n1095 dvss 9.692531f
C1449 avss.t14 dvss 13.3336f
C1450 avss.t68 dvss 10.9233f
C1451 avss.n1096 dvss 20.644001f
C1452 avss.t394 dvss 17.866999f
C1453 avss.t64 dvss 15.7068f
C1454 avss.t12 dvss 15.849701f
C1455 avss.t107 dvss 15.849701f
C1456 avss.t232 dvss 15.849701f
C1457 avss.t239 dvss 15.849701f
C1458 avss.t263 dvss 12.7259f
C1459 avss.n1097 dvss 17.8087f
C1460 avss.n1098 dvss 12.420401f
C1461 avss.t296 dvss 2.80633f
.ends

