magic
tech sky130A
magscale 1 2
timestamp 1713454396
<< dnwell >>
rect -438 -2037 10654 2526
<< nwell >>
rect -357 6707 -341 6741
rect 10311 5341 11035 7579
rect -518 2320 10734 2606
rect -518 -1831 -232 2320
rect 10448 -1831 10734 2320
rect -518 -2117 10734 -1831
<< pwell >>
rect -386 4445 -322 4606
rect -515 4381 -322 4445
rect -515 3689 -451 4337
<< nsubdiff >>
rect -481 2549 10697 2569
rect -481 2515 -401 2549
rect 10617 2515 10697 2549
rect -481 2495 10697 2515
rect -481 2489 -407 2495
rect -481 -2000 -461 2489
rect -427 -2000 -407 2489
rect -481 -2006 -407 -2000
rect 10623 2489 10697 2495
rect 10623 -2000 10643 2489
rect 10677 -2000 10697 2489
rect 10623 -2006 10697 -2000
rect -481 -2026 10697 -2006
rect -481 -2060 -401 -2026
rect 10617 -2060 10697 -2026
rect -481 -2080 10697 -2060
<< nsubdiffcont >>
rect -401 2515 10617 2549
rect -461 -2000 -427 2489
rect 10643 -2000 10677 2489
rect -401 -2060 10617 -2026
<< locali >>
rect -173 7467 -17 7501
rect -173 5839 -17 5873
rect 102 5091 166 5106
rect 102 5057 117 5091
rect 151 5057 166 5091
rect 102 5042 166 5057
rect 1760 5091 1824 5106
rect 1760 5057 1775 5091
rect 1809 5057 1824 5091
rect 1760 5042 1824 5057
rect 5076 5091 5140 5106
rect 5076 5057 5091 5091
rect 5125 5057 5140 5091
rect 5076 5042 5140 5057
rect 8392 5091 8456 5106
rect 8392 5057 8407 5091
rect 8441 5057 8456 5091
rect 8392 5042 8456 5057
rect 10050 5091 10114 5106
rect 10050 5057 10065 5091
rect 10099 5057 10114 5091
rect 10050 5042 10114 5057
rect 10739 7501 10803 7516
rect 10739 7467 10754 7501
rect 10788 7467 10803 7501
rect 10739 7452 10803 7467
rect 10739 5453 10803 5468
rect 10739 5419 10754 5453
rect 10788 5419 10803 5453
rect 10739 5404 10803 5419
rect 102 4557 166 4572
rect 5076 4557 5140 4572
rect 10050 4557 10114 4572
rect 102 4523 117 4557
rect 10099 4523 10114 4557
rect 102 4508 166 4523
rect 5076 4508 5140 4523
rect 10050 4508 10114 4523
rect 10421 4406 10485 4421
rect 10421 4288 10436 4406
rect 10470 4288 10485 4406
rect 10421 4273 10485 4288
rect 10945 4406 11009 4421
rect 10945 4288 10960 4406
rect 10994 4288 11009 4406
rect 10945 4273 11009 4288
rect 102 4168 166 4183
rect 1760 4168 1824 4183
rect 5076 4168 5140 4183
rect 8392 4168 8456 4183
rect 10050 4168 10114 4183
rect -203 4134 -17 4168
rect 102 4134 117 4168
rect 10099 4134 10114 4168
rect 102 4119 166 4134
rect 1760 4119 1824 4134
rect 5076 4119 5140 4134
rect 8392 4119 8456 4134
rect 10050 4119 10114 4134
rect 102 3288 166 3303
rect 1760 3288 1824 3303
rect 5076 3288 5140 3303
rect 8392 3288 8456 3303
rect 10050 3288 10114 3303
rect -203 3254 -17 3288
rect 102 3254 117 3288
rect 10099 3254 10114 3288
rect 102 3239 166 3254
rect 1760 3239 1824 3254
rect 5076 3239 5140 3254
rect 8392 3239 8456 3254
rect 10050 3239 10114 3254
rect 1456 2549 1520 2564
rect 5230 2549 5294 2564
rect 8696 2549 8760 2564
rect -461 2515 -401 2549
rect 10617 2515 10677 2549
rect -461 2489 -427 2515
rect 1456 2500 1520 2515
rect 5230 2500 5294 2515
rect 8696 2500 8760 2515
rect 10643 2489 10677 2515
rect -461 -2026 -427 -2000
rect 1456 -2026 1520 -2011
rect 5230 -2026 5294 -2011
rect 8696 -2026 8760 -2011
rect 10643 -2026 10677 -2000
rect -461 -2060 -401 -2026
rect 10617 -2060 10677 -2026
rect 1456 -2075 1520 -2060
rect 5230 -2075 5294 -2060
rect 8696 -2075 8760 -2060
<< viali >>
rect 79 9409 10137 9443
rect -17 4598 17 9347
rect 79 7781 10137 7815
rect 117 5057 151 5091
rect 1775 5057 1809 5091
rect 5091 5057 5125 5091
rect 8407 5057 8441 5091
rect 10065 5057 10099 5091
rect 10199 4646 10233 9347
rect 10754 7467 10788 7501
rect 10754 5419 10788 5453
rect 117 4523 10099 4557
rect 10436 4288 10470 4406
rect 10960 4288 10994 4406
rect 117 4134 10099 4168
rect 117 3254 10099 3288
rect -307 2515 10040 2549
rect -461 -1929 -427 2426
rect 79 2078 10137 2112
rect -17 -1338 17 2016
rect 10199 -1338 10233 2016
rect 79 -1434 10137 -1400
rect 10643 -1968 10677 2387
rect 50 -2060 10397 -2026
<< metal1 >>
rect -32 9443 10248 9458
rect -32 9409 79 9443
rect 10137 9409 10248 9443
rect -32 9394 10248 9409
rect -32 9347 32 9394
rect -614 7223 -550 7229
rect -614 7171 -608 7223
rect -556 7171 -550 7223
rect -614 7165 -550 7171
rect -356 7223 -292 7229
rect -356 7171 -350 7223
rect -298 7171 -292 7223
rect -356 7165 -292 7171
rect -485 7115 -421 7121
rect -485 7063 -479 7115
rect -427 7063 -421 7115
rect -485 7057 -421 7063
rect -614 6858 -550 6864
rect -614 6806 -608 6858
rect -556 6806 -550 6858
rect -614 6800 -550 6806
rect -356 6858 -292 6864
rect -356 6806 -350 6858
rect -298 6806 -292 6858
rect -356 6800 -292 6806
rect -485 6750 -421 6756
rect -485 6698 -479 6750
rect -427 6698 -421 6750
rect -485 6692 -421 6698
rect -614 6493 -550 6499
rect -614 6441 -608 6493
rect -556 6441 -550 6493
rect -614 6435 -550 6441
rect -356 6481 -292 6487
rect -356 6429 -350 6481
rect -298 6429 -292 6481
rect -356 6423 -292 6429
rect -485 6385 -421 6391
rect -485 6333 -479 6385
rect -427 6333 -421 6385
rect -485 6327 -421 6333
rect -614 6116 -550 6122
rect -614 6064 -608 6116
rect -556 6064 -550 6116
rect -614 6058 -550 6064
rect -356 6116 -292 6122
rect -356 6064 -350 6116
rect -298 6064 -292 6116
rect -356 6058 -292 6064
rect -485 6020 -421 6026
rect -485 5968 -479 6020
rect -427 5968 -421 6020
rect -485 5962 -421 5968
rect -515 5107 -451 5113
rect -515 5055 -509 5107
rect -457 5055 -451 5107
rect -515 5049 -451 5055
rect -644 5020 -580 5026
rect -644 4968 -638 5020
rect -586 4968 -580 5020
rect -644 4962 -580 4968
rect -386 5020 -322 5026
rect -386 4968 -380 5020
rect -328 4968 -322 5020
rect -386 4962 -322 4968
rect -567 4751 -503 4757
rect -567 4699 -561 4751
rect -509 4699 -503 4751
rect -567 4693 -503 4699
rect -386 4664 -322 4670
rect -386 4612 -380 4664
rect -328 4612 -322 4664
rect -386 4606 -322 4612
rect -32 4598 -17 9347
rect 17 7827 32 9347
rect 10184 9347 10248 9394
rect 6743 9169 6789 9255
rect 102 9163 166 9169
rect 102 9111 108 9163
rect 160 9111 166 9163
rect 102 9105 166 9111
rect 1760 9163 1824 9169
rect 1760 9111 1766 9163
rect 1818 9111 1824 9163
rect 1760 9105 1824 9111
rect 3418 9162 3482 9168
rect 3418 9110 3424 9162
rect 3476 9110 3482 9162
rect 3418 9104 3482 9110
rect 5076 9163 5140 9169
rect 5076 9111 5082 9163
rect 5134 9111 5140 9163
rect 5076 9105 5140 9111
rect 6734 9163 6798 9169
rect 6734 9111 6740 9163
rect 6792 9111 6798 9163
rect 6734 9105 6798 9111
rect 8392 9163 8456 9169
rect 8392 9111 8398 9163
rect 8450 9111 8456 9163
rect 8392 9105 8456 9111
rect 10050 9163 10114 9169
rect 10050 9111 10056 9163
rect 10108 9111 10114 9163
rect 10050 9105 10114 9111
rect 111 9054 157 9095
rect 3427 9054 3473 9095
rect 6743 9054 6789 9105
rect 10059 9054 10105 9095
rect 111 9022 167 9054
rect 3417 9008 3483 9054
rect 6733 9008 6799 9054
rect 10049 9022 10105 9054
rect 102 8798 166 8804
rect 102 8746 108 8798
rect 160 8746 166 8798
rect 102 8740 166 8746
rect 1760 8798 1824 8804
rect 3427 8803 3473 9008
rect 6743 8804 6789 9008
rect 1760 8746 1766 8798
rect 1818 8746 1824 8798
rect 1760 8740 1824 8746
rect 3418 8797 3482 8803
rect 3418 8745 3424 8797
rect 3476 8745 3482 8797
rect 3418 8739 3482 8745
rect 5076 8798 5140 8804
rect 5076 8746 5082 8798
rect 5134 8746 5140 8798
rect 5076 8740 5140 8746
rect 6734 8798 6798 8804
rect 6734 8746 6740 8798
rect 6792 8746 6798 8798
rect 6734 8740 6798 8746
rect 8392 8798 8456 8804
rect 8392 8746 8398 8798
rect 8450 8746 8456 8798
rect 8392 8740 8456 8746
rect 10050 8798 10114 8804
rect 10050 8746 10056 8798
rect 10108 8746 10114 8798
rect 10050 8740 10114 8746
rect 111 8689 157 8730
rect 3427 8689 3473 8739
rect 6743 8689 6789 8740
rect 10059 8689 10105 8730
rect 111 8657 167 8689
rect 3417 8643 3483 8689
rect 6733 8643 6799 8689
rect 10049 8657 10105 8689
rect 102 8433 166 8439
rect 102 8381 108 8433
rect 160 8381 166 8433
rect 102 8375 166 8381
rect 1760 8433 1824 8439
rect 3427 8438 3473 8643
rect 6743 8439 6789 8643
rect 1760 8381 1766 8433
rect 1818 8381 1824 8433
rect 1760 8375 1824 8381
rect 3418 8432 3482 8438
rect 3418 8380 3424 8432
rect 3476 8380 3482 8432
rect 3418 8374 3482 8380
rect 5076 8433 5140 8439
rect 5076 8381 5082 8433
rect 5134 8381 5140 8433
rect 5076 8375 5140 8381
rect 6734 8433 6798 8439
rect 6734 8381 6740 8433
rect 6792 8381 6798 8433
rect 6734 8375 6798 8381
rect 8392 8433 8456 8439
rect 8392 8381 8398 8433
rect 8450 8381 8456 8433
rect 8392 8375 8456 8381
rect 10050 8433 10114 8439
rect 10050 8381 10056 8433
rect 10108 8381 10114 8433
rect 10050 8375 10114 8381
rect 111 8324 157 8365
rect 3427 8324 3473 8374
rect 6743 8324 6789 8375
rect 10059 8324 10105 8365
rect 111 8292 167 8324
rect 3417 8278 3483 8324
rect 6733 8278 6799 8324
rect 10049 8292 10105 8324
rect 3427 8074 3473 8278
rect 6743 8200 6789 8278
rect 6743 8074 6789 8160
rect 102 8068 166 8074
rect 102 8016 108 8068
rect 160 8016 166 8068
rect 102 8010 166 8016
rect 1760 8068 1824 8074
rect 1760 8016 1766 8068
rect 1818 8016 1824 8068
rect 1760 8010 1824 8016
rect 3418 8068 3482 8074
rect 3418 8016 3424 8068
rect 3476 8016 3482 8068
rect 3418 8010 3482 8016
rect 5076 8068 5140 8074
rect 5076 8016 5082 8068
rect 5134 8016 5140 8068
rect 5076 8010 5140 8016
rect 6734 8068 6798 8074
rect 6734 8016 6740 8068
rect 6792 8016 6798 8068
rect 6734 8010 6798 8016
rect 8392 8068 8456 8074
rect 8392 8016 8398 8068
rect 8450 8016 8456 8068
rect 8392 8010 8456 8016
rect 10050 8068 10114 8074
rect 10050 8016 10056 8068
rect 10108 8016 10114 8068
rect 10050 8010 10114 8016
rect 111 7959 157 8000
rect 3427 7959 3473 8010
rect 6743 7959 6789 8010
rect 10059 7959 10105 8000
rect 111 7927 167 7959
rect 3417 7913 3483 7959
rect 6733 7913 6799 7959
rect 10049 7927 10105 7959
rect 10184 7827 10199 9347
rect 17 7815 10199 7827
rect 17 7781 79 7815
rect 10137 7781 10199 7815
rect 17 7769 10199 7781
rect 17 4598 32 7769
rect 102 7534 166 7540
rect 102 7482 108 7534
rect 160 7482 166 7534
rect 102 7476 166 7482
rect 1760 7534 1824 7540
rect 1760 7482 1766 7534
rect 1818 7482 1824 7534
rect 1760 7476 1824 7482
rect 3418 7534 3482 7540
rect 3418 7482 3424 7534
rect 3476 7482 3482 7534
rect 3418 7476 3482 7482
rect 5076 7534 5140 7540
rect 5076 7482 5082 7534
rect 5134 7482 5140 7534
rect 5076 7476 5140 7482
rect 6734 7534 6798 7540
rect 6734 7482 6740 7534
rect 6792 7482 6798 7534
rect 6734 7476 6798 7482
rect 8392 7534 8456 7540
rect 8392 7482 8398 7534
rect 8450 7482 8456 7534
rect 8392 7476 8456 7482
rect 10050 7534 10114 7540
rect 10050 7482 10056 7534
rect 10108 7482 10114 7534
rect 10050 7476 10114 7482
rect 111 7425 157 7466
rect 4300 7428 4364 7434
rect 111 7379 167 7425
rect 3417 7379 3483 7425
rect 4300 7376 4306 7428
rect 4358 7376 4364 7428
rect 4300 7370 4364 7376
rect 5956 7428 6020 7434
rect 5956 7376 5962 7428
rect 6014 7376 6020 7428
rect 10059 7425 10105 7466
rect 6733 7379 6799 7425
rect 10049 7379 10105 7425
rect 5956 7370 6020 7376
rect 102 7169 166 7175
rect 102 7117 108 7169
rect 160 7117 166 7169
rect 102 7111 166 7117
rect 1760 7169 1824 7175
rect 1760 7117 1766 7169
rect 1818 7117 1824 7169
rect 1760 7111 1824 7117
rect 3418 7169 3482 7175
rect 3418 7117 3424 7169
rect 3476 7117 3482 7169
rect 3418 7111 3482 7117
rect 5076 7169 5140 7175
rect 5076 7117 5082 7169
rect 5134 7117 5140 7169
rect 5076 7111 5140 7117
rect 6734 7169 6798 7175
rect 6734 7117 6740 7169
rect 6792 7117 6798 7169
rect 6734 7111 6798 7117
rect 8392 7169 8456 7175
rect 8392 7117 8398 7169
rect 8450 7117 8456 7169
rect 8392 7111 8456 7117
rect 10050 7169 10114 7175
rect 10050 7117 10056 7169
rect 10108 7117 10114 7169
rect 10050 7111 10114 7117
rect 111 7060 157 7101
rect 4300 7063 4364 7069
rect 111 7014 167 7060
rect 3417 7014 3483 7060
rect 4300 7011 4306 7063
rect 4358 7011 4364 7063
rect 4300 7005 4364 7011
rect 5956 7063 6020 7069
rect 5956 7011 5962 7063
rect 6014 7011 6020 7063
rect 10059 7060 10105 7101
rect 6733 7014 6799 7060
rect 10049 7014 10105 7060
rect 10184 7018 10199 7769
rect 5956 7005 6020 7011
rect 10169 6954 10199 7018
rect 102 6804 166 6810
rect 102 6752 108 6804
rect 160 6752 166 6804
rect 102 6746 166 6752
rect 1760 6804 1824 6810
rect 1760 6752 1766 6804
rect 1818 6752 1824 6804
rect 1760 6746 1824 6752
rect 3418 6804 3482 6810
rect 3418 6752 3424 6804
rect 3476 6752 3482 6804
rect 3418 6746 3482 6752
rect 5076 6804 5140 6810
rect 5076 6752 5082 6804
rect 5134 6752 5140 6804
rect 5076 6746 5140 6752
rect 6734 6804 6798 6810
rect 6734 6752 6740 6804
rect 6792 6752 6798 6804
rect 6734 6746 6798 6752
rect 8392 6804 8456 6810
rect 8392 6752 8398 6804
rect 8450 6752 8456 6804
rect 8392 6746 8456 6752
rect 10050 6804 10114 6810
rect 10050 6752 10056 6804
rect 10108 6752 10114 6804
rect 10050 6746 10114 6752
rect 111 6695 157 6736
rect 4300 6698 4364 6704
rect 111 6649 167 6695
rect 3417 6649 3483 6695
rect 4300 6646 4306 6698
rect 4358 6646 4364 6698
rect 4300 6640 4364 6646
rect 5956 6698 6020 6704
rect 5956 6646 5962 6698
rect 6014 6646 6020 6698
rect 10059 6695 10105 6736
rect 6733 6649 6799 6695
rect 10049 6649 10105 6695
rect 5956 6640 6020 6646
rect 102 6439 166 6445
rect 102 6387 108 6439
rect 160 6387 166 6439
rect 102 6381 166 6387
rect 1760 6439 1824 6445
rect 1760 6387 1766 6439
rect 1818 6387 1824 6439
rect 1760 6381 1824 6387
rect 3418 6439 3482 6445
rect 3418 6387 3424 6439
rect 3476 6387 3482 6439
rect 3418 6381 3482 6387
rect 5076 6439 5140 6445
rect 5076 6387 5082 6439
rect 5134 6387 5140 6439
rect 5076 6381 5140 6387
rect 6734 6439 6798 6445
rect 6734 6387 6740 6439
rect 6792 6387 6798 6439
rect 6734 6381 6798 6387
rect 8392 6439 8456 6445
rect 8392 6387 8398 6439
rect 8450 6387 8456 6439
rect 8392 6381 8456 6387
rect 10050 6439 10114 6445
rect 10050 6387 10056 6439
rect 10108 6387 10114 6439
rect 10050 6381 10114 6387
rect 111 6330 157 6371
rect 4300 6333 4364 6339
rect 111 6284 167 6330
rect 3417 6284 3483 6330
rect 4300 6281 4306 6333
rect 4358 6281 4364 6333
rect 4300 6275 4364 6281
rect 5956 6333 6020 6339
rect 5956 6281 5962 6333
rect 6014 6281 6020 6333
rect 10059 6330 10105 6371
rect 6733 6284 6799 6330
rect 10049 6284 10105 6330
rect 5956 6275 6020 6281
rect 102 6074 166 6080
rect 102 6022 108 6074
rect 160 6022 166 6074
rect 102 6016 166 6022
rect 1760 6074 1824 6080
rect 1760 6022 1766 6074
rect 1818 6022 1824 6074
rect 1760 6016 1824 6022
rect 3418 6074 3482 6080
rect 3418 6022 3424 6074
rect 3476 6022 3482 6074
rect 3418 6016 3482 6022
rect 5076 6074 5140 6080
rect 5076 6022 5082 6074
rect 5134 6022 5140 6074
rect 5076 6016 5140 6022
rect 6734 6074 6798 6080
rect 6734 6022 6740 6074
rect 6792 6022 6798 6074
rect 6734 6016 6798 6022
rect 8392 6074 8456 6080
rect 8392 6022 8398 6074
rect 8450 6022 8456 6074
rect 8392 6016 8456 6022
rect 10050 6074 10114 6080
rect 10050 6022 10056 6074
rect 10108 6022 10114 6074
rect 10050 6016 10114 6022
rect 111 5965 157 6006
rect 4300 5968 4364 5974
rect 111 5919 167 5965
rect 3417 5919 3483 5965
rect 4300 5916 4306 5968
rect 4358 5916 4364 5968
rect 4300 5910 4364 5916
rect 5956 5968 6020 5974
rect 5956 5916 5962 5968
rect 6014 5916 6020 5968
rect 10059 5965 10105 6006
rect 6733 5919 6799 5965
rect 10049 5919 10105 5965
rect 5956 5910 6020 5916
rect 102 5709 166 5715
rect 102 5657 108 5709
rect 160 5657 166 5709
rect 102 5651 166 5657
rect 1760 5709 1824 5715
rect 1760 5657 1766 5709
rect 1818 5657 1824 5709
rect 1760 5651 1824 5657
rect 3418 5709 3482 5715
rect 3418 5657 3424 5709
rect 3476 5657 3482 5709
rect 3418 5651 3482 5657
rect 5076 5709 5140 5715
rect 5076 5657 5082 5709
rect 5134 5657 5140 5709
rect 5076 5651 5140 5657
rect 6734 5709 6798 5715
rect 6734 5657 6740 5709
rect 6792 5657 6798 5709
rect 6734 5651 6798 5657
rect 8392 5709 8456 5715
rect 8392 5657 8398 5709
rect 8450 5657 8456 5709
rect 8392 5651 8456 5657
rect 10050 5709 10114 5715
rect 10050 5657 10056 5709
rect 10108 5657 10114 5709
rect 10050 5651 10114 5657
rect 111 5600 157 5641
rect 4300 5603 4364 5609
rect 111 5554 167 5600
rect 3417 5554 3483 5600
rect 4300 5551 4306 5603
rect 4358 5551 4364 5603
rect 4300 5545 4364 5551
rect 5956 5603 6020 5609
rect 5956 5551 5962 5603
rect 6014 5551 6020 5603
rect 10059 5600 10105 5641
rect 6733 5554 6799 5600
rect 10049 5554 10105 5600
rect 5956 5545 6020 5551
rect 102 5344 166 5350
rect 102 5292 108 5344
rect 160 5292 166 5344
rect 102 5286 166 5292
rect 1760 5344 1824 5350
rect 1760 5292 1766 5344
rect 1818 5292 1824 5344
rect 1760 5286 1824 5292
rect 3418 5344 3482 5350
rect 3418 5292 3424 5344
rect 3476 5292 3482 5344
rect 3418 5286 3482 5292
rect 5076 5344 5140 5350
rect 5076 5292 5082 5344
rect 5134 5292 5140 5344
rect 5076 5286 5140 5292
rect 6734 5344 6798 5350
rect 6734 5292 6740 5344
rect 6792 5292 6798 5344
rect 6734 5286 6798 5292
rect 8392 5344 8456 5350
rect 8392 5292 8398 5344
rect 8450 5292 8456 5344
rect 8392 5286 8456 5292
rect 10050 5344 10114 5350
rect 10050 5292 10056 5344
rect 10108 5292 10114 5344
rect 10050 5286 10114 5292
rect 111 5235 157 5276
rect 4300 5238 4364 5244
rect 111 5189 167 5235
rect 3417 5189 3483 5235
rect 4300 5186 4306 5238
rect 4358 5186 4364 5238
rect 4300 5180 4364 5186
rect 5956 5238 6020 5244
rect 5956 5186 5962 5238
rect 6014 5186 6020 5238
rect 10059 5235 10105 5276
rect 6733 5189 6799 5235
rect 10049 5189 10105 5235
rect 5956 5180 6020 5186
rect 102 5100 166 5106
rect 102 5048 108 5100
rect 160 5048 166 5100
rect 102 5042 166 5048
rect 1760 5100 1824 5106
rect 1760 5048 1766 5100
rect 1818 5048 1824 5100
rect 1760 5042 1824 5048
rect 5076 5100 5140 5106
rect 5076 5048 5082 5100
rect 5134 5048 5140 5100
rect 5076 5042 5140 5048
rect 8392 5100 8456 5106
rect 8392 5048 8398 5100
rect 8450 5048 8456 5100
rect 8392 5042 8456 5048
rect 10050 5100 10114 5106
rect 10050 5048 10056 5100
rect 10108 5048 10114 5100
rect 10050 5042 10114 5048
rect 102 4937 166 4943
rect 102 4885 108 4937
rect 160 4885 166 4937
rect 102 4879 166 4885
rect 1760 4937 1824 4943
rect 1760 4885 1766 4937
rect 1818 4885 1824 4937
rect 1760 4879 1824 4885
rect 5076 4937 5140 4943
rect 5076 4885 5082 4937
rect 5134 4885 5140 4937
rect 5076 4879 5140 4885
rect 8392 4937 8456 4943
rect 8392 4885 8398 4937
rect 8450 4885 8456 4937
rect 8392 4879 8456 4885
rect 10050 4937 10114 4943
rect 10050 4885 10056 4937
rect 10108 4885 10114 4937
rect 10050 4879 10114 4885
rect 3418 4807 3482 4813
rect 3418 4755 3424 4807
rect 3476 4755 3482 4807
rect 3418 4749 3482 4755
rect 6734 4807 6798 4813
rect 6734 4755 6740 4807
rect 6792 4755 6798 4807
rect 6734 4749 6798 4755
rect 111 4702 157 4743
rect 4300 4705 4364 4711
rect 111 4656 167 4702
rect 3417 4656 3483 4702
rect 4300 4653 4306 4705
rect 4358 4653 4364 4705
rect 4300 4647 4364 4653
rect 5956 4705 6020 4711
rect 5956 4653 5962 4705
rect 6014 4653 6020 4705
rect 10059 4702 10105 4743
rect 6733 4656 6799 4702
rect 10049 4656 10105 4702
rect 5956 4647 6020 4653
rect -32 4572 32 4598
rect 10184 4646 10199 6954
rect 10233 4646 10248 9347
rect 10739 7510 10803 7516
rect 10739 7458 10745 7510
rect 10797 7458 10803 7510
rect 10739 7452 10803 7458
rect 10739 7376 10803 7382
rect 10739 7324 10745 7376
rect 10797 7324 10803 7376
rect 10739 7318 10803 7324
rect 10522 6071 10568 7205
rect 10609 7198 10673 7204
rect 10609 7146 10615 7198
rect 10667 7146 10673 7198
rect 10609 7140 10673 7146
rect 10739 7020 10803 7026
rect 10739 6968 10745 7020
rect 10797 6968 10803 7020
rect 10739 6962 10803 6968
rect 10609 6842 10673 6848
rect 10609 6790 10615 6842
rect 10667 6790 10673 6842
rect 10609 6784 10673 6790
rect 10739 6664 10803 6670
rect 10739 6612 10745 6664
rect 10797 6612 10803 6664
rect 10739 6606 10803 6612
rect 10609 6486 10673 6492
rect 10609 6434 10615 6486
rect 10667 6434 10673 6486
rect 10609 6428 10673 6434
rect 10739 6308 10803 6314
rect 10739 6256 10745 6308
rect 10797 6256 10803 6308
rect 10739 6250 10803 6256
rect 10609 6130 10673 6136
rect 10609 6078 10615 6130
rect 10667 6078 10673 6130
rect 10609 6072 10673 6078
rect 10506 6007 10570 6013
rect 10506 5955 10512 6007
rect 10564 5955 10570 6007
rect 10506 5949 10570 5955
rect 10739 5952 10803 5958
rect 10739 5900 10745 5952
rect 10797 5900 10803 5952
rect 10739 5894 10803 5900
rect 10522 5715 10568 5781
rect 10609 5774 10673 5780
rect 10609 5722 10615 5774
rect 10667 5722 10673 5774
rect 10609 5716 10673 5722
rect 10508 5661 10572 5667
rect 10508 5609 10514 5661
rect 10566 5609 10572 5661
rect 10508 5603 10572 5609
rect 10739 5596 10803 5602
rect 10739 5544 10745 5596
rect 10797 5544 10803 5596
rect 10739 5538 10803 5544
rect 10739 5462 10803 5468
rect 10739 5410 10745 5462
rect 10797 5410 10803 5462
rect 10739 5404 10803 5410
rect 10774 5096 10838 5102
rect 10774 5044 10780 5096
rect 10832 5044 10838 5096
rect 10774 5038 10838 5044
rect 10184 4572 10248 4646
rect -32 4566 10248 4572
rect -644 4528 -580 4534
rect -644 4476 -638 4528
rect -586 4476 -580 4528
rect -32 4514 108 4566
rect 160 4557 1766 4566
rect 1818 4557 5082 4566
rect 5134 4557 10056 4566
rect 160 4514 1766 4523
rect 1818 4514 5082 4523
rect 5134 4514 10056 4523
rect 10108 4514 10248 4566
rect -32 4508 10248 4514
rect -644 4470 -580 4476
rect 10421 4415 10485 4421
rect -515 4395 -451 4401
rect -515 4343 -509 4395
rect -457 4343 -451 4395
rect -515 4337 -451 4343
rect 10421 4279 10427 4415
rect 10479 4279 10485 4415
rect 10421 4273 10485 4279
rect -386 4184 -322 4190
rect -644 4172 -580 4178
rect -644 4120 -638 4172
rect -586 4120 -580 4172
rect -386 4132 -380 4184
rect -328 4132 -322 4184
rect -386 4126 -322 4132
rect -32 4177 10248 4183
rect -644 4114 -580 4120
rect -32 4125 108 4177
rect 160 4168 1766 4177
rect 1818 4168 5082 4177
rect 5134 4168 8398 4177
rect 8450 4168 10056 4177
rect 160 4125 1766 4134
rect 1818 4125 5082 4134
rect 5134 4125 8398 4134
rect 8450 4125 10056 4134
rect 10108 4125 10248 4177
rect -32 4119 10248 4125
rect -515 4039 -451 4045
rect -515 3987 -509 4039
rect -457 3987 -451 4039
rect -515 3981 -451 3987
rect -386 3952 -322 3958
rect -386 3900 -380 3952
rect -328 3900 -322 3952
rect -386 3894 -322 3900
rect -644 3816 -580 3822
rect -644 3764 -638 3816
rect -586 3764 -580 3816
rect -644 3758 -580 3764
rect -515 3683 -451 3689
rect -515 3631 -509 3683
rect -457 3631 -451 3683
rect -515 3625 -451 3631
rect -386 3596 -322 3602
rect -386 3544 -380 3596
rect -327 3544 -322 3596
rect -386 3538 -322 3544
rect -644 3460 -580 3466
rect -644 3408 -638 3460
rect -586 3408 -580 3460
rect -644 3402 -580 3408
rect -32 3303 32 4119
rect 108 3990 167 4036
rect 3417 3990 3483 4036
rect 5075 3990 5141 4036
rect 6733 3990 6799 4036
rect 10049 3990 10108 4036
rect 108 3952 160 3990
rect 3427 3952 3473 3990
rect 10056 3952 10108 3990
rect 102 3946 166 3952
rect 102 3894 108 3946
rect 160 3894 166 3946
rect 102 3888 166 3894
rect 1760 3946 1824 3952
rect 1760 3894 1766 3946
rect 1818 3894 1824 3946
rect 1760 3888 1824 3894
rect 3418 3946 3482 3952
rect 3418 3894 3424 3946
rect 3476 3894 3482 3946
rect 3418 3888 3482 3894
rect 5076 3946 5140 3952
rect 5076 3894 5082 3946
rect 5134 3894 5140 3946
rect 5076 3888 5140 3894
rect 6734 3947 6798 3952
rect 6734 3894 6740 3947
rect 6792 3894 6798 3947
rect 6734 3888 6798 3894
rect 8392 3946 8456 3952
rect 8392 3894 8398 3946
rect 8450 3894 8456 3946
rect 8392 3888 8456 3894
rect 10050 3946 10114 3952
rect 10050 3894 10056 3946
rect 10108 3894 10114 3946
rect 10050 3888 10114 3894
rect 108 3634 167 3680
rect 3417 3634 3483 3680
rect 5075 3634 5141 3680
rect 6733 3634 6799 3680
rect 10049 3634 10108 3680
rect 108 3596 160 3634
rect 3427 3596 3473 3634
rect 10056 3596 10108 3634
rect 102 3590 166 3596
rect 102 3538 108 3590
rect 160 3538 166 3590
rect 102 3532 166 3538
rect 1760 3590 1824 3596
rect 1760 3538 1766 3590
rect 1818 3538 1824 3590
rect 1760 3532 1824 3538
rect 3418 3590 3482 3596
rect 3418 3538 3424 3590
rect 3476 3538 3482 3590
rect 3418 3532 3482 3538
rect 5076 3590 5140 3596
rect 5076 3538 5082 3590
rect 5134 3538 5140 3590
rect 5076 3532 5140 3538
rect 8392 3590 8456 3596
rect 8392 3538 8398 3590
rect 8450 3538 8456 3590
rect 8392 3532 8456 3538
rect 10050 3590 10114 3596
rect 10050 3538 10056 3590
rect 10108 3538 10114 3590
rect 10050 3532 10114 3538
rect 6734 3466 6798 3472
rect 6734 3414 6740 3466
rect 6792 3414 6798 3466
rect 6734 3408 6798 3414
rect 10184 3303 10248 4119
rect 10560 3791 10606 4925
rect 10643 4919 10707 4925
rect 10643 4867 10649 4919
rect 10701 4867 10707 4919
rect 10643 4861 10707 4867
rect 10774 4740 10838 4746
rect 10774 4688 10780 4740
rect 10832 4688 10838 4740
rect 10774 4682 10838 4688
rect 10643 4563 10707 4569
rect 10643 4511 10649 4563
rect 10701 4511 10707 4563
rect 10643 4505 10707 4511
rect 10945 4415 11009 4421
rect 10774 4384 10838 4390
rect 10774 4332 10780 4384
rect 10832 4332 10838 4384
rect 10774 4326 10838 4332
rect 10945 4279 10951 4415
rect 11003 4279 11009 4415
rect 10945 4273 11009 4279
rect 10643 4207 10707 4213
rect 10643 4155 10649 4207
rect 10701 4155 10707 4207
rect 10643 4149 10707 4155
rect 10774 4028 10838 4034
rect 10774 3976 10780 4028
rect 10832 3976 10838 4028
rect 10774 3970 10838 3976
rect 10643 3851 10707 3857
rect 10643 3799 10649 3851
rect 10701 3799 10707 3851
rect 10643 3793 10707 3799
rect 10539 3728 10603 3734
rect 10539 3676 10545 3728
rect 10597 3676 10603 3728
rect 10539 3670 10603 3676
rect 10774 3672 10838 3678
rect 10774 3620 10780 3672
rect 10832 3620 10838 3672
rect 10774 3614 10838 3620
rect 10545 3608 10609 3614
rect 10545 3556 10551 3608
rect 10603 3556 10609 3608
rect 10545 3550 10609 3556
rect 10560 3435 10606 3501
rect 10645 3494 10709 3500
rect 10645 3442 10651 3494
rect 10703 3442 10709 3494
rect 10645 3436 10709 3442
rect -32 3297 10248 3303
rect -32 3245 108 3297
rect 160 3288 1766 3297
rect 1818 3288 5082 3297
rect 5134 3288 8398 3297
rect 8450 3288 10056 3297
rect 160 3245 1766 3254
rect 1818 3245 5082 3254
rect 5134 3245 8398 3254
rect 8450 3245 10056 3254
rect 10108 3245 10248 3297
rect 10774 3316 10838 3322
rect 10774 3264 10780 3316
rect 10832 3264 10838 3316
rect 10774 3258 10838 3264
rect -32 3239 10248 3245
rect -476 2558 10692 2564
rect -476 2549 1462 2558
rect 1514 2549 5236 2558
rect 5288 2549 8702 2558
rect 8754 2549 10692 2558
rect -476 2515 -307 2549
rect 10040 2515 10692 2549
rect -476 2506 1462 2515
rect 1514 2506 5236 2515
rect 5288 2506 8702 2515
rect 8754 2506 10692 2515
rect -476 2500 10692 2506
rect -476 2426 -412 2500
rect -476 -1929 -461 2426
rect -427 -1929 -412 2426
rect 10628 2387 10692 2500
rect -29 2121 10245 2124
rect -29 2112 108 2121
rect 160 2112 3424 2121
rect 3476 2112 6740 2121
rect 6792 2112 10056 2121
rect 10108 2112 10245 2121
rect -29 2078 79 2112
rect 10137 2078 10245 2112
rect -29 2069 108 2078
rect 160 2069 3424 2078
rect 3476 2069 6740 2078
rect 6792 2069 10056 2078
rect 10108 2069 10245 2078
rect -29 2066 10245 2069
rect -29 2016 29 2066
rect -29 -1338 -17 2016
rect 17 -1338 29 2016
rect 10187 2016 10245 2066
rect 347 1983 411 1989
rect 9854 1983 9918 1989
rect 347 1931 353 1983
rect 405 1931 411 1983
rect 3138 1931 3144 1983
rect 3196 1931 3202 1983
rect 4725 1931 4731 1983
rect 4783 1931 4789 1983
rect 5075 1934 5141 1980
rect 6957 1931 6963 1983
rect 7015 1931 7021 1983
rect 9854 1931 9860 1983
rect 9912 1931 9918 1983
rect 347 1925 411 1931
rect 9854 1925 9918 1931
rect 102 1766 166 1772
rect 102 1714 108 1766
rect 160 1714 166 1766
rect 102 1708 166 1714
rect 1760 1766 1824 1772
rect 1760 1714 1766 1766
rect 1818 1714 1824 1766
rect 1760 1708 1824 1714
rect 3418 1766 3482 1772
rect 3418 1714 3424 1766
rect 3476 1714 3482 1766
rect 3418 1708 3482 1714
rect 5076 1766 5140 1772
rect 5076 1714 5082 1766
rect 5134 1714 5140 1766
rect 5076 1708 5140 1714
rect 6734 1766 6798 1772
rect 6734 1714 6740 1766
rect 6792 1714 6798 1766
rect 6734 1708 6798 1714
rect 8392 1766 8456 1772
rect 8392 1714 8398 1766
rect 8450 1714 8456 1766
rect 8392 1708 8456 1714
rect 10050 1766 10114 1772
rect 10050 1714 10056 1766
rect 10108 1714 10114 1766
rect 10050 1708 10114 1714
rect 347 1673 411 1679
rect 9854 1673 9918 1679
rect 347 1621 353 1673
rect 405 1621 411 1673
rect 3138 1621 3144 1673
rect 3196 1621 3202 1673
rect 4725 1621 4731 1673
rect 4783 1621 4789 1673
rect 5075 1624 5141 1670
rect 6957 1621 6963 1673
rect 7015 1621 7021 1673
rect 9854 1621 9860 1673
rect 9912 1621 9918 1673
rect 347 1615 411 1621
rect 9854 1615 9918 1621
rect 347 1565 411 1571
rect 9854 1565 9918 1571
rect 347 1513 353 1565
rect 405 1513 411 1565
rect 3138 1513 3144 1565
rect 3196 1513 3202 1565
rect 4725 1513 4731 1565
rect 4783 1513 4789 1565
rect 5075 1516 5141 1562
rect 6957 1513 6963 1565
rect 7015 1513 7021 1565
rect 9854 1513 9860 1565
rect 9912 1513 9918 1565
rect 347 1507 411 1513
rect 9854 1507 9918 1513
rect 102 1348 166 1354
rect 102 1296 108 1348
rect 160 1296 166 1348
rect 102 1290 166 1296
rect 1760 1348 1824 1354
rect 1760 1296 1766 1348
rect 1818 1296 1824 1348
rect 1760 1290 1824 1296
rect 3418 1348 3482 1354
rect 3418 1296 3424 1348
rect 3476 1296 3482 1348
rect 3418 1290 3482 1296
rect 5076 1348 5140 1354
rect 5076 1296 5082 1348
rect 5134 1296 5140 1348
rect 5076 1290 5140 1296
rect 6734 1348 6798 1354
rect 6734 1296 6740 1348
rect 6792 1296 6798 1348
rect 6734 1290 6798 1296
rect 8392 1348 8456 1354
rect 8392 1296 8398 1348
rect 8450 1296 8456 1348
rect 8392 1290 8456 1296
rect 10050 1348 10114 1354
rect 10050 1296 10056 1348
rect 10108 1296 10114 1348
rect 10050 1290 10114 1296
rect 347 1255 411 1261
rect 9854 1255 9918 1261
rect 347 1203 353 1255
rect 405 1203 411 1255
rect 3138 1203 3144 1255
rect 3196 1203 3202 1255
rect 4725 1203 4731 1255
rect 4783 1203 4789 1255
rect 5075 1206 5141 1252
rect 6957 1203 6963 1255
rect 7015 1203 7021 1255
rect 9854 1203 9860 1255
rect 9912 1203 9918 1255
rect 347 1197 411 1203
rect 9854 1197 9918 1203
rect 347 1147 411 1153
rect 9854 1147 9918 1153
rect 347 1095 353 1147
rect 405 1095 411 1147
rect 3138 1095 3144 1147
rect 3196 1095 3202 1147
rect 4725 1095 4731 1147
rect 4783 1095 4789 1147
rect 5075 1098 5141 1144
rect 6957 1095 6963 1147
rect 7015 1095 7021 1147
rect 9854 1095 9860 1147
rect 9912 1095 9918 1147
rect 347 1089 411 1095
rect 9854 1089 9918 1095
rect 102 930 166 936
rect 102 878 108 930
rect 160 878 166 930
rect 102 872 166 878
rect 1760 930 1824 936
rect 1760 878 1766 930
rect 1818 878 1824 930
rect 1760 872 1824 878
rect 3418 930 3482 936
rect 3418 878 3424 930
rect 3476 878 3482 930
rect 3418 872 3482 878
rect 5076 930 5140 936
rect 5076 878 5082 930
rect 5134 878 5140 930
rect 5076 872 5140 878
rect 6734 930 6798 936
rect 6734 878 6740 930
rect 6792 878 6798 930
rect 6734 872 6798 878
rect 8392 930 8456 936
rect 8392 878 8398 930
rect 8450 878 8456 930
rect 8392 872 8456 878
rect 10050 930 10114 936
rect 10050 878 10056 930
rect 10108 878 10114 930
rect 10050 872 10114 878
rect 347 837 411 843
rect 9854 837 9918 843
rect 347 785 353 837
rect 405 785 411 837
rect 3138 785 3144 837
rect 3196 785 3202 837
rect 4725 785 4731 837
rect 4783 785 4789 837
rect 5075 788 5141 834
rect 6957 785 6963 837
rect 7015 785 7021 837
rect 9854 785 9860 837
rect 9912 785 9918 837
rect 347 779 411 785
rect 9854 779 9918 785
rect 347 729 411 735
rect 9854 729 9918 735
rect 347 677 353 729
rect 405 677 411 729
rect 3138 677 3144 729
rect 3196 677 3202 729
rect 4725 677 4731 729
rect 4783 677 4789 729
rect 5075 680 5141 726
rect 6957 677 6963 729
rect 7015 677 7021 729
rect 9854 677 9860 729
rect 9912 677 9918 729
rect 347 671 411 677
rect 9854 671 9918 677
rect 102 512 166 518
rect 102 460 108 512
rect 160 460 166 512
rect 102 454 166 460
rect 1760 512 1824 518
rect 1760 460 1766 512
rect 1818 460 1824 512
rect 1760 454 1824 460
rect 3418 512 3482 518
rect 3418 460 3424 512
rect 3476 460 3482 512
rect 3418 454 3482 460
rect 5076 512 5140 518
rect 5076 460 5082 512
rect 5134 460 5140 512
rect 5076 454 5140 460
rect 6734 512 6798 518
rect 6734 460 6740 512
rect 6792 460 6798 512
rect 6734 454 6798 460
rect 8392 512 8456 518
rect 8392 460 8398 512
rect 8450 460 8456 512
rect 8392 454 8456 460
rect 10050 512 10114 518
rect 10050 460 10056 512
rect 10108 460 10114 512
rect 10050 454 10114 460
rect 347 419 411 425
rect 9854 419 9918 425
rect 347 367 353 419
rect 405 367 411 419
rect 3138 367 3144 419
rect 3196 367 3202 419
rect 4725 367 4731 419
rect 4783 367 4789 419
rect 5075 370 5141 416
rect 6957 367 6963 419
rect 7015 367 7021 419
rect 9854 367 9860 419
rect 9912 367 9918 419
rect 347 361 411 367
rect 9854 361 9918 367
rect 347 311 411 317
rect 9854 311 9918 317
rect 347 259 353 311
rect 405 259 411 311
rect 3138 259 3144 311
rect 3196 259 3202 311
rect 4725 259 4731 311
rect 4783 259 4789 311
rect 5075 262 5141 308
rect 6957 259 6963 311
rect 7015 259 7021 311
rect 9854 259 9860 311
rect 9912 259 9918 311
rect 347 253 411 259
rect 9854 253 9918 259
rect 102 94 166 100
rect 102 42 108 94
rect 160 42 166 94
rect 102 36 166 42
rect 1760 94 1824 100
rect 1760 42 1766 94
rect 1818 42 1824 94
rect 1760 36 1824 42
rect 3418 94 3482 100
rect 3418 42 3424 94
rect 3476 42 3482 94
rect 3418 36 3482 42
rect 5076 94 5140 100
rect 5076 42 5082 94
rect 5134 42 5140 94
rect 5076 36 5140 42
rect 6734 94 6798 100
rect 6734 42 6740 94
rect 6792 42 6798 94
rect 6734 36 6798 42
rect 8392 94 8456 100
rect 8392 42 8398 94
rect 8450 42 8456 94
rect 8392 36 8456 42
rect 10050 94 10114 100
rect 10050 42 10056 94
rect 10108 42 10114 94
rect 10050 36 10114 42
rect 347 1 411 7
rect 9854 1 9918 7
rect 347 -51 353 1
rect 405 -51 411 1
rect 3138 -51 3144 1
rect 3196 -51 3202 1
rect 4725 -51 4731 1
rect 4783 -51 4789 1
rect 5075 -48 5141 -2
rect 6957 -51 6963 1
rect 7015 -51 7021 1
rect 9854 -51 9860 1
rect 9912 -51 9918 1
rect 347 -57 411 -51
rect 9854 -57 9918 -51
rect 347 -107 411 -101
rect 9854 -107 9918 -101
rect 347 -159 353 -107
rect 405 -159 411 -107
rect 3138 -159 3144 -107
rect 3196 -159 3202 -107
rect 4725 -159 4731 -107
rect 4783 -159 4789 -107
rect 5075 -156 5141 -110
rect 6957 -159 6963 -107
rect 7015 -159 7021 -107
rect 9854 -159 9860 -107
rect 9912 -159 9918 -107
rect 347 -165 411 -159
rect 9854 -165 9918 -159
rect 102 -324 166 -318
rect 102 -376 108 -324
rect 160 -376 166 -324
rect 102 -382 166 -376
rect 1760 -324 1824 -318
rect 1760 -376 1766 -324
rect 1818 -376 1824 -324
rect 1760 -382 1824 -376
rect 3418 -324 3482 -318
rect 3418 -376 3424 -324
rect 3476 -376 3482 -324
rect 3418 -382 3482 -376
rect 5076 -324 5140 -318
rect 5076 -376 5082 -324
rect 5134 -376 5140 -324
rect 5076 -382 5140 -376
rect 6734 -324 6798 -318
rect 6734 -376 6740 -324
rect 6792 -376 6798 -324
rect 6734 -382 6798 -376
rect 8392 -324 8456 -318
rect 8392 -376 8398 -324
rect 8450 -376 8456 -324
rect 8392 -382 8456 -376
rect 10050 -324 10114 -318
rect 10050 -376 10056 -324
rect 10108 -376 10114 -324
rect 10050 -382 10114 -376
rect 347 -417 411 -411
rect 9854 -417 9918 -411
rect 347 -469 353 -417
rect 405 -469 411 -417
rect 3138 -469 3144 -417
rect 3196 -469 3202 -417
rect 4725 -469 4731 -417
rect 4783 -469 4789 -417
rect 5075 -466 5141 -420
rect 6957 -469 6963 -417
rect 7015 -469 7021 -417
rect 9854 -469 9860 -417
rect 9912 -469 9918 -417
rect 347 -475 411 -469
rect 9854 -475 9918 -469
rect 347 -525 411 -519
rect 9854 -525 9918 -519
rect 347 -577 353 -525
rect 405 -577 411 -525
rect 3138 -577 3144 -525
rect 3196 -577 3202 -525
rect 4725 -577 4731 -525
rect 4783 -577 4789 -525
rect 5075 -574 5141 -528
rect 6957 -577 6963 -525
rect 7015 -577 7021 -525
rect 9854 -577 9860 -525
rect 9912 -577 9918 -525
rect 347 -583 411 -577
rect 9854 -583 9918 -577
rect 102 -742 166 -736
rect 102 -794 108 -742
rect 160 -794 166 -742
rect 102 -800 166 -794
rect 1760 -742 1824 -736
rect 1760 -794 1766 -742
rect 1818 -794 1824 -742
rect 1760 -800 1824 -794
rect 3418 -742 3482 -736
rect 3418 -794 3424 -742
rect 3476 -794 3482 -742
rect 3418 -800 3482 -794
rect 5076 -742 5140 -736
rect 5076 -794 5082 -742
rect 5134 -794 5140 -742
rect 5076 -800 5140 -794
rect 6734 -742 6798 -736
rect 6734 -794 6740 -742
rect 6792 -794 6798 -742
rect 6734 -800 6798 -794
rect 8392 -742 8456 -736
rect 8392 -794 8398 -742
rect 8450 -794 8456 -742
rect 8392 -800 8456 -794
rect 10050 -742 10114 -736
rect 10050 -794 10056 -742
rect 10108 -794 10114 -742
rect 10050 -800 10114 -794
rect 347 -835 411 -829
rect 9854 -835 9918 -829
rect 347 -887 353 -835
rect 405 -887 411 -835
rect 3138 -887 3144 -835
rect 3196 -887 3202 -835
rect 4725 -887 4731 -835
rect 4783 -887 4789 -835
rect 5075 -884 5141 -838
rect 6957 -887 6963 -835
rect 7015 -887 7021 -835
rect 9854 -887 9860 -835
rect 9912 -887 9918 -835
rect 347 -893 411 -887
rect 9854 -893 9918 -887
rect 347 -943 411 -937
rect 9854 -943 9918 -937
rect 347 -995 353 -943
rect 405 -995 411 -943
rect 3138 -995 3144 -943
rect 3196 -995 3202 -943
rect 4725 -995 4731 -943
rect 4783 -995 4789 -943
rect 5075 -992 5141 -946
rect 6957 -995 6963 -943
rect 7015 -995 7021 -943
rect 9854 -995 9860 -943
rect 9912 -995 9918 -943
rect 347 -1001 411 -995
rect 9854 -1001 9918 -995
rect 102 -1160 166 -1154
rect 102 -1212 108 -1160
rect 160 -1212 166 -1160
rect 102 -1218 166 -1212
rect 1760 -1160 1824 -1154
rect 1760 -1212 1766 -1160
rect 1818 -1212 1824 -1160
rect 1760 -1218 1824 -1212
rect 3418 -1160 3482 -1154
rect 3418 -1212 3424 -1160
rect 3476 -1212 3482 -1160
rect 3418 -1218 3482 -1212
rect 5076 -1160 5140 -1154
rect 5076 -1212 5082 -1160
rect 5134 -1212 5140 -1160
rect 5076 -1218 5140 -1212
rect 6734 -1160 6798 -1154
rect 6734 -1212 6740 -1160
rect 6792 -1212 6798 -1160
rect 6734 -1218 6798 -1212
rect 8392 -1160 8456 -1154
rect 8392 -1212 8398 -1160
rect 8450 -1212 8456 -1160
rect 8392 -1218 8456 -1212
rect 10050 -1160 10114 -1154
rect 10050 -1212 10056 -1160
rect 10108 -1212 10114 -1160
rect 10050 -1218 10114 -1212
rect 347 -1253 411 -1247
rect 9854 -1253 9918 -1247
rect 347 -1305 353 -1253
rect 405 -1305 411 -1253
rect 3138 -1305 3144 -1253
rect 3196 -1305 3202 -1253
rect 4725 -1305 4731 -1253
rect 4783 -1305 4789 -1253
rect 5075 -1302 5141 -1256
rect 6957 -1305 6963 -1253
rect 7015 -1305 7021 -1253
rect 9854 -1305 9860 -1253
rect 9912 -1305 9918 -1253
rect 347 -1311 411 -1305
rect 9854 -1311 9918 -1305
rect -29 -1388 29 -1338
rect 10187 -1338 10199 2016
rect 10233 -1338 10245 2016
rect 10187 -1388 10245 -1338
rect -29 -1391 10245 -1388
rect -29 -1400 108 -1391
rect 160 -1400 3424 -1391
rect 3476 -1400 6740 -1391
rect 6792 -1400 10056 -1391
rect 10108 -1400 10245 -1391
rect -29 -1434 79 -1400
rect 10137 -1434 10245 -1400
rect -29 -1443 108 -1434
rect 160 -1443 3424 -1434
rect 3476 -1443 6740 -1434
rect 6792 -1443 10056 -1434
rect 10108 -1443 10245 -1434
rect -29 -1446 10245 -1443
rect -476 -2011 -412 -1929
rect 10628 -1968 10643 2387
rect 10677 -1968 10692 2387
rect 10628 -2011 10692 -1968
rect -476 -2017 10692 -2011
rect -476 -2026 1462 -2017
rect 1514 -2026 5236 -2017
rect 5288 -2026 8702 -2017
rect 8754 -2026 10692 -2017
rect -476 -2060 50 -2026
rect 10397 -2060 10692 -2026
rect -476 -2069 1462 -2060
rect 1514 -2069 5236 -2060
rect 5288 -2069 8702 -2060
rect 8754 -2069 10692 -2060
rect -476 -2075 10692 -2069
<< via1 >>
rect -608 7171 -556 7223
rect -350 7171 -298 7223
rect -479 7063 -427 7115
rect -608 6806 -556 6858
rect -350 6806 -298 6858
rect -479 6698 -427 6750
rect -608 6441 -556 6493
rect -350 6429 -298 6481
rect -479 6333 -427 6385
rect -608 6064 -556 6116
rect -350 6064 -298 6116
rect -479 5968 -427 6020
rect -509 5055 -457 5107
rect -638 4968 -586 5020
rect -380 4968 -328 5020
rect -561 4699 -509 4751
rect -380 4612 -328 4664
rect 108 9111 160 9163
rect 1766 9111 1818 9163
rect 3424 9110 3476 9162
rect 5082 9111 5134 9163
rect 6740 9111 6792 9163
rect 8398 9111 8450 9163
rect 10056 9111 10108 9163
rect 108 8746 160 8798
rect 1766 8746 1818 8798
rect 3424 8745 3476 8797
rect 5082 8746 5134 8798
rect 6740 8746 6792 8798
rect 8398 8746 8450 8798
rect 10056 8746 10108 8798
rect 108 8381 160 8433
rect 1766 8381 1818 8433
rect 3424 8380 3476 8432
rect 5082 8381 5134 8433
rect 6740 8381 6792 8433
rect 8398 8381 8450 8433
rect 10056 8381 10108 8433
rect 108 8016 160 8068
rect 1766 8016 1818 8068
rect 3424 8016 3476 8068
rect 5082 8016 5134 8068
rect 6740 8016 6792 8068
rect 8398 8016 8450 8068
rect 10056 8016 10108 8068
rect 108 7482 160 7534
rect 1766 7482 1818 7534
rect 3424 7482 3476 7534
rect 5082 7482 5134 7534
rect 6740 7482 6792 7534
rect 8398 7482 8450 7534
rect 10056 7482 10108 7534
rect 4306 7376 4358 7428
rect 5962 7376 6014 7428
rect 108 7117 160 7169
rect 1766 7117 1818 7169
rect 3424 7117 3476 7169
rect 5082 7117 5134 7169
rect 6740 7117 6792 7169
rect 8398 7117 8450 7169
rect 10056 7117 10108 7169
rect 4306 7011 4358 7063
rect 5962 7011 6014 7063
rect 108 6752 160 6804
rect 1766 6752 1818 6804
rect 3424 6752 3476 6804
rect 5082 6752 5134 6804
rect 6740 6752 6792 6804
rect 8398 6752 8450 6804
rect 10056 6752 10108 6804
rect 4306 6646 4358 6698
rect 5962 6646 6014 6698
rect 108 6387 160 6439
rect 1766 6387 1818 6439
rect 3424 6387 3476 6439
rect 5082 6387 5134 6439
rect 6740 6387 6792 6439
rect 8398 6387 8450 6439
rect 10056 6387 10108 6439
rect 4306 6281 4358 6333
rect 5962 6281 6014 6333
rect 108 6022 160 6074
rect 1766 6022 1818 6074
rect 3424 6022 3476 6074
rect 5082 6022 5134 6074
rect 6740 6022 6792 6074
rect 8398 6022 8450 6074
rect 10056 6022 10108 6074
rect 4306 5916 4358 5968
rect 5962 5916 6014 5968
rect 108 5657 160 5709
rect 1766 5657 1818 5709
rect 3424 5657 3476 5709
rect 5082 5657 5134 5709
rect 6740 5657 6792 5709
rect 8398 5657 8450 5709
rect 10056 5657 10108 5709
rect 4306 5551 4358 5603
rect 5962 5551 6014 5603
rect 108 5292 160 5344
rect 1766 5292 1818 5344
rect 3424 5292 3476 5344
rect 5082 5292 5134 5344
rect 6740 5292 6792 5344
rect 8398 5292 8450 5344
rect 10056 5292 10108 5344
rect 4306 5186 4358 5238
rect 5962 5186 6014 5238
rect 108 5091 160 5100
rect 108 5057 117 5091
rect 117 5057 151 5091
rect 151 5057 160 5091
rect 108 5048 160 5057
rect 1766 5091 1818 5100
rect 1766 5057 1775 5091
rect 1775 5057 1809 5091
rect 1809 5057 1818 5091
rect 1766 5048 1818 5057
rect 5082 5091 5134 5100
rect 5082 5057 5091 5091
rect 5091 5057 5125 5091
rect 5125 5057 5134 5091
rect 5082 5048 5134 5057
rect 8398 5091 8450 5100
rect 8398 5057 8407 5091
rect 8407 5057 8441 5091
rect 8441 5057 8450 5091
rect 8398 5048 8450 5057
rect 10056 5091 10108 5100
rect 10056 5057 10065 5091
rect 10065 5057 10099 5091
rect 10099 5057 10108 5091
rect 10056 5048 10108 5057
rect 108 4885 160 4937
rect 1766 4885 1818 4937
rect 5082 4885 5134 4937
rect 8398 4885 8450 4937
rect 10056 4885 10108 4937
rect 3424 4755 3476 4807
rect 6740 4755 6792 4807
rect 4306 4653 4358 4705
rect 5962 4653 6014 4705
rect 10745 7501 10797 7510
rect 10745 7467 10754 7501
rect 10754 7467 10788 7501
rect 10788 7467 10797 7501
rect 10745 7458 10797 7467
rect 10745 7324 10797 7376
rect 10615 7146 10667 7198
rect 10745 6968 10797 7020
rect 10615 6790 10667 6842
rect 10745 6612 10797 6664
rect 10615 6434 10667 6486
rect 10745 6256 10797 6308
rect 10615 6078 10667 6130
rect 10512 5955 10564 6007
rect 10745 5900 10797 5952
rect 10615 5722 10667 5774
rect 10514 5609 10566 5661
rect 10745 5544 10797 5596
rect 10745 5453 10797 5462
rect 10745 5419 10754 5453
rect 10754 5419 10788 5453
rect 10788 5419 10797 5453
rect 10745 5410 10797 5419
rect 10780 5044 10832 5096
rect -638 4476 -586 4528
rect 108 4557 160 4566
rect 1766 4557 1818 4566
rect 5082 4557 5134 4566
rect 10056 4557 10108 4566
rect 108 4523 117 4557
rect 117 4523 160 4557
rect 1766 4523 1818 4557
rect 5082 4523 5134 4557
rect 10056 4523 10099 4557
rect 10099 4523 10108 4557
rect 108 4514 160 4523
rect 1766 4514 1818 4523
rect 5082 4514 5134 4523
rect 10056 4514 10108 4523
rect -509 4343 -457 4395
rect 10427 4406 10479 4415
rect 10427 4288 10436 4406
rect 10436 4288 10470 4406
rect 10470 4288 10479 4406
rect 10427 4279 10479 4288
rect -638 4120 -586 4172
rect -380 4132 -328 4184
rect 108 4168 160 4177
rect 1766 4168 1818 4177
rect 5082 4168 5134 4177
rect 8398 4168 8450 4177
rect 10056 4168 10108 4177
rect 108 4134 117 4168
rect 117 4134 160 4168
rect 1766 4134 1818 4168
rect 5082 4134 5134 4168
rect 8398 4134 8450 4168
rect 10056 4134 10099 4168
rect 10099 4134 10108 4168
rect 108 4125 160 4134
rect 1766 4125 1818 4134
rect 5082 4125 5134 4134
rect 8398 4125 8450 4134
rect 10056 4125 10108 4134
rect -509 3987 -457 4039
rect -380 3900 -328 3952
rect -638 3764 -586 3816
rect -509 3631 -457 3683
rect -380 3544 -327 3596
rect -638 3408 -586 3460
rect 108 3894 160 3946
rect 1766 3894 1818 3946
rect 3424 3894 3476 3946
rect 5082 3894 5134 3946
rect 6740 3894 6792 3947
rect 8398 3894 8450 3946
rect 10056 3894 10108 3946
rect 108 3538 160 3590
rect 1766 3538 1818 3590
rect 3424 3538 3476 3590
rect 5082 3538 5134 3590
rect 8398 3538 8450 3590
rect 10056 3538 10108 3590
rect 6740 3414 6792 3466
rect 10649 4867 10701 4919
rect 10780 4688 10832 4740
rect 10649 4511 10701 4563
rect 10780 4332 10832 4384
rect 10951 4406 11003 4415
rect 10951 4288 10960 4406
rect 10960 4288 10994 4406
rect 10994 4288 11003 4406
rect 10951 4279 11003 4288
rect 10649 4155 10701 4207
rect 10780 3976 10832 4028
rect 10649 3799 10701 3851
rect 10545 3676 10597 3728
rect 10780 3620 10832 3672
rect 10551 3556 10603 3608
rect 10651 3442 10703 3494
rect 108 3288 160 3297
rect 1766 3288 1818 3297
rect 5082 3288 5134 3297
rect 8398 3288 8450 3297
rect 10056 3288 10108 3297
rect 108 3254 117 3288
rect 117 3254 160 3288
rect 1766 3254 1818 3288
rect 5082 3254 5134 3288
rect 8398 3254 8450 3288
rect 10056 3254 10099 3288
rect 10099 3254 10108 3288
rect 108 3245 160 3254
rect 1766 3245 1818 3254
rect 5082 3245 5134 3254
rect 8398 3245 8450 3254
rect 10056 3245 10108 3254
rect 10780 3264 10832 3316
rect 1462 2549 1514 2558
rect 5236 2549 5288 2558
rect 8702 2549 8754 2558
rect 1462 2515 1514 2549
rect 5236 2515 5288 2549
rect 8702 2515 8754 2549
rect 1462 2506 1514 2515
rect 5236 2506 5288 2515
rect 8702 2506 8754 2515
rect 108 2112 160 2121
rect 3424 2112 3476 2121
rect 6740 2112 6792 2121
rect 10056 2112 10108 2121
rect 108 2078 160 2112
rect 3424 2078 3476 2112
rect 6740 2078 6792 2112
rect 10056 2078 10108 2112
rect 108 2069 160 2078
rect 3424 2069 3476 2078
rect 6740 2069 6792 2078
rect 10056 2069 10108 2078
rect 353 1931 405 1983
rect 3144 1931 3196 1983
rect 4731 1931 4783 1983
rect 6963 1931 7015 1983
rect 9860 1931 9912 1983
rect 108 1714 160 1766
rect 1766 1714 1818 1766
rect 3424 1714 3476 1766
rect 5082 1714 5134 1766
rect 6740 1714 6792 1766
rect 8398 1714 8450 1766
rect 10056 1714 10108 1766
rect 353 1621 405 1673
rect 3144 1621 3196 1673
rect 4731 1621 4783 1673
rect 6963 1621 7015 1673
rect 9860 1621 9912 1673
rect 353 1513 405 1565
rect 3144 1513 3196 1565
rect 4731 1513 4783 1565
rect 6963 1513 7015 1565
rect 9860 1513 9912 1565
rect 108 1296 160 1348
rect 1766 1296 1818 1348
rect 3424 1296 3476 1348
rect 5082 1296 5134 1348
rect 6740 1296 6792 1348
rect 8398 1296 8450 1348
rect 10056 1296 10108 1348
rect 353 1203 405 1255
rect 3144 1203 3196 1255
rect 4731 1203 4783 1255
rect 6963 1203 7015 1255
rect 9860 1203 9912 1255
rect 353 1095 405 1147
rect 3144 1095 3196 1147
rect 4731 1095 4783 1147
rect 6963 1095 7015 1147
rect 9860 1095 9912 1147
rect 108 878 160 930
rect 1766 878 1818 930
rect 3424 878 3476 930
rect 5082 878 5134 930
rect 6740 878 6792 930
rect 8398 878 8450 930
rect 10056 878 10108 930
rect 353 785 405 837
rect 3144 785 3196 837
rect 4731 785 4783 837
rect 6963 785 7015 837
rect 9860 785 9912 837
rect 353 677 405 729
rect 3144 677 3196 729
rect 4731 677 4783 729
rect 6963 677 7015 729
rect 9860 677 9912 729
rect 108 460 160 512
rect 1766 460 1818 512
rect 3424 460 3476 512
rect 5082 460 5134 512
rect 6740 460 6792 512
rect 8398 460 8450 512
rect 10056 460 10108 512
rect 353 367 405 419
rect 3144 367 3196 419
rect 4731 367 4783 419
rect 6963 367 7015 419
rect 9860 367 9912 419
rect 353 259 405 311
rect 3144 259 3196 311
rect 4731 259 4783 311
rect 6963 259 7015 311
rect 9860 259 9912 311
rect 108 42 160 94
rect 1766 42 1818 94
rect 3424 42 3476 94
rect 5082 42 5134 94
rect 6740 42 6792 94
rect 8398 42 8450 94
rect 10056 42 10108 94
rect 353 -51 405 1
rect 3144 -51 3196 1
rect 4731 -51 4783 1
rect 6963 -51 7015 1
rect 9860 -51 9912 1
rect 353 -159 405 -107
rect 3144 -159 3196 -107
rect 4731 -159 4783 -107
rect 6963 -159 7015 -107
rect 9860 -159 9912 -107
rect 108 -376 160 -324
rect 1766 -376 1818 -324
rect 3424 -376 3476 -324
rect 5082 -376 5134 -324
rect 6740 -376 6792 -324
rect 8398 -376 8450 -324
rect 10056 -376 10108 -324
rect 353 -469 405 -417
rect 3144 -469 3196 -417
rect 4731 -469 4783 -417
rect 6963 -469 7015 -417
rect 9860 -469 9912 -417
rect 353 -577 405 -525
rect 3144 -577 3196 -525
rect 4731 -577 4783 -525
rect 6963 -577 7015 -525
rect 9860 -577 9912 -525
rect 108 -794 160 -742
rect 1766 -794 1818 -742
rect 3424 -794 3476 -742
rect 5082 -794 5134 -742
rect 6740 -794 6792 -742
rect 8398 -794 8450 -742
rect 10056 -794 10108 -742
rect 353 -887 405 -835
rect 3144 -887 3196 -835
rect 4731 -887 4783 -835
rect 6963 -887 7015 -835
rect 9860 -887 9912 -835
rect 353 -995 405 -943
rect 3144 -995 3196 -943
rect 4731 -995 4783 -943
rect 6963 -995 7015 -943
rect 9860 -995 9912 -943
rect 108 -1212 160 -1160
rect 1766 -1212 1818 -1160
rect 3424 -1212 3476 -1160
rect 5082 -1212 5134 -1160
rect 6740 -1212 6792 -1160
rect 8398 -1212 8450 -1160
rect 10056 -1212 10108 -1160
rect 353 -1305 405 -1253
rect 3144 -1305 3196 -1253
rect 4731 -1305 4783 -1253
rect 6963 -1305 7015 -1253
rect 9860 -1305 9912 -1253
rect 108 -1400 160 -1391
rect 3424 -1400 3476 -1391
rect 6740 -1400 6792 -1391
rect 10056 -1400 10108 -1391
rect 108 -1434 160 -1400
rect 3424 -1434 3476 -1400
rect 6740 -1434 6792 -1400
rect 10056 -1434 10108 -1400
rect 108 -1443 160 -1434
rect 3424 -1443 3476 -1434
rect 6740 -1443 6792 -1434
rect 10056 -1443 10108 -1434
rect 1462 -2026 1514 -2017
rect 5236 -2026 5288 -2017
rect 8702 -2026 8754 -2017
rect 1462 -2060 1514 -2026
rect 5236 -2060 5288 -2026
rect 8702 -2060 8754 -2026
rect 1462 -2069 1514 -2060
rect 5236 -2069 5288 -2060
rect 8702 -2069 8754 -2060
<< metal2 >>
rect -619 9746 -545 9755
rect -619 9616 -610 9746
rect -554 9616 -545 9746
rect -619 9607 -545 9616
rect 97 9746 171 9755
rect 97 9616 106 9746
rect 162 9616 171 9746
rect 97 9607 171 9616
rect 1755 9746 1829 9755
rect 1755 9616 1764 9746
rect 1820 9616 1829 9746
rect 1755 9607 1829 9616
rect 5071 9746 5145 9755
rect 5071 9616 5080 9746
rect 5136 9616 5145 9746
rect 5071 9607 5145 9616
rect 8387 9746 8461 9755
rect 8387 9616 8396 9746
rect 8452 9616 8461 9746
rect 8387 9607 8461 9616
rect 10045 9746 10119 9755
rect 10045 9616 10054 9746
rect 10110 9616 10119 9746
rect 10045 9607 10119 9616
rect 10734 9746 10808 9755
rect 10734 9616 10743 9746
rect 10799 9616 10808 9746
rect 10734 9607 10808 9616
rect -614 7223 -550 9607
rect 102 9163 166 9607
rect 102 9111 108 9163
rect 160 9111 166 9163
rect 102 8798 166 9111
rect 102 8746 108 8798
rect 160 8746 166 8798
rect 102 8433 166 8746
rect 102 8381 108 8433
rect 160 8381 166 8433
rect 102 8068 166 8381
rect 102 8016 108 8068
rect 160 8016 166 8068
rect 102 7534 166 8016
rect 102 7482 108 7534
rect 160 7482 166 7534
rect -614 7171 -608 7223
rect -556 7171 -550 7223
rect -614 6858 -550 7171
rect -361 7225 -287 7234
rect -361 7169 -352 7225
rect -296 7169 -287 7225
rect -361 7160 -287 7169
rect 102 7169 166 7482
rect -614 6806 -608 6858
rect -556 6806 -550 6858
rect -614 6493 -550 6806
rect -614 6441 -608 6493
rect -556 6441 -550 6493
rect -614 6435 -550 6441
rect -485 7115 -421 7121
rect -485 7063 -479 7115
rect -427 7063 -421 7115
rect -485 6750 -421 7063
rect 102 7117 108 7169
rect 160 7117 166 7169
rect -361 6860 -287 6869
rect -361 6804 -352 6860
rect -296 6804 -287 6860
rect -361 6795 -287 6804
rect 102 6804 166 7117
rect -485 6698 -479 6750
rect -427 6698 -421 6750
rect -485 6385 -421 6698
rect 102 6752 108 6804
rect 160 6752 166 6804
rect -356 6481 -141 6487
rect -356 6429 -350 6481
rect -298 6429 -141 6481
rect -356 6423 -141 6429
rect -485 6369 -479 6385
rect -765 6333 -479 6369
rect -427 6333 -421 6385
rect -765 6305 -421 6333
rect -765 4757 -701 6305
rect -205 6246 -141 6423
rect -485 6182 -141 6246
rect -614 6116 -550 6122
rect -614 6064 -608 6116
rect -556 6064 -550 6116
rect -614 5359 -550 6064
rect -485 6020 -421 6182
rect -485 5968 -479 6020
rect -427 5968 -421 6020
rect -485 5962 -421 5968
rect -356 6116 -292 6122
rect -356 6064 -350 6116
rect -298 6064 -292 6116
rect -624 5350 -550 5359
rect -624 5349 -615 5350
rect -644 5294 -615 5349
rect -559 5294 -550 5350
rect -356 5349 -292 6064
rect -644 5285 -550 5294
rect -386 5285 -292 5349
rect -644 5020 -580 5285
rect -644 4968 -638 5020
rect -586 4968 -580 5020
rect -644 4962 -580 4968
rect -515 5107 -451 5113
rect -515 5055 -509 5107
rect -457 5055 -451 5107
rect -515 4757 -451 5055
rect -386 5031 -322 5285
rect -391 5022 -317 5031
rect -391 4966 -382 5022
rect -326 4966 -317 5022
rect -391 4957 -317 4966
rect -205 4877 -141 6182
rect 102 6439 166 6752
rect 102 6387 108 6439
rect 160 6387 166 6439
rect 102 6074 166 6387
rect 102 6022 108 6074
rect 160 6022 166 6074
rect 102 5709 166 6022
rect 102 5657 108 5709
rect 160 5657 166 5709
rect 102 5344 166 5657
rect 102 5292 108 5344
rect 160 5292 166 5344
rect 102 5100 166 5292
rect 102 5048 108 5100
rect 160 5048 166 5100
rect -107 5015 -33 5024
rect -107 4959 -98 5015
rect -42 4959 -33 5015
rect -107 4950 -33 4959
rect -765 4751 -451 4757
rect -765 4699 -561 4751
rect -509 4699 -451 4751
rect -765 4693 -451 4699
rect -322 4813 -141 4877
rect -322 4670 -258 4813
rect -386 4664 -258 4670
rect -386 4612 -380 4664
rect -328 4612 -258 4664
rect -386 4606 -258 4612
rect -644 4528 -580 4534
rect -644 4476 -638 4528
rect -586 4476 -580 4528
rect -644 4347 -580 4476
rect -386 4445 -322 4606
rect -515 4395 -322 4445
rect -649 4338 -575 4347
rect -649 4282 -640 4338
rect -584 4282 -575 4338
rect -649 4273 -575 4282
rect -515 4343 -509 4395
rect -457 4381 -322 4395
rect -457 4343 -451 4381
rect -644 4172 -580 4273
rect -644 4120 -638 4172
rect -586 4120 -580 4172
rect -644 3816 -580 4120
rect -644 3764 -638 3816
rect -586 3764 -580 3816
rect -644 3460 -580 3764
rect -515 4039 -451 4343
rect -393 4184 -319 4193
rect -100 4187 -40 4950
rect 102 4937 166 5048
rect 102 4885 108 4937
rect 160 4885 166 4937
rect 102 4566 166 4885
rect 102 4514 108 4566
rect 160 4514 166 4566
rect 102 4508 166 4514
rect 1760 9163 1824 9607
rect 1760 9111 1766 9163
rect 1818 9111 1824 9163
rect 1760 8798 1824 9111
rect 1760 8746 1766 8798
rect 1818 8746 1824 8798
rect 1760 8433 1824 8746
rect 1760 8381 1766 8433
rect 1818 8381 1824 8433
rect 1760 8068 1824 8381
rect 1760 8016 1766 8068
rect 1818 8016 1824 8068
rect 1760 7534 1824 8016
rect 1760 7482 1766 7534
rect 1818 7482 1824 7534
rect 1760 7169 1824 7482
rect 1760 7117 1766 7169
rect 1818 7117 1824 7169
rect 1760 6804 1824 7117
rect 1760 6752 1766 6804
rect 1818 6752 1824 6804
rect 1760 6439 1824 6752
rect 1760 6387 1766 6439
rect 1818 6387 1824 6439
rect 1760 6074 1824 6387
rect 1760 6022 1766 6074
rect 1818 6022 1824 6074
rect 1760 5709 1824 6022
rect 1760 5657 1766 5709
rect 1818 5657 1824 5709
rect 1760 5344 1824 5657
rect 1760 5292 1766 5344
rect 1818 5292 1824 5344
rect 1760 5100 1824 5292
rect 1760 5048 1766 5100
rect 1818 5048 1824 5100
rect 1760 4937 1824 5048
rect 3418 9162 3482 9295
rect 3418 9110 3424 9162
rect 3476 9110 3482 9162
rect 3418 8797 3482 9110
rect 3418 8745 3424 8797
rect 3476 8745 3482 8797
rect 3418 8432 3482 8745
rect 3418 8380 3424 8432
rect 3476 8380 3482 8432
rect 3418 8068 3482 8380
rect 3418 8016 3424 8068
rect 3476 8016 3482 8068
rect 3418 7534 3482 8016
rect 5076 9163 5140 9607
rect 5076 9111 5082 9163
rect 5134 9111 5140 9163
rect 5076 8798 5140 9111
rect 5076 8746 5082 8798
rect 5134 8746 5140 8798
rect 5076 8433 5140 8746
rect 5076 8381 5082 8433
rect 5134 8381 5140 8433
rect 5076 8068 5140 8381
rect 5076 8016 5082 8068
rect 5134 8016 5140 8068
rect 3418 7482 3424 7534
rect 3476 7482 3482 7534
rect 3418 7223 3482 7482
rect 3418 7167 3422 7223
rect 3478 7167 3482 7223
rect 3418 7117 3424 7167
rect 3476 7117 3482 7167
rect 3418 6804 3482 7117
rect 3418 6752 3424 6804
rect 3476 6752 3482 6804
rect 3418 6439 3482 6752
rect 3418 6387 3424 6439
rect 3476 6387 3482 6439
rect 3418 6074 3482 6387
rect 3418 6022 3424 6074
rect 3476 6022 3482 6074
rect 3418 5709 3482 6022
rect 3418 5657 3424 5709
rect 3476 5657 3482 5709
rect 3418 5344 3482 5657
rect 3418 5292 3424 5344
rect 3476 5292 3482 5344
rect 3418 5075 3482 5292
rect 4300 7428 4364 7596
rect 4300 7376 4306 7428
rect 4358 7376 4364 7428
rect 4300 7063 4364 7376
rect 4300 7011 4306 7063
rect 4358 7011 4364 7063
rect 4300 6698 4364 7011
rect 4300 6646 4306 6698
rect 4358 6646 4364 6698
rect 4300 6333 4364 6646
rect 4300 6281 4306 6333
rect 4358 6281 4364 6333
rect 4300 5968 4364 6281
rect 4300 5916 4306 5968
rect 4358 5916 4364 5968
rect 4300 5603 4364 5916
rect 4300 5551 4306 5603
rect 4358 5551 4364 5603
rect 4300 5238 4364 5551
rect 4300 5186 4306 5238
rect 4358 5186 4364 5238
rect 3418 5011 3678 5075
rect 1760 4885 1766 4937
rect 1818 4885 1824 4937
rect 1760 4566 1824 4885
rect 3418 4807 3482 4813
rect 3418 4755 3424 4807
rect 3476 4755 3482 4807
rect 3418 4749 3482 4755
rect 1760 4514 1766 4566
rect 1818 4514 1824 4566
rect 97 4409 171 4420
rect 1760 4415 1824 4514
rect 97 4281 106 4409
rect 162 4281 171 4409
rect 97 4272 171 4281
rect 1456 4351 1824 4415
rect -393 4128 -384 4184
rect -328 4128 -319 4184
rect -393 4119 -319 4128
rect -109 4178 -35 4187
rect -109 4122 -100 4178
rect -44 4122 -35 4178
rect -109 4113 -35 4122
rect 102 4177 166 4272
rect 102 4125 108 4177
rect 160 4125 166 4177
rect -515 3987 -509 4039
rect -457 3987 -451 4039
rect -515 3683 -451 3987
rect -395 3952 -321 3960
rect -395 3951 -380 3952
rect -395 3895 -386 3951
rect -328 3900 -321 3952
rect -330 3895 -321 3900
rect -395 3886 -321 3895
rect -515 3631 -509 3683
rect -457 3631 -451 3683
rect -515 3625 -451 3631
rect -100 3603 -40 4113
rect 102 3946 166 4125
rect 102 3894 108 3946
rect 160 3894 166 3946
rect -395 3596 -321 3603
rect -395 3594 -380 3596
rect -395 3538 -386 3594
rect -327 3544 -321 3596
rect -330 3538 -321 3544
rect -395 3529 -321 3538
rect -109 3594 -35 3603
rect -109 3538 -100 3594
rect -44 3538 -35 3594
rect -109 3529 -35 3538
rect 102 3590 166 3894
rect 102 3538 108 3590
rect 160 3538 166 3590
rect -644 3408 -638 3460
rect -586 3408 -580 3460
rect -644 3402 -580 3408
rect 102 3297 166 3538
rect 102 3245 108 3297
rect 160 3245 166 3297
rect 102 2251 166 3245
rect 1456 2558 1520 4351
rect 1760 4177 1824 4183
rect 1760 4125 1766 4177
rect 1818 4125 1824 4177
rect 1760 3946 1824 4125
rect 3424 3953 3476 4749
rect 1760 3894 1766 3946
rect 1818 3894 1824 3946
rect 1760 3590 1824 3894
rect 3409 3946 3483 3953
rect 3409 3944 3424 3946
rect 3409 3888 3418 3944
rect 3476 3894 3483 3946
rect 3474 3888 3483 3894
rect 3409 3879 3483 3888
rect 1760 3538 1766 3590
rect 1818 3538 1824 3590
rect 1760 3297 1824 3538
rect 3409 3590 3483 3597
rect 3409 3588 3424 3590
rect 3409 3532 3418 3588
rect 3476 3538 3483 3590
rect 3474 3532 3483 3538
rect 3409 3523 3483 3532
rect 1760 3245 1766 3297
rect 1818 3245 1824 3297
rect 1760 3239 1824 3245
rect 3133 2915 3207 2924
rect 3133 2859 3142 2915
rect 3198 2859 3207 2915
rect 3133 2850 3207 2859
rect 1456 2506 1462 2558
rect 1514 2506 1520 2558
rect 102 2187 411 2251
rect 102 2184 166 2187
rect 102 2121 166 2124
rect 102 2069 108 2121
rect 160 2069 166 2121
rect 102 1766 166 2069
rect 102 1714 108 1766
rect 160 1714 166 1766
rect 102 1348 166 1714
rect 102 1296 108 1348
rect 160 1296 166 1348
rect 102 930 166 1296
rect 102 878 108 930
rect 160 878 166 930
rect 102 512 166 878
rect 102 460 108 512
rect 160 460 166 512
rect 102 94 166 460
rect 102 42 108 94
rect 160 42 166 94
rect 102 -324 166 42
rect 102 -376 108 -324
rect 160 -376 166 -324
rect 102 -742 166 -376
rect 102 -794 108 -742
rect 160 -794 166 -742
rect 102 -1160 166 -794
rect 102 -1212 108 -1160
rect 160 -1212 166 -1160
rect 102 -1391 166 -1212
rect 102 -1443 108 -1391
rect 160 -1443 166 -1391
rect 102 -1446 166 -1443
rect 347 1983 411 2187
rect 347 1931 353 1983
rect 405 1931 411 1983
rect 347 1673 411 1931
rect 347 1621 353 1673
rect 405 1621 411 1673
rect 347 1565 411 1621
rect 347 1513 353 1565
rect 405 1513 411 1565
rect 347 1255 411 1513
rect 347 1203 353 1255
rect 405 1203 411 1255
rect 347 1147 411 1203
rect 347 1095 353 1147
rect 405 1095 411 1147
rect 347 837 411 1095
rect 347 785 353 837
rect 405 785 411 837
rect 347 729 411 785
rect 347 677 353 729
rect 405 677 411 729
rect 347 419 411 677
rect 347 367 353 419
rect 405 367 411 419
rect 347 311 411 367
rect 347 259 353 311
rect 405 259 411 311
rect 347 1 411 259
rect 347 -51 353 1
rect 405 -51 411 1
rect 347 -107 411 -51
rect 347 -159 353 -107
rect 405 -159 411 -107
rect 347 -417 411 -159
rect 347 -469 353 -417
rect 405 -469 411 -417
rect 347 -525 411 -469
rect 347 -577 353 -525
rect 405 -577 411 -525
rect 347 -835 411 -577
rect 347 -887 353 -835
rect 405 -887 411 -835
rect 347 -943 411 -887
rect 347 -995 353 -943
rect 405 -995 411 -943
rect 347 -1253 411 -995
rect 347 -1305 353 -1253
rect 405 -1305 411 -1253
rect 347 -1676 411 -1305
rect 345 -1685 419 -1676
rect 345 -1815 354 -1685
rect 410 -1815 419 -1685
rect 345 -1824 419 -1815
rect 1456 -2017 1520 2506
rect 1755 2315 1829 2324
rect 1755 2259 1764 2315
rect 1820 2259 1829 2315
rect 1755 2250 1829 2259
rect 1766 1772 1818 2250
rect 3144 1983 3196 2850
rect 3614 2724 3678 5011
rect 4300 4705 4364 5186
rect 4300 4653 4306 4705
rect 4358 4653 4364 4705
rect 3609 2715 3683 2724
rect 3609 2659 3618 2715
rect 3674 2659 3683 2715
rect 3609 2650 3683 2659
rect 3413 2515 3487 2524
rect 3413 2459 3422 2515
rect 3478 2459 3487 2515
rect 3413 2450 3487 2459
rect 1760 1766 1824 1772
rect 1760 1714 1766 1766
rect 1818 1714 1824 1766
rect 1760 1708 1824 1714
rect 1766 1354 1818 1708
rect 3144 1673 3196 1931
rect 3424 2121 3476 2450
rect 4300 2324 4364 4653
rect 5076 7534 5140 8016
rect 6734 9255 6795 9295
rect 6734 9163 6798 9255
rect 6734 9111 6740 9163
rect 6792 9111 6798 9163
rect 6734 9022 6798 9111
rect 8392 9163 8456 9607
rect 8392 9111 8398 9163
rect 8450 9111 8456 9163
rect 6734 8890 6795 9022
rect 6734 8798 6798 8890
rect 6734 8746 6740 8798
rect 6792 8746 6798 8798
rect 6734 8657 6798 8746
rect 8392 8798 8456 9111
rect 8392 8746 8398 8798
rect 8450 8746 8456 8798
rect 6734 8525 6795 8657
rect 6734 8433 6798 8525
rect 6734 8381 6740 8433
rect 6792 8381 6798 8433
rect 6734 8292 6798 8381
rect 8392 8433 8456 8746
rect 8392 8381 8398 8433
rect 8450 8381 8456 8433
rect 6734 8160 6795 8292
rect 6734 8068 6798 8160
rect 6734 8016 6740 8068
rect 6792 8016 6798 8068
rect 6734 7927 6798 8016
rect 6736 7596 6798 7927
rect 5076 7482 5082 7534
rect 5134 7482 5140 7534
rect 5076 7169 5140 7482
rect 5076 7117 5082 7169
rect 5134 7117 5140 7169
rect 5076 6804 5140 7117
rect 5076 6752 5082 6804
rect 5134 6752 5140 6804
rect 5076 6439 5140 6752
rect 5076 6387 5082 6439
rect 5134 6387 5140 6439
rect 5076 6074 5140 6387
rect 5076 6022 5082 6074
rect 5134 6022 5140 6074
rect 5076 5709 5140 6022
rect 5076 5657 5082 5709
rect 5134 5657 5140 5709
rect 5076 5344 5140 5657
rect 5076 5292 5082 5344
rect 5134 5292 5140 5344
rect 5076 5100 5140 5292
rect 5076 5048 5082 5100
rect 5134 5048 5140 5100
rect 5076 4937 5140 5048
rect 5076 4885 5082 4937
rect 5134 4885 5140 4937
rect 5076 4572 5140 4885
rect 5956 7428 6020 7596
rect 5956 7376 5962 7428
rect 6014 7376 6020 7428
rect 5956 7063 6020 7376
rect 5956 7011 5962 7063
rect 6014 7011 6020 7063
rect 5956 6698 6020 7011
rect 5956 6646 5962 6698
rect 6014 6646 6020 6698
rect 5956 6333 6020 6646
rect 5956 6281 5962 6333
rect 6014 6281 6020 6333
rect 5956 5968 6020 6281
rect 5956 5916 5962 5968
rect 6014 5916 6020 5968
rect 5956 5603 6020 5916
rect 5956 5551 5962 5603
rect 6014 5551 6020 5603
rect 5956 5238 6020 5551
rect 5956 5186 5962 5238
rect 6014 5186 6020 5238
rect 5956 4705 6020 5186
rect 6734 7534 6798 7596
rect 6734 7482 6740 7534
rect 6792 7482 6798 7534
rect 6734 7169 6798 7482
rect 6734 7117 6740 7169
rect 6792 7117 6798 7169
rect 6734 6859 6798 7117
rect 6734 6752 6740 6859
rect 6796 6803 6798 6859
rect 6792 6752 6798 6803
rect 6734 6439 6798 6752
rect 6734 6387 6740 6439
rect 6792 6387 6798 6439
rect 6734 6074 6798 6387
rect 6734 6022 6740 6074
rect 6792 6022 6798 6074
rect 6734 5709 6798 6022
rect 6734 5657 6740 5709
rect 6792 5657 6798 5709
rect 6734 5344 6798 5657
rect 6734 5292 6740 5344
rect 6792 5292 6798 5344
rect 6734 5075 6798 5292
rect 5956 4653 5962 4705
rect 6014 4653 6020 4705
rect 5076 4566 5294 4572
rect 5076 4514 5082 4566
rect 5134 4514 5294 4566
rect 5076 4508 5294 4514
rect 5071 4410 5145 4421
rect 5071 4282 5080 4410
rect 5136 4282 5145 4410
rect 5071 4273 5145 4282
rect 5076 4177 5140 4273
rect 5076 4125 5082 4177
rect 5134 4125 5140 4177
rect 5076 3946 5140 4125
rect 5076 3894 5082 3946
rect 5134 3894 5140 3946
rect 5076 3590 5140 3894
rect 5076 3538 5082 3590
rect 5134 3538 5140 3590
rect 5076 3297 5140 3538
rect 5076 3245 5082 3297
rect 5134 3245 5140 3297
rect 5076 3239 5140 3245
rect 4720 3115 4794 3124
rect 4720 3059 4729 3115
rect 4785 3059 4794 3115
rect 4720 3050 4794 3059
rect 4295 2315 4369 2324
rect 4295 2259 4304 2315
rect 4360 2259 4369 2315
rect 4295 2250 4369 2259
rect 3424 1772 3476 2069
rect 4731 1983 4783 3050
rect 5071 2715 5145 2724
rect 5071 2659 5080 2715
rect 5136 2659 5145 2715
rect 5071 2650 5145 2659
rect 3418 1766 3482 1772
rect 3418 1714 3424 1766
rect 3476 1714 3482 1766
rect 3418 1708 3482 1714
rect 3144 1565 3196 1621
rect 1760 1348 1824 1354
rect 1760 1296 1766 1348
rect 1818 1296 1824 1348
rect 1760 1290 1824 1296
rect 1766 936 1818 1290
rect 3144 1255 3196 1513
rect 3424 1354 3476 1708
rect 4731 1673 4783 1931
rect 5082 1772 5134 2650
rect 5230 2558 5294 4508
rect 5956 2721 6020 4653
rect 6538 5011 6798 5075
rect 8392 8068 8456 8381
rect 8392 8016 8398 8068
rect 8450 8016 8456 8068
rect 8392 7534 8456 8016
rect 8392 7482 8398 7534
rect 8450 7482 8456 7534
rect 8392 7169 8456 7482
rect 8392 7117 8398 7169
rect 8450 7117 8456 7169
rect 8392 6804 8456 7117
rect 8392 6752 8398 6804
rect 8450 6752 8456 6804
rect 8392 6439 8456 6752
rect 8392 6387 8398 6439
rect 8450 6387 8456 6439
rect 8392 6074 8456 6387
rect 8392 6022 8398 6074
rect 8450 6022 8456 6074
rect 8392 5709 8456 6022
rect 8392 5657 8398 5709
rect 8450 5657 8456 5709
rect 8392 5344 8456 5657
rect 8392 5292 8398 5344
rect 8450 5292 8456 5344
rect 8392 5100 8456 5292
rect 8392 5048 8398 5100
rect 8450 5048 8456 5100
rect 5950 2712 6024 2721
rect 5950 2656 5959 2712
rect 6015 2656 6024 2712
rect 5950 2647 6024 2656
rect 5230 2506 5236 2558
rect 5288 2506 5294 2558
rect 5076 1766 5140 1772
rect 5076 1714 5082 1766
rect 5134 1714 5140 1766
rect 5076 1708 5140 1714
rect 4731 1565 4783 1621
rect 3418 1348 3482 1354
rect 3418 1296 3424 1348
rect 3476 1296 3482 1348
rect 3418 1290 3482 1296
rect 3144 1147 3196 1203
rect 1760 930 1824 936
rect 1760 878 1766 930
rect 1818 878 1824 930
rect 1760 872 1824 878
rect 1766 518 1818 872
rect 3144 837 3196 1095
rect 3424 936 3476 1290
rect 4731 1255 4783 1513
rect 5082 1354 5134 1708
rect 5076 1348 5140 1354
rect 5076 1296 5082 1348
rect 5134 1296 5140 1348
rect 5076 1290 5140 1296
rect 4731 1147 4783 1203
rect 3418 930 3482 936
rect 3418 878 3424 930
rect 3476 878 3482 930
rect 3418 872 3482 878
rect 3144 729 3196 785
rect 1760 512 1824 518
rect 1760 460 1766 512
rect 1818 460 1824 512
rect 1760 454 1824 460
rect 1766 100 1818 454
rect 3144 419 3196 677
rect 3424 518 3476 872
rect 4731 837 4783 1095
rect 5082 936 5134 1290
rect 5076 930 5140 936
rect 5076 878 5082 930
rect 5134 878 5140 930
rect 5076 872 5140 878
rect 4731 729 4783 785
rect 3418 512 3482 518
rect 3418 460 3424 512
rect 3476 460 3482 512
rect 3418 454 3482 460
rect 3144 311 3196 367
rect 1760 94 1824 100
rect 1760 42 1766 94
rect 1818 42 1824 94
rect 1760 36 1824 42
rect 1766 -318 1818 36
rect 3144 1 3196 259
rect 3424 100 3476 454
rect 4731 419 4783 677
rect 5082 518 5134 872
rect 5076 512 5140 518
rect 5076 460 5082 512
rect 5134 460 5140 512
rect 5076 454 5140 460
rect 4731 311 4783 367
rect 3418 94 3482 100
rect 3418 42 3424 94
rect 3476 42 3482 94
rect 3418 36 3482 42
rect 3144 -107 3196 -51
rect 1760 -324 1824 -318
rect 1760 -376 1766 -324
rect 1818 -376 1824 -324
rect 1760 -382 1824 -376
rect 1766 -736 1818 -382
rect 3144 -417 3196 -159
rect 3424 -318 3476 36
rect 4731 1 4783 259
rect 5082 100 5134 454
rect 5076 94 5140 100
rect 5076 42 5082 94
rect 5134 42 5140 94
rect 5076 36 5140 42
rect 4731 -107 4783 -51
rect 3418 -324 3482 -318
rect 3418 -376 3424 -324
rect 3476 -376 3482 -324
rect 3418 -382 3482 -376
rect 3144 -525 3196 -469
rect 1760 -742 1824 -736
rect 1760 -794 1766 -742
rect 1818 -794 1824 -742
rect 1760 -800 1824 -794
rect 1766 -1154 1818 -800
rect 3144 -835 3196 -577
rect 3424 -736 3476 -382
rect 4731 -417 4783 -159
rect 5082 -318 5134 36
rect 5076 -324 5140 -318
rect 5076 -376 5082 -324
rect 5134 -376 5140 -324
rect 5076 -382 5140 -376
rect 4731 -525 4783 -469
rect 3418 -742 3482 -736
rect 3418 -794 3424 -742
rect 3476 -794 3482 -742
rect 3418 -800 3482 -794
rect 3144 -943 3196 -887
rect 1760 -1160 1824 -1154
rect 1760 -1212 1766 -1160
rect 1818 -1212 1824 -1160
rect 1760 -1218 1824 -1212
rect 1766 -1224 1818 -1218
rect 3144 -1253 3196 -995
rect 3424 -1154 3476 -800
rect 4731 -835 4783 -577
rect 5082 -736 5134 -382
rect 5076 -742 5140 -736
rect 5076 -794 5082 -742
rect 5134 -794 5140 -742
rect 5076 -800 5140 -794
rect 4731 -943 4783 -887
rect 3418 -1160 3482 -1154
rect 3418 -1212 3424 -1160
rect 3476 -1212 3482 -1160
rect 3418 -1218 3482 -1212
rect 3144 -1311 3196 -1305
rect 3424 -1391 3476 -1218
rect 4731 -1253 4783 -995
rect 5082 -1154 5134 -800
rect 5076 -1160 5140 -1154
rect 5076 -1212 5082 -1160
rect 5134 -1212 5140 -1160
rect 5076 -1218 5140 -1212
rect 5082 -1224 5134 -1218
rect 4731 -1311 4783 -1305
rect 3424 -1449 3476 -1443
rect 1456 -2069 1462 -2017
rect 1514 -2069 1520 -2017
rect 1456 -2075 1520 -2069
rect 5230 -2017 5294 2506
rect 6538 2324 6602 5011
rect 8392 4937 8456 5048
rect 8392 4885 8398 4937
rect 8450 4885 8456 4937
rect 6734 4807 6798 4813
rect 6734 4755 6740 4807
rect 6792 4755 6798 4807
rect 6734 4749 6798 4755
rect 6740 3954 6792 4749
rect 8392 4415 8456 4885
rect 10050 9163 10114 9607
rect 10050 9111 10056 9163
rect 10108 9111 10114 9163
rect 10050 8798 10114 9111
rect 10050 8746 10056 8798
rect 10108 8746 10114 8798
rect 10050 8433 10114 8746
rect 10050 8381 10056 8433
rect 10108 8381 10114 8433
rect 10050 8068 10114 8381
rect 10050 8016 10056 8068
rect 10108 8016 10114 8068
rect 10050 7534 10114 8016
rect 10050 7482 10056 7534
rect 10108 7482 10114 7534
rect 10050 7169 10114 7482
rect 10739 7510 10803 9607
rect 10739 7458 10745 7510
rect 10797 7458 10803 7510
rect 10739 7376 10803 7458
rect 10739 7324 10745 7376
rect 10797 7324 10803 7376
rect 10050 7117 10056 7169
rect 10108 7117 10114 7169
rect 10050 6804 10114 7117
rect 10050 6752 10056 6804
rect 10108 6752 10114 6804
rect 10050 6439 10114 6752
rect 10050 6387 10056 6439
rect 10108 6387 10114 6439
rect 10050 6074 10114 6387
rect 10609 7198 10673 7204
rect 10609 7146 10615 7198
rect 10667 7146 10673 7198
rect 10609 6842 10673 7146
rect 10609 6790 10615 6842
rect 10667 6790 10673 6842
rect 10609 6486 10673 6790
rect 10609 6434 10615 6486
rect 10667 6434 10673 6486
rect 10609 6142 10673 6434
rect 10739 7020 10803 7324
rect 10739 6968 10745 7020
rect 10797 6968 10803 7020
rect 10739 6664 10803 6968
rect 10739 6612 10745 6664
rect 10797 6612 10803 6664
rect 10739 6308 10803 6612
rect 10739 6256 10745 6308
rect 10797 6256 10803 6308
rect 10050 6022 10056 6074
rect 10108 6022 10114 6074
rect 10050 5709 10114 6022
rect 10050 5657 10056 5709
rect 10108 5657 10114 5709
rect 10050 5344 10114 5657
rect 10050 5292 10056 5344
rect 10108 5292 10114 5344
rect 10050 5100 10114 5292
rect 10050 5048 10056 5100
rect 10108 5048 10114 5100
rect 10050 4937 10114 5048
rect 10050 4885 10056 4937
rect 10108 4885 10114 4937
rect 10186 6130 10260 6139
rect 10186 6074 10195 6130
rect 10251 6074 10260 6130
rect 10186 6065 10260 6074
rect 10602 6133 10676 6142
rect 10602 6077 10611 6133
rect 10667 6077 10676 6133
rect 10602 6068 10676 6077
rect 10186 4922 10242 6065
rect 10506 6007 10570 6013
rect 10506 5955 10512 6007
rect 10564 5995 10570 6007
rect 10564 5955 10665 5995
rect 10506 5949 10665 5955
rect 10609 5780 10665 5949
rect 10739 5952 10803 6256
rect 10739 5900 10745 5952
rect 10797 5900 10803 5952
rect 10609 5774 10673 5780
rect 10609 5722 10615 5774
rect 10667 5722 10673 5774
rect 10609 5716 10673 5722
rect 10508 5661 10572 5667
rect 10508 5656 10514 5661
rect 10312 5609 10514 5656
rect 10566 5609 10572 5661
rect 10312 5603 10572 5609
rect 10050 4566 10114 4885
rect 10174 4913 10248 4922
rect 10174 4857 10183 4913
rect 10239 4857 10248 4913
rect 10174 4848 10248 4857
rect 10050 4514 10056 4566
rect 10108 4514 10114 4566
rect 10050 4508 10114 4514
rect 8392 4351 8760 4415
rect 8392 4177 8456 4183
rect 8392 4125 8398 4177
rect 8450 4125 8456 4177
rect 6724 3947 6798 3954
rect 6724 3945 6740 3947
rect 6724 3889 6733 3945
rect 6792 3894 6798 3947
rect 6789 3889 6798 3894
rect 6724 3880 6798 3889
rect 8392 3946 8456 4125
rect 8392 3894 8398 3946
rect 8450 3894 8456 3946
rect 8392 3590 8456 3894
rect 8392 3538 8398 3590
rect 8450 3538 8456 3590
rect 6734 3466 6798 3472
rect 6734 3414 6740 3466
rect 6792 3414 6798 3466
rect 6734 3408 6798 3414
rect 6740 2524 6792 3408
rect 8392 3297 8456 3538
rect 8392 3245 8398 3297
rect 8450 3245 8456 3297
rect 8392 3239 8456 3245
rect 6952 2915 7026 2924
rect 6952 2859 6961 2915
rect 7017 2859 7026 2915
rect 6952 2850 7026 2859
rect 6729 2515 6803 2524
rect 6729 2459 6738 2515
rect 6794 2459 6803 2515
rect 6729 2450 6803 2459
rect 6533 2315 6607 2324
rect 6533 2259 6542 2315
rect 6598 2259 6607 2315
rect 6533 2250 6607 2259
rect 6740 2121 6792 2450
rect 6740 1772 6792 2069
rect 6963 1983 7015 2850
rect 8696 2558 8760 4351
rect 10045 4410 10119 4421
rect 10045 4284 10054 4410
rect 10110 4284 10119 4410
rect 10045 4273 10119 4284
rect 8696 2506 8702 2558
rect 8754 2506 8760 2558
rect 8387 2315 8461 2324
rect 8387 2259 8396 2315
rect 8452 2259 8461 2315
rect 8387 2250 8461 2259
rect 6734 1766 6798 1772
rect 6734 1714 6740 1766
rect 6792 1714 6798 1766
rect 6734 1708 6798 1714
rect 6740 1354 6792 1708
rect 6963 1673 7015 1931
rect 8398 1772 8450 2250
rect 8392 1766 8456 1772
rect 8392 1714 8398 1766
rect 8450 1714 8456 1766
rect 8392 1708 8456 1714
rect 6963 1565 7015 1621
rect 6734 1348 6798 1354
rect 6734 1296 6740 1348
rect 6792 1296 6798 1348
rect 6734 1290 6798 1296
rect 6740 936 6792 1290
rect 6963 1255 7015 1513
rect 8398 1354 8450 1708
rect 8392 1348 8456 1354
rect 8392 1296 8398 1348
rect 8450 1296 8456 1348
rect 8392 1290 8456 1296
rect 6963 1147 7015 1203
rect 6734 930 6798 936
rect 6734 878 6740 930
rect 6792 878 6798 930
rect 6734 872 6798 878
rect 6740 518 6792 872
rect 6963 837 7015 1095
rect 8398 936 8450 1290
rect 8392 930 8456 936
rect 8392 878 8398 930
rect 8450 878 8456 930
rect 8392 872 8456 878
rect 6963 729 7015 785
rect 6734 512 6798 518
rect 6734 460 6740 512
rect 6792 460 6798 512
rect 6734 454 6798 460
rect 6740 100 6792 454
rect 6963 419 7015 677
rect 8398 518 8450 872
rect 8392 512 8456 518
rect 8392 460 8398 512
rect 8450 460 8456 512
rect 8392 454 8456 460
rect 6963 311 7015 367
rect 6734 94 6798 100
rect 6734 42 6740 94
rect 6792 42 6798 94
rect 6734 36 6798 42
rect 6740 -318 6792 36
rect 6963 1 7015 259
rect 8398 100 8450 454
rect 8392 94 8456 100
rect 8392 42 8398 94
rect 8450 42 8456 94
rect 8392 36 8456 42
rect 6963 -107 7015 -51
rect 6734 -324 6798 -318
rect 6734 -376 6740 -324
rect 6792 -376 6798 -324
rect 6734 -382 6798 -376
rect 6740 -736 6792 -382
rect 6963 -417 7015 -159
rect 8398 -318 8450 36
rect 8392 -324 8456 -318
rect 8392 -376 8398 -324
rect 8450 -376 8456 -324
rect 8392 -382 8456 -376
rect 6963 -525 7015 -469
rect 6734 -742 6798 -736
rect 6734 -794 6740 -742
rect 6792 -794 6798 -742
rect 6734 -800 6798 -794
rect 6740 -1154 6792 -800
rect 6963 -835 7015 -577
rect 8398 -736 8450 -382
rect 8392 -742 8456 -736
rect 8392 -794 8398 -742
rect 8450 -794 8456 -742
rect 8392 -800 8456 -794
rect 6963 -943 7015 -887
rect 6734 -1160 6798 -1154
rect 6734 -1212 6740 -1160
rect 6792 -1212 6798 -1160
rect 6734 -1218 6798 -1212
rect 6740 -1391 6792 -1218
rect 6963 -1253 7015 -995
rect 8398 -1154 8450 -800
rect 8392 -1160 8456 -1154
rect 8392 -1212 8398 -1160
rect 8450 -1212 8456 -1160
rect 8392 -1218 8456 -1212
rect 8398 -1224 8450 -1218
rect 6963 -1311 7015 -1305
rect 6740 -1449 6792 -1443
rect 5230 -2069 5236 -2017
rect 5288 -2069 5294 -2017
rect 5230 -2079 5294 -2069
rect 8696 -2017 8760 2506
rect 10050 4177 10114 4273
rect 10050 4125 10056 4177
rect 10108 4125 10114 4177
rect 10050 3946 10114 4125
rect 10050 3894 10056 3946
rect 10108 3894 10114 3946
rect 10050 3590 10114 3894
rect 10312 3796 10368 5603
rect 10609 5569 10665 5716
rect 10539 5513 10665 5569
rect 10739 5596 10803 5900
rect 10739 5544 10745 5596
rect 10797 5544 10803 5596
rect 10416 4415 10490 4421
rect 10416 4410 10427 4415
rect 10479 4410 10490 4415
rect 10416 4284 10425 4410
rect 10481 4284 10490 4410
rect 10416 4279 10427 4284
rect 10479 4279 10490 4284
rect 10416 4273 10490 4279
rect 10303 3787 10377 3796
rect 10303 3731 10312 3787
rect 10368 3731 10377 3787
rect 10303 3722 10377 3731
rect 10539 3734 10595 5513
rect 10739 5462 10803 5544
rect 10739 5410 10745 5462
rect 10797 5410 10803 5462
rect 10739 5404 10803 5410
rect 10774 5096 10838 5102
rect 10774 5044 10780 5096
rect 10832 5044 10838 5096
rect 10635 4920 10709 4929
rect 10635 4864 10644 4920
rect 10700 4919 10709 4920
rect 10701 4867 10709 4919
rect 10700 4864 10709 4867
rect 10635 4855 10709 4864
rect 10643 4563 10707 4855
rect 10643 4511 10649 4563
rect 10701 4511 10707 4563
rect 10643 4207 10707 4511
rect 10643 4155 10649 4207
rect 10701 4155 10707 4207
rect 10643 3851 10707 4155
rect 10643 3799 10649 3851
rect 10701 3799 10707 3851
rect 10643 3793 10707 3799
rect 10774 4740 10838 5044
rect 10774 4688 10780 4740
rect 10832 4688 10838 4740
rect 10774 4421 10838 4688
rect 10774 4410 10848 4421
rect 10774 4384 10783 4410
rect 10774 4332 10780 4384
rect 10774 4284 10783 4332
rect 10839 4284 10848 4410
rect 10774 4273 10848 4284
rect 10940 4415 11014 4421
rect 10940 4410 10951 4415
rect 11003 4410 11014 4415
rect 10940 4284 10949 4410
rect 11005 4284 11014 4410
rect 10940 4279 10951 4284
rect 11003 4279 11014 4284
rect 10940 4273 11014 4279
rect 10774 4028 10838 4273
rect 10774 3976 10780 4028
rect 10832 3976 10838 4028
rect 10539 3729 10603 3734
rect 10539 3728 10704 3729
rect 10050 3538 10056 3590
rect 10108 3538 10114 3590
rect 10312 3613 10368 3722
rect 10539 3676 10545 3728
rect 10597 3676 10704 3728
rect 10539 3673 10704 3676
rect 10539 3670 10603 3673
rect 10545 3613 10609 3614
rect 10312 3608 10609 3613
rect 10312 3557 10551 3608
rect 10545 3556 10551 3557
rect 10603 3556 10609 3608
rect 10545 3550 10609 3556
rect 10050 3297 10114 3538
rect 10648 3500 10704 3673
rect 10774 3672 10838 3976
rect 10774 3620 10780 3672
rect 10832 3620 10838 3672
rect 10645 3494 10709 3500
rect 10645 3442 10651 3494
rect 10703 3442 10709 3494
rect 10645 3436 10709 3442
rect 10050 3245 10056 3297
rect 10108 3245 10114 3297
rect 10774 3316 10838 3620
rect 10774 3264 10780 3316
rect 10832 3264 10838 3316
rect 10774 3258 10838 3264
rect 10050 2248 10114 3245
rect 9854 2184 10114 2248
rect 9854 1983 9918 2184
rect 9854 1931 9860 1983
rect 9912 1931 9918 1983
rect 9854 1673 9918 1931
rect 9854 1621 9860 1673
rect 9912 1621 9918 1673
rect 9854 1565 9918 1621
rect 9854 1513 9860 1565
rect 9912 1513 9918 1565
rect 9854 1255 9918 1513
rect 9854 1203 9860 1255
rect 9912 1203 9918 1255
rect 9854 1147 9918 1203
rect 9854 1095 9860 1147
rect 9912 1095 9918 1147
rect 9854 837 9918 1095
rect 9854 785 9860 837
rect 9912 785 9918 837
rect 9854 729 9918 785
rect 9854 677 9860 729
rect 9912 677 9918 729
rect 9854 419 9918 677
rect 9854 367 9860 419
rect 9912 367 9918 419
rect 9854 311 9918 367
rect 9854 259 9860 311
rect 9912 259 9918 311
rect 9854 1 9918 259
rect 9854 -51 9860 1
rect 9912 -51 9918 1
rect 9854 -107 9918 -51
rect 9854 -159 9860 -107
rect 9912 -159 9918 -107
rect 9854 -417 9918 -159
rect 9854 -469 9860 -417
rect 9912 -469 9918 -417
rect 9854 -525 9918 -469
rect 9854 -577 9860 -525
rect 9912 -577 9918 -525
rect 9854 -835 9918 -577
rect 9854 -887 9860 -835
rect 9912 -887 9918 -835
rect 9854 -943 9918 -887
rect 9854 -995 9860 -943
rect 9912 -995 9918 -943
rect 9854 -1253 9918 -995
rect 9854 -1305 9860 -1253
rect 9912 -1305 9918 -1253
rect 9854 -1676 9918 -1305
rect 10050 2121 10114 2124
rect 10050 2069 10056 2121
rect 10108 2069 10114 2121
rect 10050 1766 10114 2069
rect 10050 1714 10056 1766
rect 10108 1714 10114 1766
rect 10050 1348 10114 1714
rect 10050 1296 10056 1348
rect 10108 1296 10114 1348
rect 10050 930 10114 1296
rect 10050 878 10056 930
rect 10108 878 10114 930
rect 10050 512 10114 878
rect 10050 460 10056 512
rect 10108 460 10114 512
rect 10050 94 10114 460
rect 10050 42 10056 94
rect 10108 42 10114 94
rect 10050 -324 10114 42
rect 10050 -376 10056 -324
rect 10108 -376 10114 -324
rect 10050 -742 10114 -376
rect 10050 -794 10056 -742
rect 10108 -794 10114 -742
rect 10050 -1160 10114 -794
rect 10050 -1212 10056 -1160
rect 10108 -1212 10114 -1160
rect 10050 -1391 10114 -1212
rect 10050 -1443 10056 -1391
rect 10108 -1443 10114 -1391
rect 10050 -1446 10114 -1443
rect 9845 -1685 9919 -1676
rect 9845 -1815 9854 -1685
rect 9910 -1815 9919 -1685
rect 9845 -1824 9919 -1815
rect 8696 -2069 8702 -2017
rect 8754 -2069 8760 -2017
rect 8696 -2075 8760 -2069
<< via2 >>
rect -610 9616 -554 9746
rect 106 9616 162 9746
rect 1764 9616 1820 9746
rect 5080 9616 5136 9746
rect 8396 9616 8452 9746
rect 10054 9616 10110 9746
rect 10743 9616 10799 9746
rect -352 7223 -296 7225
rect -352 7171 -350 7223
rect -350 7171 -298 7223
rect -298 7171 -296 7223
rect -352 7169 -296 7171
rect -352 6858 -296 6860
rect -352 6806 -350 6858
rect -350 6806 -298 6858
rect -298 6806 -296 6858
rect -352 6804 -296 6806
rect -615 5294 -559 5350
rect -382 5020 -326 5022
rect -382 4968 -380 5020
rect -380 4968 -328 5020
rect -328 4968 -326 5020
rect -382 4966 -326 4968
rect -98 4959 -42 5015
rect -640 4282 -584 4338
rect 3422 7169 3478 7223
rect 3422 7167 3424 7169
rect 3424 7167 3476 7169
rect 3476 7167 3478 7169
rect 106 4281 162 4409
rect -384 4132 -380 4184
rect -380 4132 -328 4184
rect -384 4128 -328 4132
rect -100 4122 -44 4178
rect -386 3900 -380 3951
rect -380 3900 -330 3951
rect -386 3895 -330 3900
rect -386 3544 -380 3594
rect -380 3544 -330 3594
rect -386 3538 -330 3544
rect -100 3538 -44 3594
rect 3418 3894 3424 3944
rect 3424 3894 3474 3944
rect 3418 3888 3474 3894
rect 3418 3538 3424 3588
rect 3424 3538 3474 3588
rect 3418 3532 3474 3538
rect 3142 2859 3198 2915
rect 354 -1815 410 -1685
rect 1764 2259 1820 2315
rect 3618 2659 3674 2715
rect 3422 2459 3478 2515
rect 6740 6804 6796 6859
rect 6740 6803 6792 6804
rect 6792 6803 6796 6804
rect 5080 4282 5136 4410
rect 4729 3059 4785 3115
rect 4304 2259 4360 2315
rect 5080 2659 5136 2715
rect 5959 2656 6015 2712
rect 10195 6074 10251 6130
rect 10611 6130 10667 6133
rect 10611 6078 10615 6130
rect 10615 6078 10667 6130
rect 10611 6077 10667 6078
rect 10183 4857 10239 4913
rect 6733 3894 6740 3945
rect 6740 3894 6789 3945
rect 6733 3889 6789 3894
rect 6961 2859 7017 2915
rect 6738 2459 6794 2515
rect 6542 2259 6598 2315
rect 10054 4284 10110 4410
rect 8396 2259 8452 2315
rect 10425 4284 10427 4410
rect 10427 4284 10479 4410
rect 10479 4284 10481 4410
rect 10312 3731 10368 3787
rect 10644 4919 10700 4920
rect 10644 4867 10649 4919
rect 10649 4867 10700 4919
rect 10644 4864 10700 4867
rect 10783 4384 10839 4410
rect 10783 4332 10832 4384
rect 10832 4332 10839 4384
rect 10783 4284 10839 4332
rect 10949 4284 10951 4410
rect 10951 4284 11003 4410
rect 11003 4284 11005 4410
rect 9854 -1815 9910 -1685
<< metal3 >>
rect -619 9746 10808 9755
rect -619 9616 -610 9746
rect -554 9616 106 9746
rect 162 9616 1764 9746
rect 1820 9616 5080 9746
rect 5136 9616 8396 9746
rect 8452 9616 10054 9746
rect 10110 9616 10743 9746
rect 10799 9616 10808 9746
rect -619 9607 10808 9616
rect -361 7225 -287 7234
rect 3417 7225 3483 7228
rect -361 7169 -352 7225
rect -296 7223 3483 7225
rect -296 7169 3422 7223
rect -361 7167 3422 7169
rect 3478 7167 3483 7223
rect -361 7165 3483 7167
rect -361 7160 -287 7165
rect 3417 7162 3483 7165
rect -361 6861 -287 6869
rect 6735 6861 6801 6864
rect -361 6860 6801 6861
rect -361 6804 -352 6860
rect -296 6859 6801 6860
rect -296 6804 6740 6859
rect -361 6803 6740 6804
rect 6796 6803 6801 6859
rect -361 6801 6801 6803
rect -361 6795 -287 6801
rect 6735 6798 6801 6801
rect 10186 6132 10260 6139
rect 10602 6133 10676 6142
rect 10602 6132 10611 6133
rect 10186 6130 10611 6132
rect 10186 6074 10195 6130
rect 10251 6077 10611 6130
rect 10667 6077 10676 6133
rect 10251 6074 10676 6077
rect 10186 6072 10676 6074
rect 10186 6065 10260 6072
rect 10602 6068 10676 6072
rect -701 5350 -550 5359
rect -701 5294 -615 5350
rect -559 5294 -550 5350
rect -701 5285 -550 5294
rect -391 5022 -317 5031
rect -391 4966 -382 5022
rect -326 5017 -317 5022
rect -107 5017 -33 5024
rect -326 5015 -33 5017
rect -326 4966 -98 5015
rect -391 4959 -98 4966
rect -42 4959 -33 5015
rect -391 4957 -33 4959
rect -107 4950 -33 4957
rect 10174 4920 10248 4922
rect 10635 4920 10709 4929
rect 10174 4913 10644 4920
rect 10174 4857 10183 4913
rect 10239 4864 10644 4913
rect 10700 4864 10709 4920
rect 10239 4860 10709 4864
rect 10239 4857 10248 4860
rect 10174 4848 10248 4857
rect 10635 4855 10709 4860
rect -649 4420 97 4421
rect 171 4420 11014 4421
rect -649 4410 11014 4420
rect -649 4409 5080 4410
rect -649 4338 106 4409
rect -649 4282 -640 4338
rect -584 4282 106 4338
rect -649 4281 106 4282
rect 162 4282 5080 4409
rect 5136 4284 10054 4410
rect 10110 4284 10425 4410
rect 10481 4284 10783 4410
rect 10839 4284 10949 4410
rect 11005 4284 11014 4410
rect 5136 4282 11014 4284
rect 162 4281 11014 4282
rect -649 4273 11014 4281
rect 97 4272 171 4273
rect -393 4184 -319 4193
rect -393 4128 -384 4184
rect -328 4182 -319 4184
rect -109 4182 -35 4187
rect -328 4178 -35 4182
rect -328 4128 -100 4178
rect -393 4122 -100 4128
rect -44 4122 -35 4178
rect -393 4119 -319 4122
rect -109 4113 -35 4122
rect -395 3951 -321 3960
rect 3409 3951 3483 3953
rect -395 3895 -386 3951
rect -330 3944 3483 3951
rect -330 3895 3418 3944
rect -395 3891 3418 3895
rect -395 3886 -321 3891
rect 3409 3888 3418 3891
rect 3474 3888 3483 3944
rect 3409 3879 3483 3888
rect 6724 3945 6798 3954
rect 6724 3889 6733 3945
rect 6789 3889 6798 3945
rect 6724 3880 6798 3889
rect 6724 3791 6784 3880
rect 10303 3791 10377 3796
rect -356 3787 10377 3791
rect -356 3731 10312 3787
rect 10368 3731 10377 3787
rect -356 3625 -296 3731
rect 10303 3722 10377 3731
rect -395 3594 -296 3625
rect -395 3538 -386 3594
rect -330 3565 -296 3594
rect -109 3594 -35 3603
rect 3409 3594 3483 3597
rect -330 3538 -321 3565
rect -395 3529 -321 3538
rect -109 3538 -100 3594
rect -44 3588 3483 3594
rect -44 3538 3418 3588
rect -109 3534 3418 3538
rect -109 3529 -35 3534
rect 3409 3532 3418 3534
rect 3474 3532 3483 3588
rect 3409 3523 3483 3532
rect 4720 3117 4794 3124
rect 1766 3115 8450 3117
rect 1766 3059 4729 3115
rect 4785 3059 8450 3115
rect 1766 3057 8450 3059
rect 4720 3050 4794 3057
rect 3133 2917 3207 2924
rect 6952 2917 7026 2924
rect 1766 2915 8450 2917
rect 1766 2859 3142 2915
rect 3198 2859 6961 2915
rect 7017 2859 8450 2915
rect 1766 2857 8450 2859
rect 3133 2850 3207 2857
rect 6952 2850 7026 2857
rect 3609 2717 3683 2724
rect 5071 2717 5145 2724
rect 5950 2717 6024 2721
rect 1766 2715 8450 2717
rect 1766 2659 3618 2715
rect 3674 2659 5080 2715
rect 5136 2712 8450 2715
rect 5136 2659 5959 2712
rect 1766 2657 5959 2659
rect 3609 2650 3683 2657
rect 5071 2650 5145 2657
rect 5950 2656 5959 2657
rect 6015 2657 8450 2712
rect 6015 2656 6024 2657
rect 5950 2647 6024 2656
rect 3413 2517 3487 2524
rect 6729 2517 6803 2524
rect 1766 2515 8450 2517
rect 1766 2459 3422 2515
rect 3478 2459 6738 2515
rect 6794 2459 8450 2515
rect 1766 2457 8450 2459
rect 3413 2450 3487 2457
rect 6729 2450 6803 2457
rect 1755 2317 1829 2324
rect 4295 2317 4369 2324
rect 6533 2317 6607 2324
rect 8387 2317 8461 2324
rect 1755 2315 8461 2317
rect 1755 2259 1764 2315
rect 1820 2259 4304 2315
rect 4360 2259 6542 2315
rect 6598 2259 8396 2315
rect 8452 2259 8461 2315
rect 1755 2257 8461 2259
rect 1755 2250 1829 2257
rect 4295 2250 4369 2257
rect 6533 2250 6607 2257
rect 8387 2250 8461 2257
rect 97 -1685 10045 -1676
rect 97 -1815 354 -1685
rect 410 -1815 9854 -1685
rect 9910 -1815 10045 -1685
rect 97 -1824 10045 -1815
use sky130_fd_pr__nfet_g5v0d10v5_GG9S2Z  sky130_fd_pr__nfet_g5v0d10v5_GG9S2Z_0
timestamp 1712930986
transform 1 0 -483 0 1 4245
box -328 -1039 328 1039
use sky130_fd_pr__nfet_g5v0d10v5_HZHY2Z  sky130_fd_pr__nfet_g5v0d10v5_HZHY2Z_0
timestamp 1712930986
transform 0 -1 10707 -1 0 4180
box -1089 -327 1089 327
use sky130_fd_pr__nfet_g5v0d10v5_T82T27  sky130_fd_pr__nfet_g5v0d10v5_T82T27_1
timestamp 1712930986
transform 1 0 5108 0 1 3711
box -5173 -505 5173 505
use sky130_fd_pr__nfet_g5v0d10v5_ZV8547  sky130_fd_pr__nfet_g5v0d10v5_ZV8547_0
timestamp 1712930986
transform 1 0 5108 0 1 339
box -5173 -1821 5173 1821
use sky130_fd_pr__pfet_g5v0d10v5_3HV7M9  sky130_fd_pr__pfet_g5v0d10v5_3HV7M9_0
timestamp 1712930986
transform 1 0 5108 0 1 4807
box -5203 -362 5203 362
use sky130_fd_pr__pfet_g5v0d10v5_5H9LZ4  sky130_fd_pr__pfet_g5v0d10v5_5H9LZ4_0
timestamp 1712930986
transform 1 0 -453 0 1 6670
box -358 -909 358 909
use sky130_fd_pr__pfet_g5v0d10v5_5HV9F5  sky130_fd_pr__pfet_g5v0d10v5_5HV9F5_0
timestamp 1712930986
transform 1 0 5108 0 1 8612
box -5203 -909 5203 909
use sky130_fd_pr__pfet_g5v0d10v5_5HVT2F  sky130_fd_pr__pfet_g5v0d10v5_5HVT2F_0
timestamp 1712930986
transform 1 0 5108 0 1 6436
box -5203 -1457 5203 1457
use sky130_fd_pr__pfet_g5v0d10v5_W8MWAU  sky130_fd_pr__pfet_g5v0d10v5_W8MWAU_0
timestamp 1712930986
transform 0 -1 10673 -1 0 6460
box -1119 -362 1119 362
<< labels >>
rlabel metal2 3424 4230 3424 4230 7 vm
rlabel metal2 3418 3596 3418 3596 7 vn
flabel comment s 9285 3504 9285 3504 0 FreeSans 1600 0 0 0 dum
flabel comment s 7627 3504 7627 3504 0 FreeSans 1600 0 0 0 Mta
flabel comment s 5969 3504 5969 3504 0 FreeSans 1600 0 0 0 Mta
flabel comment s 4311 3504 4311 3504 0 FreeSans 1600 0 0 0 Mb
flabel comment s 2653 3504 2653 3504 0 FreeSans 1600 0 0 0 Mb
flabel comment s 995 3504 995 3504 0 FreeSans 1600 0 0 0 dum
flabel comment s 995 3864 995 3864 0 FreeSans 1600 0 0 0 dum
flabel comment s 2653 3864 2653 3864 0 FreeSans 1600 0 0 0 Mnn0
flabel comment s 4311 3864 4311 3864 0 FreeSans 1600 0 0 0 Mnn0
flabel comment s 5969 3864 5969 3864 0 FreeSans 1600 0 0 0 Mnn1
flabel comment s 7627 3864 7627 3864 0 FreeSans 1600 0 0 0 Mnn1
flabel comment s 9285 3864 9285 3864 0 FreeSans 1600 0 0 0 dum
flabel comment s 9285 4824 9285 4824 0 FreeSans 1600 0 0 0 dum
flabel comment s 7627 4824 7627 4824 0 FreeSans 1600 0 0 0 Mpp1
flabel comment s 5969 4824 5969 4824 0 FreeSans 1600 0 0 0 Mpp1
flabel comment s 4311 4824 4311 4824 0 FreeSans 1600 0 0 0 Mpp0
flabel comment s 2653 4824 2653 4824 0 FreeSans 1600 0 0 0 Mpp0
flabel comment s 995 4824 995 4824 0 FreeSans 1600 0 0 0 dum
flabel comment s -452 6161 -452 6161 0 FreeSans 800 0 0 0 Mt0
flabel comment s -452 6526 -452 6526 0 FreeSans 800 0 0 0 Minv1
flabel comment s -452 6891 -452 6891 0 FreeSans 800 0 0 0 Ml3
flabel comment s -452 7256 -452 7256 0 FreeSans 800 0 0 0 Ml4
flabel comment s -479 3464 -479 3464 0 FreeSans 800 0 0 0 Ml2
flabel comment s -479 4559 -479 4559 0 FreeSans 800 0 0 0 Minv0
flabel comment s -479 4924 -479 4924 0 FreeSans 800 0 0 0 Mt1
flabel comment s -488 4217 -488 4217 0 FreeSans 800 0 0 0 Ml0
flabel comment s -488 3861 -488 3861 0 FreeSans 800 0 0 0 Ml1
flabel metal3 -624 5359 -624 5359 7 FreeSans 1200 0 0 0 ibias
port 2 w
flabel metal2 -765 5650 -765 5650 7 FreeSans 1200 0 0 0 ena
port 4 w
flabel metal2 -205 5718 -205 5718 7 FreeSans 800 0 0 0 ena_b
flabel metal2 6740 4230 6740 4230 7 FreeSans 800 0 0 0 n0
flabel metal3 1755 2317 1755 2317 7 FreeSans 800 0 0 0 vnn
flabel metal3 1766 2517 1766 2517 7 FreeSans 800 0 0 0 vt
flabel metal3 1766 2717 1766 2717 7 FreeSans 800 0 0 0 vpp
flabel metal3 1766 2917 1766 2917 7 FreeSans 1200 0 0 0 vinn
port 5 w
flabel metal3 1766 3117 1766 3117 7 FreeSans 1200 0 0 0 vinp
port 6 w
flabel metal2 10704 3729 10704 3729 3 FreeSans 800 0 0 0 n1
flabel metal3 10472 6132 10472 6132 1 FreeSans 1200 0 0 0 out
port 3 n
flabel metal3 97 -1676 97 -1676 7 FreeSans 1200 0 0 0 avss
port 7 w
flabel comment s 995 5324 995 5324 0 FreeSans 1600 0 0 0 dum
flabel comment s 2653 5324 2653 5324 0 FreeSans 1600 0 0 0 Mh0
flabel comment s 4311 5324 4311 5324 0 FreeSans 1600 0 0 0 Mh0
flabel comment s 5969 5324 5969 5324 0 FreeSans 1600 0 0 0 Mh1
flabel comment s 7627 5324 7627 5324 0 FreeSans 1600 0 0 0 Mh1
flabel comment s 9285 5324 9285 5324 0 FreeSans 1600 0 0 0 dum
flabel metal3 -619 9751 -619 9751 7 FreeSans 1200 0 0 0 avdd
port 1 w
flabel comment s 973 9194 973 9194 0 FreeSans 1600 0 0 0 dum
flabel comment s 2631 9194 2631 9194 0 FreeSans 1600 0 0 0 Mld1
flabel comment s 4289 9194 4289 9194 0 FreeSans 1600 0 0 0 Mld1
flabel comment s 5947 9194 5947 9194 0 FreeSans 1600 0 0 0 Mld0
flabel comment s 7605 9194 7605 9194 0 FreeSans 1600 0 0 0 Mld0
flabel comment s 9263 9194 9263 9194 0 FreeSans 1600 0 0 0 dum
flabel space 2662 -1130 2662 -1130 0 FreeSans 1600 0 0 0 Mi0
flabel space 7646 -1130 7646 -1130 0 FreeSans 1600 0 0 0 Mi0
flabel space 2634 1800 2634 1800 0 FreeSans 1600 0 0 0 Mi0
flabel space 7618 1790 7618 1790 0 FreeSans 1600 0 0 0 Mi0
flabel space 4324 1808 4324 1808 0 FreeSans 1600 0 0 0 Mi1
flabel space 6022 1808 6022 1808 0 FreeSans 1600 0 0 0 Mi1
flabel space 4332 -1130 4332 -1130 0 FreeSans 1600 0 0 0 Mi1
flabel space 5986 -1110 5986 -1110 0 FreeSans 1600 0 0 0 Mi1
flabel space 10720 7260 10720 7260 0 FreeSans 480 0 0 0 Minv5
flabel space 10698 6192 10698 6192 0 FreeSans 480 0 0 0 Minv5
flabel space 10688 6008 10688 6008 0 FreeSans 480 0 0 0 Minv5
flabel space 10698 5834 10698 5834 0 FreeSans 480 0 0 0 Minv3
flabel space 10702 5664 10702 5664 0 FreeSans 480 0 0 0 Minv3
flabel space 10720 4972 10720 4972 0 FreeSans 480 0 0 0 Minv4
flabel space 10734 3898 10734 3898 0 FreeSans 480 0 0 0 Minv4
flabel space 10734 3554 10734 3554 0 FreeSans 480 0 0 0 Minv2
flabel space 10730 3380 10730 3380 0 FreeSans 480 0 0 0 Minv2
flabel space 10734 4092 10734 4092 0 FreeSans 480 0 0 0 Minv4
<< end >>
