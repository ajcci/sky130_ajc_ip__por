magic
tech sky130A
magscale 1 2
timestamp 1713026247
<< dnwell >>
rect -2387 -2578 25767 1958
<< nwell >>
rect -2467 1752 25847 2038
rect -2467 -2372 -2181 1752
rect -1877 385 2073 1482
rect 25561 -2372 25847 1752
rect -2467 -2658 25847 -2372
<< pwell >>
rect -1874 -496 2076 227
<< nmos >>
rect -619 -266 -499 -66
rect -441 -266 -321 -66
rect -262 -266 -226 -66
rect -166 -266 -130 -66
rect -71 -266 29 -66
rect 87 -266 187 -66
rect 245 -266 445 -66
rect 503 -266 603 -66
rect 661 -266 761 -66
rect 819 -266 919 -66
rect 977 -266 1077 -66
<< ndiff >>
rect -677 -78 -619 -66
rect -677 -254 -665 -78
rect -631 -254 -619 -78
rect -677 -266 -619 -254
rect -499 -78 -441 -66
rect -499 -254 -487 -78
rect -453 -254 -441 -78
rect -499 -266 -441 -254
rect -321 -78 -262 -66
rect -321 -254 -309 -78
rect -275 -254 -262 -78
rect -321 -266 -262 -254
rect -226 -78 -166 -66
rect -226 -254 -213 -78
rect -179 -254 -166 -78
rect -226 -266 -166 -254
rect -130 -78 -71 -66
rect -130 -254 -117 -78
rect -83 -254 -71 -78
rect -130 -266 -71 -254
rect 29 -78 87 -66
rect 29 -254 41 -78
rect 75 -254 87 -78
rect 29 -266 87 -254
rect 187 -78 245 -66
rect 187 -254 199 -78
rect 233 -254 245 -78
rect 187 -266 245 -254
rect 445 -78 503 -66
rect 445 -254 457 -78
rect 491 -254 503 -78
rect 445 -266 503 -254
rect 603 -78 661 -66
rect 603 -254 615 -78
rect 649 -254 661 -78
rect 603 -266 661 -254
rect 761 -78 819 -66
rect 761 -254 773 -78
rect 807 -254 819 -78
rect 761 -266 819 -254
rect 919 -78 977 -66
rect 919 -254 931 -78
rect 965 -254 977 -78
rect 919 -266 977 -254
rect 1077 -78 1135 -66
rect 1077 -254 1089 -78
rect 1123 -254 1135 -78
rect 1077 -266 1135 -254
<< ndiffc >>
rect -665 -254 -631 -78
rect -487 -254 -453 -78
rect -309 -254 -275 -78
rect -213 -254 -179 -78
rect -117 -254 -83 -78
rect 41 -254 75 -78
rect 199 -254 233 -78
rect 457 -254 491 -78
rect 615 -254 649 -78
rect 773 -254 807 -78
rect 931 -254 965 -78
rect 1089 -254 1123 -78
<< psubdiff >>
rect -1838 157 -1778 191
rect 1980 157 2040 191
rect -1838 131 -1804 157
rect 2006 131 2040 157
rect -1838 -426 -1804 -400
rect 2006 -426 2040 -400
rect -1838 -460 -1778 -426
rect 1980 -460 2040 -426
<< nsubdiff >>
rect -2430 1981 25810 2001
rect -2430 1947 -2350 1981
rect 25730 1947 25810 1981
rect -2430 1927 25810 1947
rect -2430 1921 -2356 1927
rect -2430 -2541 -2410 1921
rect -2376 -2541 -2356 1921
rect 25736 1921 25810 1927
rect -1841 1412 -1781 1446
rect 1977 1412 2037 1446
rect -1841 1386 -1807 1412
rect 2003 1386 2037 1412
rect -1841 455 -1807 481
rect 2003 455 2037 481
rect -1841 421 -1781 455
rect 1977 421 2037 455
rect -2430 -2547 -2356 -2541
rect 25736 -2541 25756 1921
rect 25790 -2541 25810 1921
rect 25736 -2547 25810 -2541
rect -2430 -2567 25810 -2547
rect -2430 -2601 -2350 -2567
rect 25730 -2601 25810 -2567
rect -2430 -2621 25810 -2601
<< psubdiffcont >>
rect -1778 157 1980 191
rect -1838 -400 -1804 131
rect 2006 -400 2040 131
rect -1778 -460 1980 -426
<< nsubdiffcont >>
rect -2350 1947 25730 1981
rect -2410 -2541 -2376 1921
rect -1781 1412 1977 1446
rect -1841 481 -1807 1386
rect 2003 481 2037 1386
rect -1781 421 1977 455
rect 25756 -2541 25790 1921
rect -2350 -2601 25730 -2567
<< poly >>
rect -1653 821 -1623 837
rect -1689 805 -1623 821
rect -1689 771 -1673 805
rect -1639 771 -1623 805
rect -1689 755 -1623 771
rect -619 6 -499 22
rect -619 -28 -603 6
rect -515 -28 -499 6
rect -619 -66 -499 -28
rect -277 6 -211 22
rect -277 -28 -261 6
rect -227 -28 -211 6
rect -441 -66 -321 -40
rect -277 -44 -211 -28
rect -71 6 29 22
rect -71 -28 -55 6
rect 13 -28 29 6
rect -262 -66 -226 -44
rect -166 -66 -130 -40
rect -71 -66 29 -28
rect 87 6 187 22
rect 87 -28 103 6
rect 171 -28 187 6
rect 87 -66 187 -28
rect 245 6 445 22
rect 245 -28 261 6
rect 429 -28 445 6
rect 245 -66 445 -28
rect 503 6 603 22
rect 503 -28 519 6
rect 587 -28 603 6
rect 503 -66 603 -28
rect 661 6 761 22
rect 661 -28 677 6
rect 745 -28 761 6
rect 661 -66 761 -28
rect 819 6 919 22
rect 819 -28 835 6
rect 903 -28 919 6
rect 819 -66 919 -28
rect 977 6 1077 22
rect 977 -28 993 6
rect 1061 -28 1077 6
rect 977 -66 1077 -28
rect -619 -292 -499 -266
rect -441 -304 -321 -266
rect -262 -292 -226 -266
rect -166 -288 -130 -266
rect -441 -338 -425 -304
rect -337 -338 -321 -304
rect -441 -354 -321 -338
rect -181 -304 -115 -288
rect -71 -292 29 -266
rect 87 -292 187 -266
rect 245 -292 445 -266
rect 503 -292 603 -266
rect 661 -292 761 -266
rect 819 -292 919 -266
rect 977 -292 1077 -266
rect -181 -338 -165 -304
rect -131 -338 -115 -304
rect -181 -354 -115 -338
<< polycont >>
rect -1673 771 -1639 805
rect -603 -28 -515 6
rect -261 -28 -227 6
rect -55 -28 13 6
rect 103 -28 171 6
rect 261 -28 429 6
rect 519 -28 587 6
rect 677 -28 745 6
rect 835 -28 903 6
rect 993 -28 1061 6
rect -425 -338 -337 -304
rect -165 -338 -131 -304
<< locali >>
rect -2410 1947 -2350 1981
rect 25730 1947 25790 1981
rect -2410 1921 -2376 1947
rect 25756 1921 25790 1947
rect -1841 1412 -1781 1446
rect 1977 1412 2037 1446
rect -1841 1386 -1807 1412
rect 2003 1386 2037 1412
rect -1689 805 -1623 821
rect -1689 771 -1673 805
rect -1639 771 -1623 805
rect -1689 755 -1623 771
rect -1841 455 -1807 481
rect 2003 455 2037 481
rect -1841 421 -1781 455
rect 1977 421 2037 455
rect -1838 157 -1778 191
rect 1980 157 2040 191
rect -1838 131 -1804 157
rect 2006 131 2040 157
rect -619 -28 -603 6
rect -515 -28 -499 6
rect -277 -28 -261 6
rect -227 -28 -211 6
rect -71 -28 -55 6
rect 13 -28 29 6
rect 87 -28 103 6
rect 171 -28 187 6
rect 245 -28 261 6
rect 429 -28 445 6
rect 503 -28 519 6
rect 587 -28 603 6
rect 661 -28 677 6
rect 745 -28 761 6
rect 819 -28 835 6
rect 903 -28 919 6
rect 977 -28 993 6
rect 1061 -28 1077 6
rect -665 -78 -631 -62
rect -665 -270 -631 -254
rect -487 -78 -453 -62
rect -487 -270 -453 -254
rect -309 -78 -275 -62
rect -309 -270 -275 -254
rect -213 -78 -179 -62
rect -213 -270 -179 -254
rect -117 -78 -83 -62
rect -117 -270 -83 -254
rect 41 -78 75 -62
rect 41 -270 75 -254
rect 199 -78 233 -62
rect 199 -270 233 -254
rect 457 -78 491 -62
rect 457 -270 491 -254
rect 615 -78 649 -62
rect 615 -270 649 -254
rect 773 -78 807 -62
rect 773 -270 807 -254
rect 931 -78 965 -62
rect 931 -270 965 -254
rect 1089 -78 1123 -62
rect 1089 -270 1123 -254
rect -441 -338 -425 -304
rect -337 -338 -321 -304
rect -181 -338 -165 -304
rect -131 -338 -115 -304
rect -1838 -426 -1804 -400
rect 2006 -426 2040 -400
rect -1838 -460 -1778 -426
rect 1980 -460 2040 -426
rect -2410 -2567 -2376 -2541
rect 25756 -2567 25790 -2541
rect -2410 -2601 -2350 -2567
rect 25730 -2601 25790 -2567
<< viali >>
rect -2350 1947 25730 1981
rect 2230 1614 25330 1648
rect -41 1446 -7 1447
rect -1781 1412 1977 1446
rect -1673 771 -1639 805
rect -1781 421 1977 455
rect -1778 157 1980 191
rect -603 -28 -515 6
rect -261 -28 -227 6
rect -55 -28 13 6
rect 103 -28 171 6
rect 261 -28 429 6
rect 519 -28 587 6
rect 677 -28 745 6
rect 835 -28 903 6
rect 993 -28 1061 6
rect -665 -254 -631 -78
rect -487 -254 -453 -78
rect -309 -254 -275 -78
rect -213 -254 -179 -78
rect -117 -254 -83 -78
rect 41 -254 75 -78
rect 199 -254 233 -78
rect 457 -254 491 -78
rect 615 -254 649 -78
rect 773 -254 807 -78
rect 931 -254 965 -78
rect 1089 -254 1123 -78
rect -425 -338 -337 -304
rect -165 -338 -131 -304
rect -1778 -460 1980 -426
rect 2134 -2200 2168 1552
rect 25392 -2200 25426 1552
rect 2230 -2296 25330 -2262
rect -2350 -2601 25730 -2567
<< metal1 >>
rect -2430 1981 25810 2001
rect -2430 1947 -2350 1981
rect 25730 1947 25810 1981
rect -2430 1927 25810 1947
rect -2430 -2547 -2356 1927
rect -47 1457 -1 1459
rect 1993 1457 2049 1927
rect -1851 1447 2049 1457
rect -1851 1446 -41 1447
rect -7 1446 2049 1447
rect -1851 1412 -1781 1446
rect 1977 1412 2049 1446
rect -1851 1401 2049 1412
rect -1851 1288 -1795 1401
rect -47 1288 -1 1401
rect 1993 1288 2049 1401
rect -1851 1206 2049 1288
rect -1851 466 -1795 1206
rect -1741 1073 -1667 1084
rect -1741 1021 -1730 1073
rect -1678 1021 -1667 1073
rect -1617 1063 -1576 1150
rect -1572 1144 -1524 1206
rect -1523 1063 -1476 1150
rect -1251 1149 -1199 1206
rect -995 1063 -949 1206
rect -679 1063 -633 1206
rect -363 1063 -317 1206
rect -47 1063 -1 1206
rect 469 1063 515 1206
rect -1741 1010 -1667 1021
rect -1093 1054 -1029 1060
rect -1093 1002 -1087 1054
rect -1035 1002 -1029 1054
rect -1093 996 -1029 1002
rect -851 1052 -777 1063
rect -851 1000 -840 1052
rect -788 1000 -777 1052
rect -851 989 -777 1000
rect -535 1052 -461 1063
rect -535 1000 -524 1052
rect -472 1000 -461 1052
rect -535 989 -461 1000
rect -219 1052 -145 1063
rect -219 1000 -208 1052
rect -156 1000 -145 1052
rect -219 989 -145 1000
rect 197 1052 271 1063
rect 197 1000 208 1052
rect 260 1000 271 1052
rect 197 989 271 1000
rect 699 1052 773 1063
rect 699 1000 710 1052
rect 762 1000 773 1052
rect 699 989 773 1000
rect -1363 966 -1299 972
rect -1363 914 -1357 966
rect -1305 914 -1299 966
rect -1363 908 -1299 914
rect -1202 957 -1138 963
rect -1202 905 -1196 957
rect -1144 905 -1138 957
rect -1202 899 -1138 905
rect -115 829 -51 835
rect -1689 805 -1668 821
rect -1608 810 -1602 821
rect -1117 820 -1053 826
rect -1608 808 -1467 810
rect -1689 771 -1673 805
rect -1689 761 -1668 771
rect -1608 761 -1430 808
rect -1117 768 -1111 820
rect -1059 768 -1053 820
rect -847 776 -149 822
rect -115 777 -109 829
rect -57 777 -51 829
rect 805 822 853 1206
rect 1043 1063 1089 1206
rect 1359 1063 1405 1206
rect 1675 1063 1721 1206
rect 885 1052 959 1063
rect 885 1000 896 1052
rect 948 1000 959 1052
rect 885 989 959 1000
rect 1187 1052 1261 1063
rect 1187 1000 1198 1052
rect 1250 1000 1261 1052
rect 1187 989 1261 1000
rect 1503 1052 1577 1063
rect 1503 1000 1514 1052
rect 1566 1000 1577 1052
rect 1503 989 1577 1000
rect 1819 1052 1893 1063
rect 1819 1000 1830 1052
rect 1882 1000 1893 1052
rect 1819 989 1893 1000
rect 1425 823 1489 829
rect -115 771 -51 777
rect 201 811 525 822
rect 201 776 310 811
rect -1117 762 -1053 768
rect -1689 760 -1608 761
rect -1689 755 -1623 760
rect 304 759 310 776
rect 362 776 525 811
rect 957 808 1021 814
rect 362 759 368 776
rect 304 753 368 759
rect 957 756 963 808
rect 1015 756 1021 808
rect 1033 776 1257 822
rect 1425 771 1431 823
rect 1483 771 1489 823
rect 1507 776 1731 822
rect 1425 765 1489 771
rect 957 750 1021 756
rect 1993 466 2049 1206
rect -1851 455 2049 466
rect -1851 421 -1781 455
rect 1977 421 2049 455
rect -1851 410 2049 421
rect 2105 1648 24342 1699
rect 24441 1648 25469 1699
rect 2105 1614 2230 1648
rect 25330 1614 25469 1648
rect 2105 1600 24342 1614
rect 24441 1600 25469 1614
rect 2105 1552 2204 1600
rect -1848 191 2052 202
rect -1848 157 -1778 191
rect 1980 157 2052 191
rect -1848 146 2052 157
rect -1848 -381 -1792 146
rect 673 45 737 51
rect -550 34 -239 45
rect 53 39 117 45
rect -550 28 -207 34
rect -550 12 -265 28
rect -615 6 -265 12
rect -615 -28 -603 6
rect -515 -3 -265 6
rect -515 -28 -503 -3
rect -615 -34 -503 -28
rect -273 -24 -265 -3
rect -213 -24 -207 28
rect 53 12 59 39
rect -273 -28 -261 -24
rect -227 -28 -207 -24
rect -273 -30 -207 -28
rect -67 6 59 12
rect 111 12 117 39
rect 322 36 386 42
rect 322 12 328 36
rect 111 6 183 12
rect -67 -28 -55 6
rect 13 -13 59 6
rect 13 -28 103 -13
rect 171 -28 183 6
rect -273 -34 -215 -30
rect -67 -34 183 -28
rect 249 6 328 12
rect 380 12 386 36
rect 673 12 679 45
rect 380 6 441 12
rect 249 -28 261 6
rect 429 -28 441 6
rect 249 -34 441 -28
rect 507 6 599 12
rect 507 -28 519 6
rect 587 -28 599 6
rect 507 -34 599 -28
rect 665 6 679 12
rect 731 12 737 45
rect 997 33 1061 39
rect 997 12 1003 33
rect 731 6 757 12
rect 665 -28 677 6
rect 745 -28 757 6
rect 665 -34 757 -28
rect 823 6 915 12
rect 823 -28 835 6
rect 903 -28 915 6
rect 823 -34 915 -28
rect 981 6 1003 12
rect 1055 12 1061 33
rect 1055 6 1073 12
rect 981 -28 993 6
rect 1061 -28 1073 6
rect 981 -34 1073 -28
rect -671 -78 -625 -66
rect -671 -132 -665 -78
rect -681 -138 -665 -132
rect -631 -132 -625 -78
rect -493 -78 -447 -66
rect -631 -138 -617 -132
rect -681 -190 -675 -138
rect -623 -190 -617 -138
rect -681 -196 -665 -190
rect -671 -254 -665 -196
rect -631 -196 -617 -190
rect -631 -254 -625 -196
rect -671 -266 -625 -254
rect -493 -254 -487 -78
rect -453 -254 -447 -78
rect -315 -78 -269 -66
rect -315 -189 -309 -78
rect -336 -195 -309 -189
rect -336 -247 -330 -195
rect -336 -253 -309 -247
rect -493 -298 -447 -254
rect -315 -254 -309 -253
rect -275 -254 -269 -78
rect -219 -78 -173 -66
rect -219 -182 -213 -78
rect -222 -188 -213 -182
rect -179 -182 -173 -78
rect -123 -78 -77 -66
rect -179 -188 -158 -182
rect -222 -240 -216 -188
rect -164 -240 -158 -188
rect -222 -246 -213 -240
rect -315 -266 -269 -254
rect -219 -254 -213 -246
rect -179 -246 -158 -240
rect -179 -254 -173 -246
rect -219 -266 -173 -254
rect -123 -254 -117 -78
rect -83 -254 -77 -78
rect 35 -78 81 -66
rect 35 -192 41 -78
rect -123 -298 -77 -254
rect 21 -203 41 -192
rect 75 -192 81 -78
rect 193 -78 239 -66
rect 75 -203 95 -192
rect 21 -255 32 -203
rect 84 -255 95 -203
rect 21 -266 95 -255
rect 193 -254 199 -78
rect 233 -254 239 -78
rect 451 -78 497 -66
rect 451 -192 457 -78
rect -493 -304 -325 -298
rect -493 -338 -425 -304
rect -337 -338 -325 -304
rect -177 -304 -77 -298
rect -177 -338 -165 -304
rect -131 -338 -77 -304
rect -493 -344 -322 -338
rect -177 -344 -77 -338
rect -373 -381 -322 -344
rect -123 -381 -77 -344
rect 193 -381 239 -254
rect 423 -203 457 -192
rect 423 -255 434 -203
rect 491 -254 497 -78
rect 486 -255 497 -254
rect 423 -266 497 -255
rect 530 -381 578 -34
rect 609 -78 655 -66
rect 609 -254 615 -78
rect 649 -254 655 -78
rect 767 -78 813 -66
rect 767 -192 773 -78
rect 609 -381 655 -254
rect 739 -203 773 -192
rect 739 -255 750 -203
rect 807 -254 813 -78
rect 802 -255 813 -254
rect 739 -266 813 -255
rect 845 -381 893 -34
rect 925 -78 971 -66
rect 925 -254 931 -78
rect 965 -254 971 -78
rect 1083 -78 1129 -66
rect 1083 -192 1089 -78
rect 925 -381 971 -254
rect 1069 -203 1089 -192
rect 1123 -192 1129 -78
rect 1123 -203 1143 -192
rect 1069 -255 1080 -203
rect 1132 -255 1143 -203
rect 1069 -266 1143 -255
rect 1996 -381 2052 146
rect 2105 -381 2134 1552
rect -1848 -426 2134 -381
rect -1848 -460 -1778 -426
rect 1980 -460 2134 -426
rect -1848 -480 2134 -460
rect 2094 -2200 2134 -480
rect 2168 -638 2204 1552
rect 25370 1552 25469 1600
rect 25146 1130 25290 1246
rect 2270 752 2691 868
rect 25146 374 25290 490
rect 2270 -4 2691 112
rect 25146 -382 25290 -266
rect 2168 -2200 2193 -638
rect 2270 -760 2691 -644
rect 25146 -1138 25290 -1022
rect 2270 -1516 2691 -1400
rect 25146 -1894 25290 -1778
rect 2514 -2141 2520 -2008
rect 2653 -2141 2659 -2008
rect 2094 -2228 2193 -2200
rect 25370 -2200 25392 1552
rect 25426 -2200 25469 1552
rect 25370 -2228 25469 -2200
rect 2094 -2262 25469 -2228
rect 2094 -2296 2230 -2262
rect 25330 -2296 25469 -2262
rect 2094 -2327 25469 -2296
rect 25736 -2547 25810 1927
rect -2430 -2567 25810 -2547
rect -2430 -2601 -2350 -2567
rect 25730 -2601 25810 -2567
rect -2430 -2621 25810 -2601
<< via1 >>
rect -1730 1021 -1678 1073
rect -1087 1002 -1035 1054
rect -840 1000 -788 1052
rect -524 1000 -472 1052
rect -208 1000 -156 1052
rect 208 1000 260 1052
rect 710 1000 762 1052
rect -1357 914 -1305 966
rect -1196 905 -1144 957
rect -1668 805 -1608 821
rect -1668 771 -1639 805
rect -1639 771 -1608 805
rect -1668 761 -1608 771
rect -1111 768 -1059 820
rect -109 777 -57 829
rect 896 1000 948 1052
rect 1198 1000 1250 1052
rect 1514 1000 1566 1052
rect 1830 1000 1882 1052
rect 310 759 362 811
rect 963 756 1015 808
rect 1431 771 1483 823
rect 24342 1648 24441 1699
rect 24342 1614 24441 1648
rect 24342 1600 24441 1614
rect -265 6 -213 28
rect -265 -24 -261 6
rect -261 -24 -227 6
rect -227 -24 -213 6
rect 59 6 111 39
rect 59 -13 103 6
rect 103 -13 111 6
rect 328 6 380 36
rect 328 -16 380 6
rect 679 6 731 45
rect 679 -7 731 6
rect 1003 6 1055 33
rect 1003 -19 1055 6
rect -675 -190 -665 -138
rect -665 -190 -631 -138
rect -631 -190 -623 -138
rect -330 -247 -309 -195
rect -309 -247 -278 -195
rect -216 -240 -213 -188
rect -213 -240 -179 -188
rect -179 -240 -164 -188
rect 32 -254 41 -203
rect 41 -254 75 -203
rect 75 -254 84 -203
rect 32 -255 84 -254
rect 434 -254 457 -203
rect 457 -254 486 -203
rect 434 -255 486 -254
rect 750 -254 773 -203
rect 773 -254 802 -203
rect 750 -255 802 -254
rect 1080 -254 1089 -203
rect 1089 -254 1123 -203
rect 1123 -254 1132 -203
rect 1080 -255 1132 -254
rect 2315 1320 2375 1380
rect 2520 -2141 2653 -2008
<< metal2 >>
rect 24337 1699 24446 1710
rect 24337 1600 24342 1699
rect 24441 1600 24446 1699
rect 24337 1589 24446 1600
rect -676 1380 -620 1387
rect 2309 1380 2381 1387
rect -678 1378 -618 1380
rect -678 1322 -676 1378
rect -620 1322 -618 1378
rect -1741 1075 -1667 1084
rect -1741 1019 -1732 1075
rect -1676 1019 -1667 1075
rect -1741 1010 -1667 1019
rect -1093 1057 -1029 1060
rect -1093 1054 -923 1057
rect -1093 1002 -1087 1054
rect -1035 1002 -923 1054
rect -1093 997 -923 1002
rect -1093 996 -1029 997
rect -1363 966 -1299 972
rect -1363 914 -1357 966
rect -1305 914 -1299 966
rect -1202 958 -1138 963
rect -1363 908 -1299 914
rect -1240 957 -1138 958
rect -1668 821 -1608 827
rect -1668 154 -1608 761
rect -1363 760 -1307 908
rect -1378 751 -1307 760
rect -1322 695 -1307 751
rect -1378 686 -1307 695
rect -1668 98 -1666 154
rect -1610 98 -1608 154
rect -1668 96 -1608 98
rect -1666 89 -1610 96
rect -1363 -126 -1307 686
rect -1240 905 -1196 957
rect -1144 905 -1138 957
rect -1240 899 -1138 905
rect -1240 617 -1184 899
rect -983 884 -923 997
rect -851 1054 -777 1063
rect -851 998 -842 1054
rect -786 998 -777 1054
rect -851 989 -777 998
rect -983 828 -981 884
rect -925 828 -923 884
rect -983 826 -923 828
rect -1117 820 -1053 826
rect -1117 768 -1111 820
rect -1059 798 -1053 820
rect -981 819 -925 826
rect -1059 768 -1051 798
rect -1117 762 -1051 768
rect -1118 753 -1040 762
rect -1118 693 -1109 753
rect -1049 693 -1040 753
rect -1118 684 -1040 693
rect -1242 608 -1182 617
rect -1242 539 -1182 548
rect -839 606 -765 615
rect -839 550 -830 606
rect -774 550 -765 606
rect -839 545 -765 550
rect -678 608 -618 1322
rect 2309 1320 2315 1380
rect 2375 1320 2381 1380
rect 2309 1313 2381 1320
rect -111 1248 -55 1255
rect -113 1246 -53 1248
rect -113 1190 -111 1246
rect -55 1190 -53 1246
rect -535 1054 -461 1063
rect -535 998 -526 1054
rect -470 998 -461 1054
rect -535 989 -461 998
rect -413 1060 -353 1069
rect -1365 -135 -1305 -126
rect -1365 -204 -1305 -195
rect -832 -243 -772 545
rect -678 539 -618 548
rect -413 -87 -353 1000
rect -219 1054 -145 1063
rect -219 998 -210 1054
rect -154 998 -145 1054
rect -219 989 -145 998
rect -227 886 -167 895
rect -113 835 -53 1190
rect 435 1063 495 1072
rect 197 1054 271 1063
rect 197 998 206 1054
rect 262 998 271 1054
rect 197 989 271 998
rect 699 1060 773 1063
rect 435 994 495 1003
rect 676 1054 773 1060
rect 676 998 708 1054
rect 764 998 773 1054
rect -227 817 -167 826
rect -115 829 -51 835
rect -225 169 -169 817
rect -115 777 -109 829
rect -57 777 -51 829
rect -115 771 -51 777
rect 304 811 368 817
rect -113 329 -53 771
rect 304 759 310 811
rect 362 796 368 811
rect 362 759 384 796
rect 304 753 384 759
rect 328 479 384 753
rect 316 470 384 479
rect 372 414 384 470
rect 316 405 384 414
rect -113 273 -111 329
rect -55 273 -53 329
rect -113 271 -53 273
rect 55 331 115 340
rect -111 264 -55 271
rect 55 262 115 271
rect -225 113 -95 169
rect -292 43 -218 52
rect -292 -13 -283 43
rect -227 34 -218 43
rect -227 28 -207 34
rect -292 -22 -265 -13
rect -271 -24 -265 -22
rect -213 -24 -207 28
rect -271 -30 -207 -24
rect -690 -132 -634 -128
rect -690 -137 -617 -132
rect -634 -138 -617 -137
rect -623 -190 -617 -138
rect -413 -143 -411 -87
rect -355 -143 -353 -87
rect -151 -99 -95 113
rect 57 149 113 262
rect 57 93 245 149
rect 57 45 113 93
rect 53 39 117 45
rect 53 -13 59 39
rect 111 -13 117 39
rect 53 -19 117 -13
rect 21 -87 30 -85
rect -413 -145 -353 -143
rect -411 -152 -355 -145
rect -201 -155 -95 -99
rect 17 -143 30 -87
rect 21 -145 30 -143
rect 90 -145 99 -85
rect -201 -182 -145 -155
rect -222 -188 -145 -182
rect -634 -193 -617 -190
rect -690 -196 -617 -193
rect -336 -195 -272 -189
rect -690 -202 -634 -196
rect -336 -205 -330 -195
rect -483 -243 -330 -205
rect -832 -247 -330 -243
rect -278 -247 -272 -195
rect -222 -240 -216 -188
rect -164 -226 -145 -188
rect 30 -192 86 -145
rect 21 -203 95 -192
rect -164 -235 -144 -226
rect -222 -246 -200 -240
rect -832 -253 -272 -247
rect -832 -265 -306 -253
rect -832 -303 -392 -265
rect 21 -255 32 -203
rect 84 -255 95 -203
rect 21 -266 95 -255
rect -200 -300 -144 -291
rect 189 -391 245 93
rect 328 42 384 405
rect 322 36 386 42
rect 322 -16 328 36
rect 380 -16 386 36
rect 322 -22 386 -16
rect 437 -192 493 994
rect 676 989 773 998
rect 885 1054 959 1063
rect 885 998 894 1054
rect 950 998 959 1054
rect 885 989 959 998
rect 1187 1054 1261 1063
rect 1187 998 1196 1054
rect 1252 998 1261 1054
rect 1187 989 1261 998
rect 1503 1054 1577 1063
rect 1503 998 1512 1054
rect 1568 998 1577 1054
rect 1503 989 1577 998
rect 1666 1057 1726 1066
rect 676 655 732 989
rect 888 921 944 989
rect 799 865 944 921
rect 674 646 734 655
rect 674 577 734 586
rect 676 51 732 577
rect 799 481 855 865
rect 1425 823 1489 829
rect 957 808 1021 814
rect 957 756 963 808
rect 1015 756 1021 808
rect 1425 771 1431 823
rect 1483 771 1489 823
rect 1425 765 1489 771
rect 957 750 1021 756
rect 957 644 1017 750
rect 957 588 959 644
rect 1015 588 1017 644
rect 957 586 1017 588
rect 1206 648 1266 657
rect 959 579 1015 586
rect 1206 579 1266 588
rect 797 472 857 481
rect 797 403 857 412
rect 999 455 1059 464
rect 673 45 737 51
rect 673 -7 679 45
rect 731 -7 737 45
rect 673 -13 737 -7
rect 799 -122 855 403
rect 999 386 1059 395
rect 1001 39 1057 386
rect 997 33 1061 39
rect 997 -19 1003 33
rect 1055 -19 1061 33
rect 997 -25 1061 -19
rect 1208 -120 1264 579
rect 1427 453 1487 765
rect 1666 646 1726 997
rect 1819 1054 1893 1063
rect 1819 998 1828 1054
rect 1884 998 1893 1054
rect 1819 989 1893 998
rect 1666 590 1668 646
rect 1724 590 1726 646
rect 1666 588 1726 590
rect 1668 581 1724 588
rect 1427 397 1429 453
rect 1485 397 1487 453
rect 1427 395 1487 397
rect 1429 388 1485 395
rect 745 -178 855 -122
rect 1076 -176 1264 -120
rect 745 -192 813 -178
rect 1076 -192 1143 -176
rect 423 -203 497 -192
rect 423 -255 434 -203
rect 486 -255 497 -203
rect 423 -266 497 -255
rect 739 -203 813 -192
rect 739 -255 750 -203
rect 802 -255 813 -203
rect 739 -266 813 -255
rect 1069 -203 1143 -192
rect 1069 -233 1080 -203
rect 1132 -233 1143 -203
rect 1069 -266 1076 -233
rect 1136 -266 1143 -233
rect 1076 -302 1136 -293
rect 187 -400 247 -391
rect 2535 -400 2591 -393
rect 187 -469 247 -460
rect 2533 -402 2593 -400
rect 2533 -458 2535 -402
rect 2591 -458 2593 -402
rect 2533 -2002 2593 -458
rect 2520 -2008 2653 -2002
rect 2520 -2329 2653 -2141
rect 2520 -2452 2525 -2329
rect 2648 -2452 2653 -2329
rect 2520 -2456 2653 -2452
rect 2525 -2461 2648 -2456
<< via2 >>
rect 24342 1600 24441 1699
rect -676 1322 -620 1378
rect -1732 1073 -1676 1075
rect -1732 1021 -1730 1073
rect -1730 1021 -1678 1073
rect -1678 1021 -1676 1073
rect -1732 1019 -1676 1021
rect -1378 695 -1322 751
rect -1666 98 -1610 154
rect -842 1052 -786 1054
rect -842 1000 -840 1052
rect -840 1000 -788 1052
rect -788 1000 -786 1052
rect -842 998 -786 1000
rect -981 828 -925 884
rect -1109 693 -1049 753
rect -1242 548 -1182 608
rect -830 550 -774 606
rect 2317 1322 2373 1378
rect -111 1190 -55 1246
rect -526 1052 -470 1054
rect -526 1000 -524 1052
rect -524 1000 -472 1052
rect -472 1000 -470 1052
rect -526 998 -470 1000
rect -413 1000 -353 1060
rect -678 548 -618 608
rect -1365 -195 -1305 -135
rect -210 1052 -154 1054
rect -210 1000 -208 1052
rect -208 1000 -156 1052
rect -156 1000 -154 1052
rect -210 998 -154 1000
rect -227 826 -167 886
rect 206 1052 262 1054
rect 206 1000 208 1052
rect 208 1000 260 1052
rect 260 1000 262 1052
rect 206 998 262 1000
rect 435 1003 495 1063
rect 708 1052 764 1054
rect 708 1000 710 1052
rect 710 1000 762 1052
rect 762 1000 764 1052
rect 708 998 764 1000
rect 316 414 372 470
rect -111 273 -55 329
rect 55 271 115 331
rect -283 28 -227 43
rect -283 -13 -265 28
rect -265 -13 -227 28
rect -690 -138 -634 -137
rect -690 -190 -675 -138
rect -675 -190 -634 -138
rect -411 -143 -355 -87
rect 30 -145 90 -85
rect -690 -193 -634 -190
rect -200 -240 -164 -235
rect -164 -240 -144 -235
rect -200 -291 -144 -240
rect 894 1052 950 1054
rect 894 1000 896 1052
rect 896 1000 948 1052
rect 948 1000 950 1052
rect 894 998 950 1000
rect 1196 1052 1252 1054
rect 1196 1000 1198 1052
rect 1198 1000 1250 1052
rect 1250 1000 1252 1052
rect 1196 998 1252 1000
rect 1512 1052 1568 1054
rect 1512 1000 1514 1052
rect 1514 1000 1566 1052
rect 1566 1000 1568 1052
rect 1512 998 1568 1000
rect 1666 997 1726 1057
rect 674 586 734 646
rect 959 588 1015 644
rect 1206 588 1266 648
rect 797 412 857 472
rect 999 395 1059 455
rect 1828 1052 1884 1054
rect 1828 1000 1830 1052
rect 1830 1000 1882 1052
rect 1882 1000 1884 1052
rect 1828 998 1884 1000
rect 1668 590 1724 646
rect 1429 397 1485 453
rect 1076 -255 1080 -233
rect 1080 -255 1132 -233
rect 1132 -255 1136 -233
rect 1076 -293 1136 -255
rect 187 -460 247 -400
rect 2535 -458 2591 -402
rect 2525 -2452 2648 -2329
<< metal3 >>
rect 24337 1704 24446 1710
rect 24337 1589 24446 1595
rect -681 1380 -615 1383
rect 2312 1380 2378 1383
rect -681 1378 2378 1380
rect -681 1322 -676 1378
rect -620 1322 2317 1378
rect 2373 1322 2378 1378
rect -681 1320 2378 1322
rect -681 1317 -615 1320
rect 2312 1317 2378 1320
rect -116 1248 -50 1251
rect -1727 1246 -50 1248
rect -1727 1190 -111 1246
rect -55 1190 -50 1246
rect -1727 1188 -50 1190
rect -1727 1084 -1667 1188
rect -116 1185 -50 1188
rect -1741 1075 -1667 1084
rect -1741 1019 -1732 1075
rect -1676 1019 -1667 1075
rect -418 1063 -348 1065
rect 430 1063 500 1068
rect -1741 1010 -1667 1019
rect -851 1060 435 1063
rect -851 1054 -413 1060
rect -851 998 -842 1054
rect -786 998 -526 1054
rect -470 1000 -413 1054
rect -353 1054 435 1060
rect -353 1000 -210 1054
rect -470 998 -210 1000
rect -154 998 206 1054
rect 262 1003 435 1054
rect 495 1054 773 1063
rect 495 1003 708 1054
rect 262 998 708 1003
rect 764 998 773 1054
rect -851 989 773 998
rect 885 1054 1261 1063
rect 885 998 894 1054
rect 950 998 1196 1054
rect 1252 998 1261 1054
rect 885 989 1261 998
rect 1503 1057 1893 1063
rect 1503 1054 1666 1057
rect 1503 998 1512 1054
rect 1568 998 1666 1054
rect 1503 997 1666 998
rect 1726 1054 1893 1057
rect 1726 998 1828 1054
rect 1884 998 1893 1054
rect 1726 997 1893 998
rect 1503 989 1893 997
rect -986 886 -920 889
rect -232 886 -162 891
rect -986 884 -227 886
rect -986 828 -981 884
rect -925 828 -227 884
rect -986 826 -227 828
rect -167 826 -162 886
rect -986 823 -920 826
rect -232 821 -162 826
rect -1383 753 -1317 756
rect -1114 753 -1044 758
rect -1383 751 -1109 753
rect -1383 695 -1378 751
rect -1322 695 -1109 751
rect -1383 693 -1109 695
rect -1049 693 -1044 753
rect -1383 690 -1317 693
rect -1114 688 -1044 693
rect 669 646 739 651
rect 954 646 1020 649
rect -1247 608 -1177 613
rect -835 608 -769 611
rect -683 608 -613 613
rect -1247 548 -1242 608
rect -1182 606 -678 608
rect -1182 550 -830 606
rect -774 550 -678 606
rect -1182 548 -678 550
rect -618 548 -613 608
rect 669 586 674 646
rect 734 644 1020 646
rect 734 588 959 644
rect 1015 588 1020 644
rect 734 586 1020 588
rect 669 581 739 586
rect 954 583 1020 586
rect 1201 648 1271 653
rect 1663 648 1729 651
rect 1201 588 1206 648
rect 1266 646 1729 648
rect 1266 590 1668 646
rect 1724 590 1729 646
rect 1266 588 1729 590
rect 1201 583 1271 588
rect 1663 585 1729 588
rect -1247 543 -1177 548
rect -835 545 -769 548
rect -683 543 -613 548
rect 311 472 377 475
rect 792 472 862 477
rect 311 470 797 472
rect 311 414 316 470
rect 372 414 797 470
rect 311 412 797 414
rect 857 460 1058 472
rect 857 455 1064 460
rect 1424 455 1490 458
rect 857 412 999 455
rect 311 409 377 412
rect 792 407 862 412
rect 994 395 999 412
rect 1059 453 1490 455
rect 1059 397 1429 453
rect 1485 397 1490 453
rect 1059 395 1490 397
rect 994 390 1064 395
rect 1424 392 1490 395
rect -116 331 -50 334
rect 50 331 120 336
rect -116 329 55 331
rect -116 273 -111 329
rect -55 273 55 329
rect -116 271 55 273
rect 115 271 120 331
rect -116 268 -50 271
rect 50 266 120 271
rect -1671 156 -1605 159
rect -1671 154 -232 156
rect -1671 98 -1666 154
rect -1610 98 -232 154
rect -1671 96 -232 98
rect -1671 93 -1605 96
rect -292 52 -232 96
rect -292 43 -218 52
rect -292 -13 -283 43
rect -227 -13 -218 43
rect -292 -22 -218 -13
rect -416 -85 -350 -82
rect 25 -85 95 -80
rect -416 -87 30 -85
rect -1370 -135 -1300 -130
rect -695 -135 -629 -132
rect -1370 -195 -1365 -135
rect -1305 -137 -629 -135
rect -1305 -193 -690 -137
rect -634 -193 -629 -137
rect -416 -143 -411 -87
rect -355 -143 30 -87
rect -416 -145 30 -143
rect 90 -145 95 -85
rect -416 -148 -350 -145
rect 25 -150 95 -145
rect -1305 -195 -629 -193
rect -1370 -200 -1300 -195
rect -695 -198 -629 -195
rect -205 -233 -139 -230
rect 1071 -233 1141 -228
rect -205 -235 1076 -233
rect -205 -291 -200 -235
rect -144 -291 1076 -235
rect -205 -293 1076 -291
rect 1136 -293 1141 -233
rect -205 -296 -139 -293
rect 1071 -298 1141 -293
rect 182 -400 252 -395
rect 2530 -400 2596 -397
rect 182 -460 187 -400
rect 247 -402 2596 -400
rect 247 -458 2535 -402
rect 2591 -458 2596 -402
rect 247 -460 2596 -458
rect 182 -465 252 -460
rect 2530 -463 2596 -460
rect 2520 -2326 24523 -2324
rect 2520 -2329 24391 -2326
rect 2520 -2452 2525 -2329
rect 2648 -2452 24391 -2329
rect 2520 -2457 24391 -2452
rect 24522 -2457 24528 -2326
<< via3 >>
rect 24337 1699 24446 1704
rect 24337 1600 24342 1699
rect 24342 1600 24441 1699
rect 24441 1600 24446 1699
rect 24337 1595 24446 1600
rect 24391 -2457 24522 -2326
<< metal4 >>
rect 24342 1705 24441 3852
rect 24336 1704 24447 1705
rect 24336 1595 24337 1704
rect 24446 1595 24447 1704
rect 24336 1594 24447 1595
rect 24390 -2326 24523 361
rect 24390 -2457 24391 -2326
rect 24522 -2457 24523 -2326
rect 24390 -2458 24523 -2457
<< via4 >>
rect 24317 3852 24589 4124
rect 24203 361 24523 681
<< metal5 >>
rect 24108 4124 24613 4148
rect 24108 3852 24317 4124
rect 24589 3852 24613 4124
rect 24108 3828 24613 3852
rect 23952 681 24547 705
rect 23952 361 24203 681
rect 24523 361 24547 681
rect 23952 337 24547 361
use sky130_fd_pr__cap_mim_m3_2_LUWKLG  sky130_fd_pr__cap_mim_m3_2_LUWKLG_0
timestamp 1712463840
transform 0 -1 4968 1 0 777
box -3349 -19200 3371 19200
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_0
timestamp 1712858885
transform 1 0 -1638 0 1 963
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_9QCJ55  sky130_fd_pr__pfet_01v8_9QCJ55_0
timestamp 1712722749
transform 1 0 363 0 1 927
box -452 -164 452 198
use sky130_fd_pr__pfet_01v8_C6GQGA  sky130_fd_pr__pfet_01v8_C6GQGA_0
timestamp 1712784588
transform 1 0 -1411 0 1 927
box -154 -164 154 198
use sky130_fd_pr__pfet_01v8_C64SS5  sky130_fd_pr__pfet_01v8_C64SS5_0
timestamp 1712722749
transform 1 0 -498 0 1 927
box -539 -164 539 198
use sky130_fd_pr__pfet_01v8_C68ZY6  sky130_fd_pr__pfet_01v8_C68ZY6_0
timestamp 1712722749
transform 1 0 1303 0 1 927
box -618 -164 618 198
use sky130_fd_pr__pfet_01v8_LAUYMQ  sky130_fd_pr__pfet_01v8_LAUYMQ_0
timestamp 1712784155
transform -1 0 -1068 0 -1 963
box -161 -200 161 200
use sky130_fd_pr__pfet_01v8_MA8JJJ  sky130_fd_pr__pfet_01v8_MA8JJJ_0
timestamp 1712784588
transform 1 0 -1547 0 1 999
box -112 -198 112 164
use sky130_fd_pr__pfet_01v8_MLERZ7  sky130_fd_pr__pfet_01v8_MLERZ7_0
timestamp 1712784588
transform 1 0 -1243 0 1 999
box -144 -198 144 164
use sky130_fd_pr__res_xhigh_po_1p41_ZB8LT7  sky130_fd_pr__res_xhigh_po_1p41_ZB8LT7_0
timestamp 1712975145
transform 0 1 13780 -1 0 -324
box -2008 -11682 2008 11682
<< labels >>
flabel metal3 s 1729 585 1729 585 0 FreeSans 1200 0 0 0 out
port 2 nsew
flabel metal1 s -1038 1288 -1038 1288 0 FreeSans 1200 0 0 0 dvdd
port 1 nsew
flabel metal1 s -1015 -381 -1015 -381 0 FreeSans 1200 0 0 0 dvss
port 4 nsew
flabel comment s 1460 954 1460 954 0 FreeSans 480 0 0 0 M8
flabel comment s 1618 954 1618 954 0 FreeSans 480 0 0 0 M8
flabel comment s 1778 958 1778 958 0 FreeSans 480 0 0 0 M8
flabel comment s 1304 952 1304 952 0 FreeSans 480 0 0 0 M6
flabel comment s 1148 952 1148 952 0 FreeSans 480 0 0 0 M6
flabel comment s 988 958 988 958 0 FreeSans 480 0 0 0 M6
flabel comment s 830 954 830 954 0 FreeSans 480 0 0 0 dum
flabel comment s 602 954 602 954 0 FreeSans 480 0 0 0 M4
flabel comment s 350 952 350 952 0 FreeSans 480 0 0 0 M4
flabel comment s 104 954 104 954 0 FreeSans 480 0 0 0 M4
flabel comment s -104 952 -104 952 0 FreeSans 480 0 0 0 M3
flabel comment s -266 958 -266 958 0 FreeSans 480 0 0 0 M3
flabel comment s -418 958 -418 958 0 FreeSans 480 0 0 0 M3
flabel comment s -574 954 -574 954 0 FreeSans 480 0 0 0 M3
flabel comment s -734 960 -734 960 0 FreeSans 480 0 0 0 M3
flabel comment s -886 960 -886 960 0 FreeSans 480 0 0 0 M3
flabel comment s -1022 960 -1022 960 0 FreeSans 480 0 0 0 dum
flabel comment s -1246 948 -1246 948 0 FreeSans 480 0 0 0 dum
flabel comment s -1410 1012 -1410 1012 0 FreeSans 480 0 0 0 M13
flabel comment s -1546 952 -1546 952 0 FreeSans 480 0 0 0 dum
flabel comment s -1638 1014 -1638 1014 0 FreeSans 480 0 0 0 M12
flabel comment s 1026 -156 1026 -156 0 FreeSans 480 0 0 0 M7
flabel comment s 870 -152 870 -152 0 FreeSans 480 0 0 0 dum
flabel comment s 708 -152 708 -152 0 FreeSans 480 0 0 0 M5
flabel comment s 552 -152 552 -152 0 FreeSans 480 0 0 0 dum
flabel comment s 338 -168 338 -168 0 FreeSans 480 0 0 0 M2
flabel comment s 136 -168 136 -168 0 FreeSans 480 0 0 0 M1
flabel comment s -26 -170 -26 -170 0 FreeSans 480 0 0 0 M1
flabel comment s -152 -182 -152 -182 0 FreeSans 480 0 0 0 dum
flabel comment s -246 -112 -246 -112 0 FreeSans 480 0 0 0 M9
flabel comment s -382 -176 -382 -176 0 FreeSans 480 0 0 0 dum
flabel comment s -566 -156 -566 -156 0 FreeSans 480 0 0 0 M11
flabel comment s -1118 1018 -1118 1018 0 FreeSans 480 0 0 0 M10
flabel metal2 s -1666 89 -1666 89 0 FreeSans 1200 0 0 0 ena
port 3 nsew
flabel metal2 s -1363 269 -1363 269 0 FreeSans 800 0 0 0 ena_b
flabel metal2 s -53 591 -53 591 0 FreeSans 800 0 0 0 in
flabel metal3 s 72 1063 72 1063 0 FreeSans 800 0 0 0 m
flabel metal2 s 1057 278 1057 278 0 FreeSans 800 0 0 0 n
flabel metal2 s -772 260 -772 260 0 FreeSans 800 0 0 0 vr
<< end >>
