* NGSPICE file created from por_dig.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

.subckt por_dig VGND VPWR force_pdn force_pdnb force_rc_osc force_short_oneshot osc_ck
+ osc_ena otrip[0] otrip[1] otrip[2] otrip_decoded[0] otrip_decoded[1] otrip_decoded[2]
+ otrip_decoded[3] otrip_decoded[4] otrip_decoded[5] otrip_decoded[6] otrip_decoded[7]
+ por_timed_out por_unbuf pwup_filt startup_timed_out
X_062_ net6 net4 net5 VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__nor3b_1
XFILLER_0_4_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_114_ clknet_1_1__leaf_osc_ck _005_ net23 VGND VGND VPWR VPWR cnt_por\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_7_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput20 net20 VGND VGND VPWR VPWR startup_timed_out sky130_fd_sc_hd__buf_2
XFILLER_0_13_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_12_Right_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_8_45 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_113_ clknet_1_1__leaf_osc_ck _004_ net23 VGND VGND VPWR VPWR cnt_st\[4\] sky130_fd_sc_hd__dfrtp_1
X_061_ net6 net5 net4 VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__nor3b_1
Xoutput8 net8 VGND VGND VPWR VPWR force_pdnb sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput10 net10 VGND VGND VPWR VPWR otrip_decoded[0] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_2_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_46 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_060_ net6 net5 net4 VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__nor3_1
XFILLER_0_4_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_112_ clknet_1_1__leaf_osc_ck _003_ net23 VGND VGND VPWR VPWR cnt_st\[3\] sky130_fd_sc_hd__dfrtp_1
Xhold10 cnt_por\[8\] VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_15_56 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput9 net9 VGND VGND VPWR VPWR osc_ena sky130_fd_sc_hd__buf_2
XFILLER_0_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput11 net11 VGND VGND VPWR VPWR otrip_decoded[1] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_2_37 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_10 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_12_Left_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_111_ clknet_1_1__leaf_osc_ck _002_ net23 VGND VGND VPWR VPWR cnt_st\[2\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_15_57 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold11 cnt_por\[1\] VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__dlygate4sd3_1
Xoutput12 net12 VGND VGND VPWR VPWR otrip_decoded[2] sky130_fd_sc_hd__buf_2
XFILLER_0_1_64 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_15_Left_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_0_Left_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_125__24 VGND VGND VPWR VPWR net24 _125__24/LO sky130_fd_sc_hd__conb_1
Xhold12 cnt_st\[4\] VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__dlygate4sd3_1
X_110_ clknet_1_1__leaf_osc_ck _001_ net22 VGND VGND VPWR VPWR cnt_st\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_76 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_58 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput13 net13 VGND VGND VPWR VPWR otrip_decoded[3] sky130_fd_sc_hd__buf_2
Xhold13 cnt_por\[0\] VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput14 net14 VGND VGND VPWR VPWR otrip_decoded[4] sky130_fd_sc_hd__buf_2
XFILLER_0_10_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_099_ _017_ _018_ VGND VGND VPWR VPWR _010_ sky130_fd_sc_hd__nor2_1
XFILLER_0_7_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput15 net15 VGND VGND VPWR VPWR otrip_decoded[5] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_098_ net21 _016_ net32 VGND VGND VPWR VPWR _018_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_7_Left_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_15_Right_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput16 net16 VGND VGND VPWR VPWR otrip_decoded[6] sky130_fd_sc_hd__buf_2
XFILLER_0_4_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_097_ cnt_por\[5\] net21 _016_ VGND VGND VPWR VPWR _017_ sky130_fd_sc_hd__and3_1
Xoutput17 net17 VGND VGND VPWR VPWR otrip_decoded[7] sky130_fd_sc_hd__buf_2
XFILLER_0_14_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_096_ cnt_por\[4\] _026_ _027_ net3 VGND VGND VPWR VPWR _016_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_6_42 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput18 net18 VGND VGND VPWR VPWR por_timed_out sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_079_ net31 _035_ _037_ VGND VGND VPWR VPWR _003_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_4_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_095_ net3 net21 _047_ VGND VGND VPWR VPWR _009_ sky130_fd_sc_hd__a21o_1
XFILLER_0_1_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput19 net19 VGND VGND VPWR VPWR por_unbuf sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_6_43 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_70 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_078_ net31 _035_ net20 VGND VGND VPWR VPWR _037_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_13_53 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout21 net19 VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_0_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_094_ cnt_por\[4\] _046_ VGND VGND VPWR VPWR _047_ sky130_fd_sc_hd__xor2_1
XPHY_EDGE_ROW_11_Left_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_077_ _035_ _036_ net20 VGND VGND VPWR VPWR _002_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_14_Left_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_093_ _045_ _046_ net3 net21 VGND VGND VPWR VPWR _008_ sky130_fd_sc_hd__a2bb2o_1
Xfanout22 net25 VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_3_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput1 force_pdn VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_076_ cnt_st\[2\] _032_ VGND VGND VPWR VPWR _036_ sky130_fd_sc_hd__or2_1
X_059_ _028_ _031_ VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout23 net25 VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_11_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_092_ _028_ _031_ net20 _026_ _027_ VGND VGND VPWR VPWR _046_ sky130_fd_sc_hd__o2111a_1
Xinput2 force_rc_osc VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__clkbuf_1
X_058_ _029_ _030_ VGND VGND VPWR VPWR _031_ sky130_fd_sc_hd__nand2_1
X_127_ clknet_1_0__leaf_osc_ck net27 net7 VGND VGND VPWR VPWR cnt_rsb sky130_fd_sc_hd__dfrtp_1
X_075_ cnt_st\[2\] _032_ VGND VGND VPWR VPWR _035_ sky130_fd_sc_hd__nand2_1
X_091_ cnt_por\[2\] _026_ net21 cnt_por\[3\] VGND VGND VPWR VPWR _045_ sky130_fd_sc_hd__a31oi_1
XFILLER_0_11_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput3 force_short_oneshot VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__clkbuf_2
X_074_ _033_ _034_ net20 VGND VGND VPWR VPWR _001_ sky130_fd_sc_hd__a21o_1
X_126_ clknet_1_0__leaf_osc_ck net26 net7 VGND VGND VPWR VPWR cnt_rsb_stg2 sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_057_ cnt_por\[7\] cnt_por\[9\] cnt_por\[8\] cnt_por\[10\] VGND VGND VPWR VPWR _030_
+ sky130_fd_sc_hd__and4_1
XFILLER_0_14_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_10 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_109_ clknet_1_1__leaf_osc_ck _000_ net22 VGND VGND VPWR VPWR cnt_st\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_8_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_090_ net3 net19 _043_ _044_ VGND VGND VPWR VPWR _007_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_9_47 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput4 otrip[0] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__dlymetal6s2s_1
XPHY_EDGE_ROW_3_Left_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_056_ cnt_por\[5\] cnt_por\[6\] VGND VGND VPWR VPWR _029_ sky130_fd_sc_hd__and2_1
X_125_ clknet_1_0__leaf_osc_ck net24 net7 VGND VGND VPWR VPWR cnt_rsb_stg1 sky130_fd_sc_hd__dfrtp_1
X_073_ cnt_st\[1\] cnt_st\[0\] net3 VGND VGND VPWR VPWR _034_ sky130_fd_sc_hd__or3_1
XPHY_EDGE_ROW_6_Left_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_108_ net29 _022_ VGND VGND VPWR VPWR _015_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_3_38 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_10_48 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput5 otrip[1] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__dlymetal6s2s_1
X_072_ _032_ VGND VGND VPWR VPWR _033_ sky130_fd_sc_hd__inv_2
X_055_ cnt_por\[4\] _026_ _027_ VGND VGND VPWR VPWR _028_ sky130_fd_sc_hd__nand3_1
X_124_ clknet_1_1__leaf_osc_ck _015_ net22 VGND VGND VPWR VPWR cnt_por\[10\] sky130_fd_sc_hd__dfrtp_1
X_107_ net30 _020_ VGND VGND VPWR VPWR _014_ sky130_fd_sc_hd__xor2_1
XPHY_EDGE_ROW_14_Right_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_49 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput6 otrip[2] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__dlymetal6s2s_1
X_071_ cnt_st\[0\] net3 cnt_st\[1\] VGND VGND VPWR VPWR _032_ sky130_fd_sc_hd__o21a_1
X_054_ cnt_por\[3\] cnt_por\[2\] VGND VGND VPWR VPWR _027_ sky130_fd_sc_hd__and2_1
XFILLER_0_8_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_123_ clknet_1_0__leaf_osc_ck _014_ net22 VGND VGND VPWR VPWR cnt_por\[9\] sky130_fd_sc_hd__dfrtp_1
X_106_ cnt_por\[7\] cnt_por\[9\] cnt_por\[8\] _019_ VGND VGND VPWR VPWR _022_ sky130_fd_sc_hd__and4_1
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput7 pwup_filt VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_070_ net3 net20 cnt_st\[0\] VGND VGND VPWR VPWR _000_ sky130_fd_sc_hd__or3b_1
X_053_ cnt_por\[1\] cnt_por\[0\] VGND VGND VPWR VPWR _026_ sky130_fd_sc_hd__and2_2
XFILLER_0_2_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_122_ clknet_1_0__leaf_osc_ck _013_ net22 VGND VGND VPWR VPWR cnt_por\[8\] sky130_fd_sc_hd__dfrtp_1
X_105_ _020_ _021_ VGND VGND VPWR VPWR _013_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_4_40 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_50 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_1__f_osc_ck clknet_0_osc_ck VGND VGND VPWR VPWR clknet_1_1__leaf_osc_ck
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_2_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_10_Left_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_052_ cnt_st\[4\] _025_ VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__and2_2
X_121_ clknet_1_0__leaf_osc_ck _012_ net22 VGND VGND VPWR VPWR cnt_por\[7\] sky130_fd_sc_hd__dfrtp_1
X_104_ cnt_por\[7\] _019_ net34 VGND VGND VPWR VPWR _021_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_15_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_120_ clknet_1_0__leaf_osc_ck _011_ net22 VGND VGND VPWR VPWR cnt_por\[6\] sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_051_ cnt_st\[1\] cnt_st\[0\] cnt_st\[2\] cnt_st\[3\] VGND VGND VPWR VPWR _025_ sky130_fd_sc_hd__and4_1
XFILLER_0_2_58 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_103_ cnt_por\[7\] cnt_por\[8\] _019_ VGND VGND VPWR VPWR _020_ sky130_fd_sc_hd__and3_1
XFILLER_0_15_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1 cnt_rsb VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_0_osc_ck osc_ck VGND VGND VPWR VPWR clknet_0_osc_ck sky130_fd_sc_hd__clkbuf_16
X_050_ net7 VGND VGND VPWR VPWR _024_ sky130_fd_sc_hd__inv_2
X_102_ net33 _019_ VGND VGND VPWR VPWR _012_ sky130_fd_sc_hd__xor2_1
Xhold2 cnt_rsb_stg1 VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_101_ net28 _017_ VGND VGND VPWR VPWR _011_ sky130_fd_sc_hd__xor2_1
XFILLER_0_8_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold3 cnt_rsb_stg2 VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_2_Left_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_100_ _028_ _031_ _016_ _029_ net20 VGND VGND VPWR VPWR _019_ sky130_fd_sc_hd__o2111a_1
XTAP_TAPCELL_ROW_7_44 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4 cnt_por\[6\] VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_5_Left_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_14_54 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold5 cnt_por\[10\] VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_15_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_55 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_089_ _026_ net19 cnt_por\[2\] VGND VGND VPWR VPWR _044_ sky130_fd_sc_hd__a21o_1
XFILLER_0_8_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold6 cnt_por\[9\] VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_15_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_088_ cnt_por\[2\] _026_ net19 VGND VGND VPWR VPWR _043_ sky130_fd_sc_hd__nand3_1
XPHY_EDGE_ROW_9_Left_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold7 cnt_st\[3\] VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_13_Right_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold8 cnt_por\[5\] VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__dlygate4sd3_1
X_087_ net3 net21 _041_ _042_ VGND VGND VPWR VPWR _006_ sky130_fd_sc_hd__a22o_1
Xclkbuf_1_0__f_osc_ck clknet_0_osc_ck VGND VGND VPWR VPWR clknet_1_0__leaf_osc_ck
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_4_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_086_ cnt_por\[0\] net21 net35 VGND VGND VPWR VPWR _042_ sky130_fd_sc_hd__a21o_1
XFILLER_0_3_43 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_069_ _028_ _031_ net20 VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__o21a_1
Xhold9 cnt_por\[7\] VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_4_39 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_085_ _026_ net21 VGND VGND VPWR VPWR _041_ sky130_fd_sc_hd__nand2_1
XFILLER_0_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_068_ _024_ net18 net2 VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__o21bai_1
XFILLER_0_9_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_13_Left_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_084_ net21 _040_ net37 VGND VGND VPWR VPWR _005_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_067_ net6 net5 net4 VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__and3_1
X_119_ clknet_1_0__leaf_osc_ck _010_ net22 VGND VGND VPWR VPWR cnt_por\[5\] sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_1_Left_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_083_ net3 net21 VGND VGND VPWR VPWR _040_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_3_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_049_ net1 VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__inv_2
XFILLER_0_10_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_118_ clknet_1_1__leaf_osc_ck _009_ net22 VGND VGND VPWR VPWR cnt_por\[4\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_5_41 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_066_ net4 net5 net6 VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__and3b_1
XPHY_EDGE_ROW_4_Left_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_51 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_082_ _023_ _038_ _039_ VGND VGND VPWR VPWR _004_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_0_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_065_ net5 net4 net6 VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__and3b_1
XFILLER_0_15_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_117_ clknet_1_1__leaf_osc_ck _008_ net22 VGND VGND VPWR VPWR cnt_por\[3\] sky130_fd_sc_hd__dfrtp_1
X_048_ net36 VGND VGND VPWR VPWR _023_ sky130_fd_sc_hd__inv_2
XFILLER_0_10_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_12_52 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_081_ _023_ _038_ _025_ VGND VGND VPWR VPWR _039_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_3_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_064_ net5 net4 net6 VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__nor3b_1
X_116_ clknet_1_1__leaf_osc_ck _007_ net23 VGND VGND VPWR VPWR cnt_por\[2\] sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_080_ cnt_st\[1\] cnt_st\[2\] cnt_st\[3\] net3 VGND VGND VPWR VPWR _038_ sky130_fd_sc_hd__and4_1
XFILLER_0_0_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_063_ net6 net5 net4 VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__and3b_1
XFILLER_0_15_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_115_ clknet_1_1__leaf_osc_ck _006_ net23 VGND VGND VPWR VPWR cnt_por\[1\] sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_8_Left_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
.ends

