magic
tech sky130A
magscale 1 2
timestamp 1713020960
<< viali >>
rect 6469 11305 6503 11339
rect 6101 11237 6135 11271
rect 4169 11101 4203 11135
rect 4353 11101 4387 11135
rect 5825 11101 5859 11135
rect 6653 11101 6687 11135
rect 6101 11033 6135 11067
rect 4261 10965 4295 10999
rect 5917 10965 5951 10999
rect 5841 10761 5875 10795
rect 5641 10693 5675 10727
rect 4813 10625 4847 10659
rect 5090 10625 5124 10659
rect 6377 10625 6411 10659
rect 2789 10557 2823 10591
rect 3065 10557 3099 10591
rect 4905 10557 4939 10591
rect 4997 10557 5031 10591
rect 6653 10557 6687 10591
rect 4629 10489 4663 10523
rect 4537 10421 4571 10455
rect 5825 10421 5859 10455
rect 6009 10421 6043 10455
rect 6469 10421 6503 10455
rect 6561 10421 6595 10455
rect 2605 10217 2639 10251
rect 5089 10217 5123 10251
rect 7573 10081 7607 10115
rect 2789 10013 2823 10047
rect 3065 10013 3099 10047
rect 3341 10013 3375 10047
rect 3617 10013 3651 10047
rect 4077 10013 4111 10047
rect 4169 10013 4203 10047
rect 4537 10013 4571 10047
rect 4629 10013 4663 10047
rect 4813 10013 4847 10047
rect 5181 10013 5215 10047
rect 5457 10013 5491 10047
rect 5549 10013 5583 10047
rect 5825 9945 5859 9979
rect 2973 9877 3007 9911
rect 3157 9877 3191 9911
rect 3525 9877 3559 9911
rect 3893 9877 3927 9911
rect 4353 9877 4387 9911
rect 4445 9877 4479 9911
rect 4537 9673 4571 9707
rect 4997 9673 5031 9707
rect 6193 9673 6227 9707
rect 3065 9605 3099 9639
rect 5089 9605 5123 9639
rect 5273 9605 5307 9639
rect 6653 9605 6687 9639
rect 2789 9537 2823 9571
rect 4905 9537 4939 9571
rect 5825 9537 5859 9571
rect 6377 9537 6411 9571
rect 5549 9469 5583 9503
rect 5733 9469 5767 9503
rect 8125 9469 8159 9503
rect 4721 9401 4755 9435
rect 4353 9129 4387 9163
rect 5273 9129 5307 9163
rect 4261 8993 4295 9027
rect 4629 8925 4663 8959
rect 5089 8925 5123 8959
rect 5243 8925 5277 8959
rect 9505 8925 9539 8959
rect 5549 8857 5583 8891
rect 4445 8789 4479 8823
rect 4537 8789 4571 8823
rect 6837 8789 6871 8823
rect 8953 8789 8987 8823
rect 3985 8585 4019 8619
rect 4829 8585 4863 8619
rect 4997 8585 5031 8619
rect 5549 8585 5583 8619
rect 6101 8585 6135 8619
rect 9597 8585 9631 8619
rect 3157 8517 3191 8551
rect 4353 8517 4387 8551
rect 4629 8517 4663 8551
rect 6561 8517 6595 8551
rect 1409 8449 1443 8483
rect 2973 8449 3007 8483
rect 3249 8449 3283 8483
rect 3341 8449 3375 8483
rect 3525 8449 3559 8483
rect 3801 8449 3835 8483
rect 4252 8471 4286 8505
rect 4537 8449 4571 8483
rect 5089 8449 5123 8483
rect 5181 8449 5215 8483
rect 5825 8449 5859 8483
rect 5917 8449 5951 8483
rect 6101 8449 6135 8483
rect 7113 8449 7147 8483
rect 8953 8449 8987 8483
rect 9130 8449 9164 8483
rect 9221 8449 9255 8483
rect 9413 8439 9447 8473
rect 9505 8449 9539 8483
rect 9689 8449 9723 8483
rect 1961 8381 1995 8415
rect 3617 8381 3651 8415
rect 5365 8381 5399 8415
rect 5549 8381 5583 8415
rect 7389 8381 7423 8415
rect 9045 8381 9079 8415
rect 1593 8313 1627 8347
rect 3433 8313 3467 8347
rect 4537 8313 4571 8347
rect 6377 8313 6411 8347
rect 8861 8313 8895 8347
rect 2789 8245 2823 8279
rect 4813 8245 4847 8279
rect 5273 8245 5307 8279
rect 5733 8245 5767 8279
rect 9321 8245 9355 8279
rect 3341 8041 3375 8075
rect 5089 7973 5123 8007
rect 3157 7905 3191 7939
rect 4353 7905 4387 7939
rect 4537 7905 4571 7939
rect 4721 7905 4755 7939
rect 4813 7905 4847 7939
rect 6561 7905 6595 7939
rect 6837 7905 6871 7939
rect 6929 7905 6963 7939
rect 9689 7905 9723 7939
rect 3249 7837 3283 7871
rect 3341 7837 3375 7871
rect 3617 7837 3651 7871
rect 3801 7837 3835 7871
rect 3985 7837 4019 7871
rect 4169 7837 4203 7871
rect 4261 7837 4295 7871
rect 4629 7837 4663 7871
rect 8953 7837 8987 7871
rect 10057 7837 10091 7871
rect 2881 7769 2915 7803
rect 7205 7769 7239 7803
rect 9873 7769 9907 7803
rect 1409 7701 1443 7735
rect 3433 7701 3467 7735
rect 8677 7701 8711 7735
rect 9597 7701 9631 7735
rect 8953 7497 8987 7531
rect 2789 7429 2823 7463
rect 4353 7429 4387 7463
rect 6377 7361 6411 7395
rect 6561 7361 6595 7395
rect 6653 7361 6687 7395
rect 6929 7361 6963 7395
rect 9137 7361 9171 7395
rect 9229 7361 9263 7395
rect 9413 7361 9447 7395
rect 9505 7361 9539 7395
rect 9873 7361 9907 7395
rect 1593 7293 1627 7327
rect 2513 7293 2547 7327
rect 7205 7293 7239 7327
rect 9597 7293 9631 7327
rect 6377 7225 6411 7259
rect 9689 7225 9723 7259
rect 2237 7157 2271 7191
rect 4261 7157 4295 7191
rect 5825 7157 5859 7191
rect 8677 7157 8711 7191
rect 9781 7157 9815 7191
rect 2040 6953 2074 6987
rect 3525 6953 3559 6987
rect 5825 6953 5859 6987
rect 6285 6953 6319 6987
rect 6653 6953 6687 6987
rect 8607 6953 8641 6987
rect 9597 6953 9631 6987
rect 1501 6885 1535 6919
rect 6101 6885 6135 6919
rect 9505 6885 9539 6919
rect 3801 6817 3835 6851
rect 4261 6817 4295 6851
rect 4721 6817 4755 6851
rect 5181 6817 5215 6851
rect 1685 6749 1719 6783
rect 1777 6749 1811 6783
rect 3985 6749 4019 6783
rect 4077 6749 4111 6783
rect 4169 6749 4203 6783
rect 4813 6749 4847 6783
rect 6929 6749 6963 6783
rect 7113 6749 7147 6783
rect 9137 6749 9171 6783
rect 9321 6749 9355 6783
rect 9597 6749 9631 6783
rect 9873 6749 9907 6783
rect 5779 6715 5813 6749
rect 5457 6681 5491 6715
rect 5983 6681 6017 6715
rect 6469 6681 6503 6715
rect 6745 6681 6779 6715
rect 8401 6681 8435 6715
rect 8617 6681 8651 6715
rect 9781 6681 9815 6715
rect 4445 6613 4479 6647
rect 5641 6613 5675 6647
rect 6269 6613 6303 6647
rect 7021 6613 7055 6647
rect 8769 6613 8803 6647
rect 8953 6613 8987 6647
rect 9229 6613 9263 6647
rect 3709 6409 3743 6443
rect 4445 6409 4479 6443
rect 4721 6409 4755 6443
rect 4905 6409 4939 6443
rect 5825 6409 5859 6443
rect 6377 6409 6411 6443
rect 9321 6409 9355 6443
rect 9965 6409 9999 6443
rect 3617 6341 3651 6375
rect 5365 6341 5399 6375
rect 3433 6273 3467 6307
rect 3709 6273 3743 6307
rect 3893 6273 3927 6307
rect 4537 6273 4571 6307
rect 4629 6273 4663 6307
rect 4905 6273 4939 6307
rect 5273 6273 5307 6307
rect 5457 6273 5491 6307
rect 5825 6273 5859 6307
rect 6101 6273 6135 6307
rect 6561 6273 6595 6307
rect 6653 6273 6687 6307
rect 6745 6273 6779 6307
rect 6837 6273 6871 6307
rect 7021 6273 7055 6307
rect 7941 6273 7975 6307
rect 9137 6273 9171 6307
rect 9689 6273 9723 6307
rect 9781 6273 9815 6307
rect 1409 6205 1443 6239
rect 1685 6205 1719 6239
rect 5733 6205 5767 6239
rect 7665 6205 7699 6239
rect 8953 6205 8987 6239
rect 5917 6137 5951 6171
rect 7757 6137 7791 6171
rect 3157 6069 3191 6103
rect 4997 6069 5031 6103
rect 5641 6069 5675 6103
rect 8125 6069 8159 6103
rect 9505 6069 9539 6103
rect 1409 5865 1443 5899
rect 3433 5865 3467 5899
rect 3525 5865 3559 5899
rect 7205 5865 7239 5899
rect 9045 5865 9079 5899
rect 3341 5729 3375 5763
rect 7021 5729 7055 5763
rect 8033 5729 8067 5763
rect 8677 5729 8711 5763
rect 3157 5661 3191 5695
rect 3617 5661 3651 5695
rect 4077 5661 4111 5695
rect 4169 5661 4203 5695
rect 4261 5661 4295 5695
rect 4445 5661 4479 5695
rect 4537 5661 4571 5695
rect 5273 5661 5307 5695
rect 7113 5661 7147 5695
rect 7573 5661 7607 5695
rect 7665 5661 7699 5695
rect 8953 5661 8987 5695
rect 9229 5661 9263 5695
rect 9505 5661 9539 5695
rect 9689 5661 9723 5695
rect 9965 5661 9999 5695
rect 2881 5593 2915 5627
rect 5549 5593 5583 5627
rect 8125 5593 8159 5627
rect 3801 5525 3835 5559
rect 5181 5525 5215 5559
rect 7389 5525 7423 5559
rect 9413 5525 9447 5559
rect 9873 5525 9907 5559
rect 3985 5321 4019 5355
rect 8493 5321 8527 5355
rect 8769 5321 8803 5355
rect 9873 5321 9907 5355
rect 5825 5253 5859 5287
rect 7021 5253 7055 5287
rect 9689 5253 9723 5287
rect 1777 5185 1811 5219
rect 2145 5185 2179 5219
rect 2237 5185 2271 5219
rect 8585 5185 8619 5219
rect 8769 5185 8803 5219
rect 9505 5185 9539 5219
rect 2513 5117 2547 5151
rect 6745 5117 6779 5151
rect 4537 5049 4571 5083
rect 1593 4981 1627 5015
rect 2053 4981 2087 5015
rect 2237 4777 2271 4811
rect 6009 4777 6043 4811
rect 8769 4777 8803 4811
rect 4261 4641 4295 4675
rect 6745 4641 6779 4675
rect 7021 4641 7055 4675
rect 7297 4641 7331 4675
rect 1807 4573 1841 4607
rect 1961 4573 1995 4607
rect 2053 4573 2087 4607
rect 4537 4505 4571 4539
rect 1593 4437 1627 4471
rect 6101 4437 6135 4471
rect 1501 4233 1535 4267
rect 1777 4233 1811 4267
rect 6469 4165 6503 4199
rect 1685 4097 1719 4131
rect 1961 4097 1995 4131
rect 4077 4097 4111 4131
rect 4721 4097 4755 4131
rect 3985 4029 4019 4063
rect 4445 4029 4479 4063
rect 4813 4029 4847 4063
rect 5089 4029 5123 4063
rect 5733 4029 5767 4063
rect 6653 4029 6687 4063
rect 5181 3961 5215 3995
rect 5825 3621 5859 3655
rect 5917 3621 5951 3655
rect 1685 3485 1719 3519
rect 4997 3485 5031 3519
rect 5089 3485 5123 3519
rect 5181 3485 5215 3519
rect 5641 3485 5675 3519
rect 5917 3485 5951 3519
rect 6009 3485 6043 3519
rect 1501 3349 1535 3383
rect 4813 3349 4847 3383
rect 6193 3349 6227 3383
rect 1869 3145 1903 3179
rect 4215 3145 4249 3179
rect 5549 3145 5583 3179
rect 6193 3145 6227 3179
rect 5365 3077 5399 3111
rect 6009 3077 6043 3111
rect 6561 3077 6595 3111
rect 1409 3009 1443 3043
rect 1777 3009 1811 3043
rect 2973 3009 3007 3043
rect 4997 3009 5031 3043
rect 5641 3009 5675 3043
rect 3249 2941 3283 2975
rect 3341 2941 3375 2975
rect 3433 2941 3467 2975
rect 3985 2941 4019 2975
rect 6929 2941 6963 2975
rect 1593 2873 1627 2907
rect 2789 2805 2823 2839
rect 3617 2805 3651 2839
rect 5365 2805 5399 2839
rect 6009 2805 6043 2839
rect 6377 2805 6411 2839
rect 6561 2805 6595 2839
rect 3157 2601 3191 2635
rect 6009 2601 6043 2635
rect 3341 2465 3375 2499
rect 3433 2465 3467 2499
rect 4905 2465 4939 2499
rect 2053 2397 2087 2431
rect 2329 2397 2363 2431
rect 3525 2397 3559 2431
rect 3801 2397 3835 2431
rect 4537 2397 4571 2431
rect 4629 2397 4663 2431
rect 6561 2397 6595 2431
rect 7205 2397 7239 2431
rect 7849 2397 7883 2431
rect 8493 2397 8527 2431
rect 5825 2329 5859 2363
rect 6025 2329 6059 2363
rect 3985 2261 4019 2295
rect 4353 2261 4387 2295
rect 6193 2261 6227 2295
rect 6745 2261 6779 2295
rect 7389 2261 7423 2295
rect 8033 2261 8067 2295
rect 8677 2261 8711 2295
<< metal1 >>
rect 1104 11450 10396 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 10396 11450
rect 1104 11376 10396 11398
rect 5810 11296 5816 11348
rect 5868 11336 5874 11348
rect 6457 11339 6515 11345
rect 6457 11336 6469 11339
rect 5868 11308 6469 11336
rect 5868 11296 5874 11308
rect 6457 11305 6469 11308
rect 6503 11305 6515 11339
rect 6457 11299 6515 11305
rect 6086 11228 6092 11280
rect 6144 11228 6150 11280
rect 4798 11200 4804 11212
rect 4356 11172 4804 11200
rect 4356 11141 4384 11172
rect 4798 11160 4804 11172
rect 4856 11200 4862 11212
rect 4856 11172 6684 11200
rect 4856 11160 4862 11172
rect 4157 11135 4215 11141
rect 4157 11101 4169 11135
rect 4203 11101 4215 11135
rect 4157 11095 4215 11101
rect 4341 11135 4399 11141
rect 4341 11101 4353 11135
rect 4387 11101 4399 11135
rect 4341 11095 4399 11101
rect 4172 11064 4200 11095
rect 5810 11092 5816 11144
rect 5868 11092 5874 11144
rect 6656 11141 6684 11172
rect 6641 11135 6699 11141
rect 6641 11101 6653 11135
rect 6687 11132 6699 11135
rect 6730 11132 6736 11144
rect 6687 11104 6736 11132
rect 6687 11101 6699 11104
rect 6641 11095 6699 11101
rect 6730 11092 6736 11104
rect 6788 11092 6794 11144
rect 5258 11064 5264 11076
rect 4172 11036 5264 11064
rect 5258 11024 5264 11036
rect 5316 11024 5322 11076
rect 5626 11024 5632 11076
rect 5684 11064 5690 11076
rect 6089 11067 6147 11073
rect 6089 11064 6101 11067
rect 5684 11036 6101 11064
rect 5684 11024 5690 11036
rect 6089 11033 6101 11036
rect 6135 11033 6147 11067
rect 6089 11027 6147 11033
rect 4249 10999 4307 11005
rect 4249 10965 4261 10999
rect 4295 10996 4307 10999
rect 4706 10996 4712 11008
rect 4295 10968 4712 10996
rect 4295 10965 4307 10968
rect 4249 10959 4307 10965
rect 4706 10956 4712 10968
rect 4764 10956 4770 11008
rect 5902 10956 5908 11008
rect 5960 10956 5966 11008
rect 1104 10906 10396 10928
rect 1104 10854 4874 10906
rect 4926 10854 4938 10906
rect 4990 10854 5002 10906
rect 5054 10854 5066 10906
rect 5118 10854 5130 10906
rect 5182 10854 10396 10906
rect 1104 10832 10396 10854
rect 5810 10792 5816 10804
rect 5868 10801 5874 10804
rect 5868 10795 5887 10801
rect 4816 10764 5816 10792
rect 4154 10616 4160 10668
rect 4212 10616 4218 10668
rect 4816 10665 4844 10764
rect 5810 10752 5816 10764
rect 5875 10792 5887 10795
rect 5994 10792 6000 10804
rect 5875 10764 6000 10792
rect 5875 10761 5887 10764
rect 5868 10755 5887 10761
rect 5868 10752 5874 10755
rect 5994 10752 6000 10764
rect 6052 10752 6058 10804
rect 6086 10752 6092 10804
rect 6144 10752 6150 10804
rect 5626 10684 5632 10736
rect 5684 10684 5690 10736
rect 4801 10659 4859 10665
rect 4801 10625 4813 10659
rect 4847 10625 4859 10659
rect 4801 10619 4859 10625
rect 5074 10616 5080 10668
rect 5132 10616 5138 10668
rect 6104 10656 6132 10752
rect 6365 10659 6423 10665
rect 6365 10656 6377 10659
rect 6104 10628 6377 10656
rect 6365 10625 6377 10628
rect 6411 10625 6423 10659
rect 6365 10619 6423 10625
rect 2774 10548 2780 10600
rect 2832 10548 2838 10600
rect 3050 10548 3056 10600
rect 3108 10548 3114 10600
rect 4893 10591 4951 10597
rect 4893 10557 4905 10591
rect 4939 10557 4951 10591
rect 4893 10551 4951 10557
rect 4985 10591 5043 10597
rect 4985 10557 4997 10591
rect 5031 10588 5043 10591
rect 5626 10588 5632 10600
rect 5031 10560 5632 10588
rect 5031 10557 5043 10560
rect 4985 10551 5043 10557
rect 4617 10523 4675 10529
rect 4617 10520 4629 10523
rect 4080 10492 4629 10520
rect 3510 10412 3516 10464
rect 3568 10452 3574 10464
rect 4080 10452 4108 10492
rect 4617 10489 4629 10492
rect 4663 10489 4675 10523
rect 4908 10520 4936 10551
rect 5626 10548 5632 10560
rect 5684 10548 5690 10600
rect 6638 10548 6644 10600
rect 6696 10548 6702 10600
rect 4908 10492 5856 10520
rect 4617 10483 4675 10489
rect 3568 10424 4108 10452
rect 3568 10412 3574 10424
rect 4522 10412 4528 10464
rect 4580 10452 4586 10464
rect 5074 10452 5080 10464
rect 4580 10424 5080 10452
rect 4580 10412 4586 10424
rect 5074 10412 5080 10424
rect 5132 10412 5138 10464
rect 5828 10461 5856 10492
rect 5813 10455 5871 10461
rect 5813 10421 5825 10455
rect 5859 10452 5871 10455
rect 5902 10452 5908 10464
rect 5859 10424 5908 10452
rect 5859 10421 5871 10424
rect 5813 10415 5871 10421
rect 5902 10412 5908 10424
rect 5960 10412 5966 10464
rect 5997 10455 6055 10461
rect 5997 10421 6009 10455
rect 6043 10452 6055 10455
rect 6457 10455 6515 10461
rect 6457 10452 6469 10455
rect 6043 10424 6469 10452
rect 6043 10421 6055 10424
rect 5997 10415 6055 10421
rect 6457 10421 6469 10424
rect 6503 10421 6515 10455
rect 6457 10415 6515 10421
rect 6546 10412 6552 10464
rect 6604 10412 6610 10464
rect 1104 10362 10396 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 10396 10362
rect 1104 10288 10396 10310
rect 2593 10251 2651 10257
rect 2593 10217 2605 10251
rect 2639 10248 2651 10251
rect 3050 10248 3056 10260
rect 2639 10220 3056 10248
rect 2639 10217 2651 10220
rect 2593 10211 2651 10217
rect 3050 10208 3056 10220
rect 3108 10208 3114 10260
rect 4338 10208 4344 10260
rect 4396 10248 4402 10260
rect 4798 10248 4804 10260
rect 4396 10220 4804 10248
rect 4396 10208 4402 10220
rect 4798 10208 4804 10220
rect 4856 10208 4862 10260
rect 5077 10251 5135 10257
rect 5077 10217 5089 10251
rect 5123 10248 5135 10251
rect 6178 10248 6184 10260
rect 5123 10220 6184 10248
rect 5123 10217 5135 10220
rect 5077 10211 5135 10217
rect 6178 10208 6184 10220
rect 6236 10208 6242 10260
rect 2774 10140 2780 10192
rect 2832 10180 2838 10192
rect 5534 10180 5540 10192
rect 2832 10152 5540 10180
rect 2832 10140 2838 10152
rect 5534 10140 5540 10152
rect 5592 10140 5598 10192
rect 3510 10112 3516 10124
rect 3068 10084 3516 10112
rect 3068 10053 3096 10084
rect 3510 10072 3516 10084
rect 3568 10072 3574 10124
rect 4706 10112 4712 10124
rect 3620 10084 4712 10112
rect 3620 10053 3648 10084
rect 4706 10072 4712 10084
rect 4764 10072 4770 10124
rect 5350 10112 5356 10124
rect 5184 10084 5356 10112
rect 2777 10047 2835 10053
rect 2777 10013 2789 10047
rect 2823 10013 2835 10047
rect 2777 10007 2835 10013
rect 3053 10047 3111 10053
rect 3053 10013 3065 10047
rect 3099 10013 3111 10047
rect 3053 10007 3111 10013
rect 3329 10047 3387 10053
rect 3329 10013 3341 10047
rect 3375 10013 3387 10047
rect 3329 10007 3387 10013
rect 3605 10047 3663 10053
rect 3605 10013 3617 10047
rect 3651 10013 3663 10047
rect 3605 10007 3663 10013
rect 4065 10047 4123 10053
rect 4065 10013 4077 10047
rect 4111 10013 4123 10047
rect 4065 10007 4123 10013
rect 4157 10047 4215 10053
rect 4157 10013 4169 10047
rect 4203 10044 4215 10047
rect 4246 10044 4252 10056
rect 4203 10016 4252 10044
rect 4203 10013 4215 10016
rect 4157 10007 4215 10013
rect 2792 9976 2820 10007
rect 2866 9976 2872 9988
rect 2792 9948 2872 9976
rect 2866 9936 2872 9948
rect 2924 9976 2930 9988
rect 3344 9976 3372 10007
rect 2924 9948 3372 9976
rect 4080 9976 4108 10007
rect 4246 10004 4252 10016
rect 4304 10004 4310 10056
rect 4338 10004 4344 10056
rect 4396 10044 4402 10056
rect 4525 10047 4583 10053
rect 4525 10044 4537 10047
rect 4396 10016 4537 10044
rect 4396 10004 4402 10016
rect 4525 10013 4537 10016
rect 4571 10013 4583 10047
rect 4525 10007 4583 10013
rect 4614 10004 4620 10056
rect 4672 10004 4678 10056
rect 5184 10053 5212 10084
rect 5350 10072 5356 10084
rect 5408 10112 5414 10124
rect 5902 10112 5908 10124
rect 5408 10084 5908 10112
rect 5408 10072 5414 10084
rect 5902 10072 5908 10084
rect 5960 10112 5966 10124
rect 7561 10115 7619 10121
rect 7561 10112 7573 10115
rect 5960 10084 7573 10112
rect 5960 10072 5966 10084
rect 7561 10081 7573 10084
rect 7607 10081 7619 10115
rect 7561 10075 7619 10081
rect 4801 10047 4859 10053
rect 4801 10013 4813 10047
rect 4847 10013 4859 10047
rect 4801 10007 4859 10013
rect 5169 10047 5227 10053
rect 5169 10013 5181 10047
rect 5215 10013 5227 10047
rect 5169 10007 5227 10013
rect 5445 10047 5503 10053
rect 5445 10013 5457 10047
rect 5491 10013 5503 10047
rect 5445 10007 5503 10013
rect 4816 9976 4844 10007
rect 4080 9948 4844 9976
rect 2924 9936 2930 9948
rect 4540 9920 4568 9948
rect 2958 9868 2964 9920
rect 3016 9868 3022 9920
rect 3142 9868 3148 9920
rect 3200 9868 3206 9920
rect 3513 9911 3571 9917
rect 3513 9877 3525 9911
rect 3559 9908 3571 9911
rect 3881 9911 3939 9917
rect 3881 9908 3893 9911
rect 3559 9880 3893 9908
rect 3559 9877 3571 9880
rect 3513 9871 3571 9877
rect 3881 9877 3893 9880
rect 3927 9877 3939 9911
rect 3881 9871 3939 9877
rect 4338 9868 4344 9920
rect 4396 9868 4402 9920
rect 4430 9868 4436 9920
rect 4488 9868 4494 9920
rect 4522 9868 4528 9920
rect 4580 9868 4586 9920
rect 5460 9908 5488 10007
rect 5534 10004 5540 10056
rect 5592 10004 5598 10056
rect 6914 10004 6920 10056
rect 6972 10004 6978 10056
rect 5810 9936 5816 9988
rect 5868 9936 5874 9988
rect 5902 9936 5908 9988
rect 5960 9936 5966 9988
rect 5626 9908 5632 9920
rect 5460 9880 5632 9908
rect 5626 9868 5632 9880
rect 5684 9908 5690 9920
rect 5920 9908 5948 9936
rect 5684 9880 5948 9908
rect 5684 9868 5690 9880
rect 1104 9818 10396 9840
rect 1104 9766 4874 9818
rect 4926 9766 4938 9818
rect 4990 9766 5002 9818
rect 5054 9766 5066 9818
rect 5118 9766 5130 9818
rect 5182 9766 10396 9818
rect 1104 9744 10396 9766
rect 4522 9664 4528 9716
rect 4580 9704 4586 9716
rect 4985 9707 5043 9713
rect 4985 9704 4997 9707
rect 4580 9676 4997 9704
rect 4580 9664 4586 9676
rect 4985 9673 4997 9676
rect 5031 9673 5043 9707
rect 4985 9667 5043 9673
rect 5350 9664 5356 9716
rect 5408 9664 5414 9716
rect 5810 9664 5816 9716
rect 5868 9704 5874 9716
rect 6181 9707 6239 9713
rect 6181 9704 6193 9707
rect 5868 9676 6193 9704
rect 5868 9664 5874 9676
rect 6181 9673 6193 9676
rect 6227 9673 6239 9707
rect 6181 9667 6239 9673
rect 7006 9664 7012 9716
rect 7064 9664 7070 9716
rect 3053 9639 3111 9645
rect 3053 9605 3065 9639
rect 3099 9636 3111 9639
rect 3142 9636 3148 9648
rect 3099 9608 3148 9636
rect 3099 9605 3111 9608
rect 3053 9599 3111 9605
rect 3142 9596 3148 9608
rect 3200 9596 3206 9648
rect 4614 9596 4620 9648
rect 4672 9636 4678 9648
rect 5077 9639 5135 9645
rect 5077 9636 5089 9639
rect 4672 9608 5089 9636
rect 4672 9596 4678 9608
rect 5077 9605 5089 9608
rect 5123 9605 5135 9639
rect 5077 9599 5135 9605
rect 5258 9596 5264 9648
rect 5316 9596 5322 9648
rect 2774 9528 2780 9580
rect 2832 9528 2838 9580
rect 4154 9528 4160 9580
rect 4212 9528 4218 9580
rect 4338 9528 4344 9580
rect 4396 9568 4402 9580
rect 4893 9571 4951 9577
rect 4893 9568 4905 9571
rect 4396 9540 4905 9568
rect 4396 9528 4402 9540
rect 4893 9537 4905 9540
rect 4939 9568 4951 9571
rect 5368 9568 5396 9664
rect 5534 9596 5540 9648
rect 5592 9636 5598 9648
rect 5592 9608 6408 9636
rect 5592 9596 5598 9608
rect 6380 9580 6408 9608
rect 6546 9596 6552 9648
rect 6604 9636 6610 9648
rect 6641 9639 6699 9645
rect 6641 9636 6653 9639
rect 6604 9608 6653 9636
rect 6604 9596 6610 9608
rect 6641 9605 6653 9608
rect 6687 9605 6699 9639
rect 7024 9636 7052 9664
rect 7024 9608 7130 9636
rect 6641 9599 6699 9605
rect 5813 9571 5871 9577
rect 4939 9540 5580 9568
rect 4939 9537 4951 9540
rect 4893 9531 4951 9537
rect 4172 9364 4200 9528
rect 5552 9509 5580 9540
rect 5813 9537 5825 9571
rect 5859 9568 5871 9571
rect 5994 9568 6000 9580
rect 5859 9540 6000 9568
rect 5859 9537 5871 9540
rect 5813 9531 5871 9537
rect 5994 9528 6000 9540
rect 6052 9528 6058 9580
rect 6362 9528 6368 9580
rect 6420 9528 6426 9580
rect 5537 9503 5595 9509
rect 5537 9469 5549 9503
rect 5583 9500 5595 9503
rect 5626 9500 5632 9512
rect 5583 9472 5632 9500
rect 5583 9469 5595 9472
rect 5537 9463 5595 9469
rect 5626 9460 5632 9472
rect 5684 9460 5690 9512
rect 5718 9460 5724 9512
rect 5776 9460 5782 9512
rect 5902 9460 5908 9512
rect 5960 9500 5966 9512
rect 8113 9503 8171 9509
rect 8113 9500 8125 9503
rect 5960 9472 8125 9500
rect 5960 9460 5966 9472
rect 8113 9469 8125 9472
rect 8159 9469 8171 9503
rect 8113 9463 8171 9469
rect 4246 9392 4252 9444
rect 4304 9432 4310 9444
rect 4709 9435 4767 9441
rect 4709 9432 4721 9435
rect 4304 9404 4721 9432
rect 4304 9392 4310 9404
rect 4709 9401 4721 9404
rect 4755 9432 4767 9435
rect 5920 9432 5948 9460
rect 4755 9404 5948 9432
rect 4755 9401 4767 9404
rect 4709 9395 4767 9401
rect 5442 9364 5448 9376
rect 4172 9336 5448 9364
rect 5442 9324 5448 9336
rect 5500 9364 5506 9376
rect 7006 9364 7012 9376
rect 5500 9336 7012 9364
rect 5500 9324 5506 9336
rect 7006 9324 7012 9336
rect 7064 9324 7070 9376
rect 1104 9274 10396 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 10396 9274
rect 1104 9200 10396 9222
rect 2958 9120 2964 9172
rect 3016 9160 3022 9172
rect 4341 9163 4399 9169
rect 4341 9160 4353 9163
rect 3016 9132 4353 9160
rect 3016 9120 3022 9132
rect 4341 9129 4353 9132
rect 4387 9129 4399 9163
rect 4341 9123 4399 9129
rect 5261 9163 5319 9169
rect 5261 9129 5273 9163
rect 5307 9160 5319 9163
rect 5718 9160 5724 9172
rect 5307 9132 5724 9160
rect 5307 9129 5319 9132
rect 5261 9123 5319 9129
rect 5718 9120 5724 9132
rect 5776 9120 5782 9172
rect 4632 9064 5488 9092
rect 4154 8984 4160 9036
rect 4212 9024 4218 9036
rect 4249 9027 4307 9033
rect 4249 9024 4261 9027
rect 4212 8996 4261 9024
rect 4212 8984 4218 8996
rect 4249 8993 4261 8996
rect 4295 8993 4307 9027
rect 4249 8987 4307 8993
rect 4632 8965 4660 9064
rect 5350 9024 5356 9036
rect 5099 8996 5356 9024
rect 5099 8966 5127 8996
rect 5350 8984 5356 8996
rect 5408 8984 5414 9036
rect 5092 8965 5127 8966
rect 4617 8959 4675 8965
rect 4617 8925 4629 8959
rect 4663 8925 4675 8959
rect 4617 8919 4675 8925
rect 5077 8959 5135 8965
rect 5077 8925 5089 8959
rect 5123 8925 5135 8959
rect 5077 8919 5135 8925
rect 5231 8959 5289 8965
rect 5231 8925 5243 8959
rect 5277 8956 5289 8959
rect 5460 8956 5488 9064
rect 5994 8956 6000 8968
rect 5277 8928 6000 8956
rect 5277 8925 5289 8928
rect 5231 8919 5289 8925
rect 5994 8916 6000 8928
rect 6052 8916 6058 8968
rect 9398 8916 9404 8968
rect 9456 8956 9462 8968
rect 9493 8959 9551 8965
rect 9493 8956 9505 8959
rect 9456 8928 9505 8956
rect 9456 8916 9462 8928
rect 9493 8925 9505 8928
rect 9539 8925 9551 8959
rect 9493 8919 9551 8925
rect 5537 8891 5595 8897
rect 4448 8860 5396 8888
rect 4448 8829 4476 8860
rect 4433 8823 4491 8829
rect 4433 8789 4445 8823
rect 4479 8789 4491 8823
rect 4433 8783 4491 8789
rect 4525 8823 4583 8829
rect 4525 8789 4537 8823
rect 4571 8820 4583 8823
rect 4614 8820 4620 8832
rect 4571 8792 4620 8820
rect 4571 8789 4583 8792
rect 4525 8783 4583 8789
rect 4614 8780 4620 8792
rect 4672 8780 4678 8832
rect 5368 8820 5396 8860
rect 5537 8857 5549 8891
rect 5583 8888 5595 8891
rect 5810 8888 5816 8900
rect 5583 8860 5816 8888
rect 5583 8857 5595 8860
rect 5537 8851 5595 8857
rect 5810 8848 5816 8860
rect 5868 8848 5874 8900
rect 5626 8820 5632 8832
rect 5368 8792 5632 8820
rect 5626 8780 5632 8792
rect 5684 8780 5690 8832
rect 6362 8780 6368 8832
rect 6420 8820 6426 8832
rect 6822 8820 6828 8832
rect 6420 8792 6828 8820
rect 6420 8780 6426 8792
rect 6822 8780 6828 8792
rect 6880 8780 6886 8832
rect 8938 8780 8944 8832
rect 8996 8780 9002 8832
rect 1104 8730 10396 8752
rect 1104 8678 4874 8730
rect 4926 8678 4938 8730
rect 4990 8678 5002 8730
rect 5054 8678 5066 8730
rect 5118 8678 5130 8730
rect 5182 8678 10396 8730
rect 1104 8656 10396 8678
rect 3970 8616 3976 8628
rect 2976 8588 3976 8616
rect 1394 8440 1400 8492
rect 1452 8440 1458 8492
rect 2866 8440 2872 8492
rect 2924 8480 2930 8492
rect 2976 8489 3004 8588
rect 3970 8576 3976 8588
rect 4028 8576 4034 8628
rect 4817 8619 4875 8625
rect 4817 8616 4829 8619
rect 4218 8588 4829 8616
rect 3145 8551 3203 8557
rect 3145 8517 3157 8551
rect 3191 8548 3203 8551
rect 3418 8548 3424 8560
rect 3191 8520 3424 8548
rect 3191 8517 3203 8520
rect 3145 8511 3203 8517
rect 3418 8508 3424 8520
rect 3476 8508 3482 8560
rect 4218 8548 4246 8588
rect 4817 8585 4829 8588
rect 4863 8585 4875 8619
rect 4817 8579 4875 8585
rect 4985 8619 5043 8625
rect 4985 8585 4997 8619
rect 5031 8585 5043 8619
rect 4985 8579 5043 8585
rect 3896 8520 4246 8548
rect 3896 8492 3924 8520
rect 4218 8511 4246 8520
rect 4341 8551 4399 8557
rect 4341 8517 4353 8551
rect 4387 8517 4399 8551
rect 4341 8511 4399 8517
rect 4617 8551 4675 8557
rect 4617 8517 4629 8551
rect 4663 8548 4675 8551
rect 5000 8548 5028 8579
rect 5534 8576 5540 8628
rect 5592 8576 5598 8628
rect 6089 8619 6147 8625
rect 6089 8585 6101 8619
rect 6135 8616 6147 8619
rect 6638 8616 6644 8628
rect 6135 8588 6644 8616
rect 6135 8585 6147 8588
rect 6089 8579 6147 8585
rect 6104 8548 6132 8579
rect 6638 8576 6644 8588
rect 6696 8576 6702 8628
rect 8938 8576 8944 8628
rect 8996 8576 9002 8628
rect 9585 8619 9643 8625
rect 9585 8616 9597 8619
rect 9048 8588 9597 8616
rect 6549 8551 6607 8557
rect 6549 8548 6561 8551
rect 4663 8520 4752 8548
rect 5000 8520 5212 8548
rect 4663 8517 4675 8520
rect 4617 8511 4675 8517
rect 4218 8505 4298 8511
rect 2961 8483 3019 8489
rect 2961 8480 2973 8483
rect 2924 8452 2973 8480
rect 2924 8440 2930 8452
rect 2961 8449 2973 8452
rect 3007 8449 3019 8483
rect 2961 8443 3019 8449
rect 3234 8440 3240 8492
rect 3292 8440 3298 8492
rect 3329 8483 3387 8489
rect 3329 8449 3341 8483
rect 3375 8449 3387 8483
rect 3329 8443 3387 8449
rect 1949 8415 2007 8421
rect 1949 8381 1961 8415
rect 1995 8412 2007 8415
rect 1995 8384 2774 8412
rect 1995 8381 2007 8384
rect 1949 8375 2007 8381
rect 1581 8347 1639 8353
rect 1581 8313 1593 8347
rect 1627 8344 1639 8347
rect 1670 8344 1676 8356
rect 1627 8316 1676 8344
rect 1627 8313 1639 8316
rect 1581 8307 1639 8313
rect 1670 8304 1676 8316
rect 1728 8304 1734 8356
rect 2746 8344 2774 8384
rect 2958 8344 2964 8356
rect 2746 8316 2964 8344
rect 2958 8304 2964 8316
rect 3016 8304 3022 8356
rect 2777 8279 2835 8285
rect 2777 8245 2789 8279
rect 2823 8276 2835 8279
rect 2866 8276 2872 8288
rect 2823 8248 2872 8276
rect 2823 8245 2835 8248
rect 2777 8239 2835 8245
rect 2866 8236 2872 8248
rect 2924 8236 2930 8288
rect 3344 8276 3372 8443
rect 3510 8440 3516 8492
rect 3568 8480 3574 8492
rect 3789 8483 3847 8489
rect 3789 8480 3801 8483
rect 3568 8452 3801 8480
rect 3568 8440 3574 8452
rect 3789 8449 3801 8452
rect 3835 8449 3847 8483
rect 3789 8443 3847 8449
rect 3602 8372 3608 8424
rect 3660 8372 3666 8424
rect 3804 8412 3832 8443
rect 3878 8440 3884 8492
rect 3936 8440 3942 8492
rect 4218 8474 4252 8505
rect 4240 8471 4252 8474
rect 4286 8471 4298 8505
rect 4240 8465 4298 8471
rect 4356 8412 4384 8511
rect 4525 8483 4583 8489
rect 4525 8449 4537 8483
rect 4571 8480 4583 8483
rect 4724 8480 4752 8520
rect 4890 8480 4896 8492
rect 4571 8452 4896 8480
rect 4571 8449 4583 8452
rect 4525 8443 4583 8449
rect 4890 8440 4896 8452
rect 4948 8440 4954 8492
rect 5184 8489 5212 8520
rect 5552 8520 6132 8548
rect 6196 8520 6561 8548
rect 5077 8483 5135 8489
rect 5077 8449 5089 8483
rect 5123 8449 5135 8483
rect 5077 8443 5135 8449
rect 5169 8483 5227 8489
rect 5169 8449 5181 8483
rect 5215 8449 5227 8483
rect 5169 8443 5227 8449
rect 5092 8412 5120 8443
rect 5552 8421 5580 8520
rect 5626 8440 5632 8492
rect 5684 8480 5690 8492
rect 5813 8483 5871 8489
rect 5813 8480 5825 8483
rect 5684 8452 5825 8480
rect 5684 8440 5690 8452
rect 5813 8449 5825 8452
rect 5859 8449 5871 8483
rect 5813 8443 5871 8449
rect 5905 8483 5963 8489
rect 5905 8449 5917 8483
rect 5951 8449 5963 8483
rect 5905 8443 5963 8449
rect 3804 8384 4384 8412
rect 4540 8384 5120 8412
rect 5353 8415 5411 8421
rect 3421 8347 3479 8353
rect 3421 8313 3433 8347
rect 3467 8344 3479 8347
rect 4062 8344 4068 8356
rect 3467 8316 4068 8344
rect 3467 8313 3479 8316
rect 3421 8307 3479 8313
rect 4062 8304 4068 8316
rect 4120 8304 4126 8356
rect 3878 8276 3884 8288
rect 3344 8248 3884 8276
rect 3878 8236 3884 8248
rect 3936 8236 3942 8288
rect 4264 8276 4292 8384
rect 4540 8353 4568 8384
rect 5353 8381 5365 8415
rect 5399 8412 5411 8415
rect 5537 8415 5595 8421
rect 5537 8412 5549 8415
rect 5399 8384 5549 8412
rect 5399 8381 5411 8384
rect 5353 8375 5411 8381
rect 5537 8381 5549 8384
rect 5583 8381 5595 8415
rect 5537 8375 5595 8381
rect 4525 8347 4583 8353
rect 4525 8313 4537 8347
rect 4571 8313 4583 8347
rect 5920 8344 5948 8443
rect 5994 8440 6000 8492
rect 6052 8440 6058 8492
rect 6086 8440 6092 8492
rect 6144 8440 6150 8492
rect 6012 8412 6040 8440
rect 6196 8412 6224 8520
rect 6549 8517 6561 8520
rect 6595 8517 6607 8551
rect 6549 8511 6607 8517
rect 8386 8508 8392 8560
rect 8444 8508 8450 8560
rect 6822 8440 6828 8492
rect 6880 8480 6886 8492
rect 8956 8489 8984 8576
rect 9048 8560 9076 8588
rect 9585 8585 9597 8588
rect 9631 8585 9643 8619
rect 9585 8579 9643 8585
rect 9030 8508 9036 8560
rect 9088 8508 9094 8560
rect 9398 8508 9404 8560
rect 9456 8508 9462 8560
rect 7101 8483 7159 8489
rect 7101 8480 7113 8483
rect 6880 8452 7113 8480
rect 6880 8440 6886 8452
rect 7101 8449 7113 8452
rect 7147 8449 7159 8483
rect 7101 8443 7159 8449
rect 8941 8483 8999 8489
rect 8941 8449 8953 8483
rect 8987 8449 8999 8483
rect 9048 8480 9076 8508
rect 9214 8489 9220 8492
rect 9118 8483 9176 8489
rect 9118 8480 9130 8483
rect 9048 8452 9130 8480
rect 8941 8443 8999 8449
rect 9118 8449 9130 8452
rect 9164 8449 9176 8483
rect 9118 8443 9176 8449
rect 9209 8443 9220 8489
rect 9272 8480 9278 8492
rect 9272 8452 9309 8480
rect 9416 8479 9444 8508
rect 9401 8473 9459 8479
rect 9214 8440 9220 8443
rect 9272 8440 9278 8452
rect 9401 8439 9413 8473
rect 9447 8439 9459 8473
rect 9490 8440 9496 8492
rect 9548 8440 9554 8492
rect 9674 8440 9680 8492
rect 9732 8440 9738 8492
rect 9401 8433 9459 8439
rect 6012 8384 6224 8412
rect 7377 8415 7435 8421
rect 7377 8381 7389 8415
rect 7423 8412 7435 8415
rect 9033 8415 9091 8421
rect 9033 8412 9045 8415
rect 7423 8384 9045 8412
rect 7423 8381 7435 8384
rect 7377 8375 7435 8381
rect 9033 8381 9045 8384
rect 9079 8381 9091 8415
rect 9033 8375 9091 8381
rect 6365 8347 6423 8353
rect 6365 8344 6377 8347
rect 4525 8307 4583 8313
rect 4816 8316 6377 8344
rect 4816 8288 4844 8316
rect 6365 8313 6377 8316
rect 6411 8313 6423 8347
rect 6365 8307 6423 8313
rect 8478 8304 8484 8356
rect 8536 8344 8542 8356
rect 8849 8347 8907 8353
rect 8849 8344 8861 8347
rect 8536 8316 8861 8344
rect 8536 8304 8542 8316
rect 8849 8313 8861 8316
rect 8895 8344 8907 8347
rect 9416 8344 9444 8433
rect 8895 8316 9444 8344
rect 8895 8313 8907 8316
rect 8849 8307 8907 8313
rect 4798 8276 4804 8288
rect 4264 8248 4804 8276
rect 4798 8236 4804 8248
rect 4856 8236 4862 8288
rect 5258 8236 5264 8288
rect 5316 8236 5322 8288
rect 5718 8236 5724 8288
rect 5776 8236 5782 8288
rect 9306 8236 9312 8288
rect 9364 8236 9370 8288
rect 1104 8186 10396 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 10396 8186
rect 1104 8112 10396 8134
rect 3234 8032 3240 8084
rect 3292 8072 3298 8084
rect 3329 8075 3387 8081
rect 3329 8072 3341 8075
rect 3292 8044 3341 8072
rect 3292 8032 3298 8044
rect 3329 8041 3341 8044
rect 3375 8041 3387 8075
rect 4798 8072 4804 8084
rect 3329 8035 3387 8041
rect 4540 8044 4804 8072
rect 2774 7896 2780 7948
rect 2832 7936 2838 7948
rect 3145 7939 3203 7945
rect 3145 7936 3157 7939
rect 2832 7908 3157 7936
rect 2832 7896 2838 7908
rect 3145 7905 3157 7908
rect 3191 7905 3203 7939
rect 3878 7936 3884 7948
rect 3145 7899 3203 7905
rect 3252 7908 3884 7936
rect 3252 7877 3280 7908
rect 3878 7896 3884 7908
rect 3936 7896 3942 7948
rect 4540 7945 4568 8044
rect 4798 8032 4804 8044
rect 4856 8032 4862 8084
rect 5534 8032 5540 8084
rect 5592 8032 5598 8084
rect 4614 7964 4620 8016
rect 4672 8004 4678 8016
rect 5077 8007 5135 8013
rect 5077 8004 5089 8007
rect 4672 7976 5089 8004
rect 4672 7964 4678 7976
rect 4724 7945 4752 7976
rect 5077 7973 5089 7976
rect 5123 7973 5135 8007
rect 5077 7967 5135 7973
rect 4341 7939 4399 7945
rect 4341 7905 4353 7939
rect 4387 7905 4399 7939
rect 4341 7899 4399 7905
rect 4525 7939 4583 7945
rect 4525 7905 4537 7939
rect 4571 7905 4583 7939
rect 4525 7899 4583 7905
rect 4709 7939 4767 7945
rect 4709 7905 4721 7939
rect 4755 7905 4767 7939
rect 4709 7899 4767 7905
rect 3237 7871 3295 7877
rect 3237 7837 3249 7871
rect 3283 7837 3295 7871
rect 3237 7831 3295 7837
rect 3329 7871 3387 7877
rect 3329 7837 3341 7871
rect 3375 7868 3387 7871
rect 3510 7868 3516 7880
rect 3375 7840 3516 7868
rect 3375 7837 3387 7840
rect 3329 7831 3387 7837
rect 3510 7828 3516 7840
rect 3568 7828 3574 7880
rect 3602 7828 3608 7880
rect 3660 7828 3666 7880
rect 3786 7828 3792 7880
rect 3844 7828 3850 7880
rect 3970 7828 3976 7880
rect 4028 7828 4034 7880
rect 4154 7828 4160 7880
rect 4212 7828 4218 7880
rect 4249 7871 4307 7877
rect 4249 7837 4261 7871
rect 4295 7868 4307 7871
rect 4356 7868 4384 7899
rect 4798 7896 4804 7948
rect 4856 7896 4862 7948
rect 5166 7896 5172 7948
rect 5224 7936 5230 7948
rect 5350 7936 5356 7948
rect 5224 7908 5356 7936
rect 5224 7896 5230 7908
rect 5350 7896 5356 7908
rect 5408 7896 5414 7948
rect 5552 7936 5580 8032
rect 6549 7939 6607 7945
rect 6549 7936 6561 7939
rect 5552 7908 6561 7936
rect 6549 7905 6561 7908
rect 6595 7905 6607 7939
rect 6549 7899 6607 7905
rect 6822 7896 6828 7948
rect 6880 7936 6886 7948
rect 6917 7939 6975 7945
rect 6917 7936 6929 7939
rect 6880 7908 6929 7936
rect 6880 7896 6886 7908
rect 6917 7905 6929 7908
rect 6963 7905 6975 7939
rect 6917 7899 6975 7905
rect 8386 7896 8392 7948
rect 8444 7896 8450 7948
rect 9122 7896 9128 7948
rect 9180 7936 9186 7948
rect 9677 7939 9735 7945
rect 9677 7936 9689 7939
rect 9180 7908 9689 7936
rect 9180 7896 9186 7908
rect 9677 7905 9689 7908
rect 9723 7905 9735 7939
rect 9677 7899 9735 7905
rect 4295 7840 4384 7868
rect 4617 7871 4675 7877
rect 4295 7837 4307 7840
rect 4249 7831 4307 7837
rect 4617 7837 4629 7871
rect 4663 7868 4675 7871
rect 5184 7868 5212 7896
rect 4663 7840 5212 7868
rect 4663 7837 4675 7840
rect 4617 7831 4675 7837
rect 5258 7828 5264 7880
rect 5316 7828 5322 7880
rect 5442 7828 5448 7880
rect 5500 7828 5506 7880
rect 8404 7868 8432 7896
rect 8326 7840 8432 7868
rect 8938 7828 8944 7880
rect 8996 7828 9002 7880
rect 9398 7828 9404 7880
rect 9456 7868 9462 7880
rect 10045 7871 10103 7877
rect 10045 7868 10057 7871
rect 9456 7840 10057 7868
rect 9456 7828 9462 7840
rect 10045 7837 10057 7840
rect 10091 7837 10103 7871
rect 10045 7831 10103 7837
rect 2774 7800 2780 7812
rect 2438 7772 2780 7800
rect 2774 7760 2780 7772
rect 2832 7760 2838 7812
rect 2869 7803 2927 7809
rect 2869 7769 2881 7803
rect 2915 7800 2927 7803
rect 5276 7800 5304 7828
rect 2915 7772 5304 7800
rect 2915 7769 2927 7772
rect 2869 7763 2927 7769
rect 1397 7735 1455 7741
rect 1397 7701 1409 7735
rect 1443 7732 1455 7735
rect 3421 7735 3479 7741
rect 3421 7732 3433 7735
rect 1443 7704 3433 7732
rect 1443 7701 1455 7704
rect 1397 7695 1455 7701
rect 3421 7701 3433 7704
rect 3467 7732 3479 7735
rect 4062 7732 4068 7744
rect 3467 7704 4068 7732
rect 3467 7701 3479 7704
rect 3421 7695 3479 7701
rect 4062 7692 4068 7704
rect 4120 7732 4126 7744
rect 4890 7732 4896 7744
rect 4120 7704 4896 7732
rect 4120 7692 4126 7704
rect 4890 7692 4896 7704
rect 4948 7692 4954 7744
rect 5258 7692 5264 7744
rect 5316 7732 5322 7744
rect 5460 7732 5488 7828
rect 7190 7760 7196 7812
rect 7248 7760 7254 7812
rect 9214 7800 9220 7812
rect 8680 7772 9220 7800
rect 8680 7744 8708 7772
rect 9214 7760 9220 7772
rect 9272 7800 9278 7812
rect 9861 7803 9919 7809
rect 9861 7800 9873 7803
rect 9272 7772 9873 7800
rect 9272 7760 9278 7772
rect 9861 7769 9873 7772
rect 9907 7769 9919 7803
rect 9861 7763 9919 7769
rect 5316 7704 5488 7732
rect 5316 7692 5322 7704
rect 8662 7692 8668 7744
rect 8720 7692 8726 7744
rect 9582 7692 9588 7744
rect 9640 7692 9646 7744
rect 1104 7642 10396 7664
rect 1104 7590 4874 7642
rect 4926 7590 4938 7642
rect 4990 7590 5002 7642
rect 5054 7590 5066 7642
rect 5118 7590 5130 7642
rect 5182 7590 10396 7642
rect 1104 7568 10396 7590
rect 3786 7528 3792 7540
rect 2792 7500 3792 7528
rect 2792 7469 2820 7500
rect 3786 7488 3792 7500
rect 3844 7488 3850 7540
rect 5994 7488 6000 7540
rect 6052 7528 6058 7540
rect 6546 7528 6552 7540
rect 6052 7500 6552 7528
rect 6052 7488 6058 7500
rect 6546 7488 6552 7500
rect 6604 7528 6610 7540
rect 6604 7500 6684 7528
rect 6604 7488 6610 7500
rect 2777 7463 2835 7469
rect 2777 7429 2789 7463
rect 2823 7429 2835 7463
rect 2777 7423 2835 7429
rect 3050 7420 3056 7472
rect 3108 7460 3114 7472
rect 4341 7463 4399 7469
rect 3108 7432 3266 7460
rect 3108 7420 3114 7432
rect 4341 7429 4353 7463
rect 4387 7460 4399 7463
rect 4706 7460 4712 7472
rect 4387 7432 4712 7460
rect 4387 7429 4399 7432
rect 4341 7423 4399 7429
rect 4706 7420 4712 7432
rect 4764 7420 4770 7472
rect 5350 7420 5356 7472
rect 5408 7460 5414 7472
rect 5408 7432 6500 7460
rect 5408 7420 5414 7432
rect 6472 7404 6500 7432
rect 4614 7352 4620 7404
rect 4672 7392 4678 7404
rect 5994 7392 6000 7404
rect 4672 7364 6000 7392
rect 4672 7352 4678 7364
rect 5994 7352 6000 7364
rect 6052 7392 6058 7404
rect 6365 7395 6423 7401
rect 6365 7392 6377 7395
rect 6052 7364 6377 7392
rect 6052 7352 6058 7364
rect 6365 7361 6377 7364
rect 6411 7361 6423 7395
rect 6365 7355 6423 7361
rect 6454 7352 6460 7404
rect 6512 7392 6518 7404
rect 6656 7401 6684 7500
rect 7006 7488 7012 7540
rect 7064 7488 7070 7540
rect 7190 7488 7196 7540
rect 7248 7528 7254 7540
rect 8941 7531 8999 7537
rect 8941 7528 8953 7531
rect 7248 7500 8953 7528
rect 7248 7488 7254 7500
rect 8941 7497 8953 7500
rect 8987 7497 8999 7531
rect 9122 7528 9128 7540
rect 8941 7491 8999 7497
rect 9048 7500 9128 7528
rect 7024 7460 7052 7488
rect 7024 7432 7682 7460
rect 6549 7395 6607 7401
rect 6549 7392 6561 7395
rect 6512 7364 6561 7392
rect 6512 7352 6518 7364
rect 6549 7361 6561 7364
rect 6595 7361 6607 7395
rect 6549 7355 6607 7361
rect 6641 7395 6699 7401
rect 6641 7361 6653 7395
rect 6687 7361 6699 7395
rect 6641 7355 6699 7361
rect 6822 7352 6828 7404
rect 6880 7392 6886 7404
rect 6917 7395 6975 7401
rect 6917 7392 6929 7395
rect 6880 7364 6929 7392
rect 6880 7352 6886 7364
rect 6917 7361 6929 7364
rect 6963 7361 6975 7395
rect 9048 7392 9076 7500
rect 9122 7488 9128 7500
rect 9180 7488 9186 7540
rect 9674 7528 9680 7540
rect 9416 7500 9680 7528
rect 9125 7395 9183 7401
rect 9125 7392 9137 7395
rect 9048 7364 9137 7392
rect 6917 7355 6975 7361
rect 9125 7361 9137 7364
rect 9171 7361 9183 7395
rect 9125 7355 9183 7361
rect 9217 7395 9275 7401
rect 9217 7361 9229 7395
rect 9263 7392 9275 7395
rect 9306 7392 9312 7404
rect 9263 7364 9312 7392
rect 9263 7361 9275 7364
rect 9217 7355 9275 7361
rect 9306 7352 9312 7364
rect 9364 7352 9370 7404
rect 9416 7401 9444 7500
rect 9674 7488 9680 7500
rect 9732 7488 9738 7540
rect 9401 7395 9459 7401
rect 9401 7361 9413 7395
rect 9447 7361 9459 7395
rect 9401 7355 9459 7361
rect 9490 7352 9496 7404
rect 9548 7352 9554 7404
rect 9858 7352 9864 7404
rect 9916 7352 9922 7404
rect 1578 7284 1584 7336
rect 1636 7284 1642 7336
rect 1762 7284 1768 7336
rect 1820 7324 1826 7336
rect 2501 7327 2559 7333
rect 2501 7324 2513 7327
rect 1820 7296 2513 7324
rect 1820 7284 1826 7296
rect 2501 7293 2513 7296
rect 2547 7293 2559 7327
rect 2501 7287 2559 7293
rect 2774 7284 2780 7336
rect 2832 7324 2838 7336
rect 3142 7324 3148 7336
rect 2832 7296 3148 7324
rect 2832 7284 2838 7296
rect 3142 7284 3148 7296
rect 3200 7324 3206 7336
rect 5074 7324 5080 7336
rect 3200 7296 5080 7324
rect 3200 7284 3206 7296
rect 5074 7284 5080 7296
rect 5132 7284 5138 7336
rect 5718 7284 5724 7336
rect 5776 7284 5782 7336
rect 7193 7327 7251 7333
rect 7193 7293 7205 7327
rect 7239 7324 7251 7327
rect 7239 7296 8524 7324
rect 7239 7293 7251 7296
rect 7193 7287 7251 7293
rect 5736 7256 5764 7284
rect 6365 7259 6423 7265
rect 6365 7256 6377 7259
rect 5736 7228 6377 7256
rect 6365 7225 6377 7228
rect 6411 7225 6423 7259
rect 8496 7256 8524 7296
rect 9030 7284 9036 7336
rect 9088 7324 9094 7336
rect 9585 7327 9643 7333
rect 9585 7324 9597 7327
rect 9088 7296 9597 7324
rect 9088 7284 9094 7296
rect 9585 7293 9597 7296
rect 9631 7293 9643 7327
rect 9585 7287 9643 7293
rect 9677 7259 9735 7265
rect 9677 7256 9689 7259
rect 8496 7228 9689 7256
rect 6365 7219 6423 7225
rect 9677 7225 9689 7228
rect 9723 7225 9735 7259
rect 9677 7219 9735 7225
rect 2222 7148 2228 7200
rect 2280 7148 2286 7200
rect 4249 7191 4307 7197
rect 4249 7157 4261 7191
rect 4295 7188 4307 7191
rect 4798 7188 4804 7200
rect 4295 7160 4804 7188
rect 4295 7157 4307 7160
rect 4249 7151 4307 7157
rect 4798 7148 4804 7160
rect 4856 7188 4862 7200
rect 5258 7188 5264 7200
rect 4856 7160 5264 7188
rect 4856 7148 4862 7160
rect 5258 7148 5264 7160
rect 5316 7148 5322 7200
rect 5810 7148 5816 7200
rect 5868 7148 5874 7200
rect 8665 7191 8723 7197
rect 8665 7157 8677 7191
rect 8711 7188 8723 7191
rect 8938 7188 8944 7200
rect 8711 7160 8944 7188
rect 8711 7157 8723 7160
rect 8665 7151 8723 7157
rect 8938 7148 8944 7160
rect 8996 7148 9002 7200
rect 9766 7148 9772 7200
rect 9824 7148 9830 7200
rect 1104 7098 10396 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 10396 7098
rect 1104 7024 10396 7046
rect 2028 6987 2086 6993
rect 2028 6953 2040 6987
rect 2074 6984 2086 6987
rect 2774 6984 2780 6996
rect 2074 6956 2780 6984
rect 2074 6953 2086 6956
rect 2028 6947 2086 6953
rect 2774 6944 2780 6956
rect 2832 6944 2838 6996
rect 3513 6987 3571 6993
rect 3513 6953 3525 6987
rect 3559 6984 3571 6987
rect 3602 6984 3608 6996
rect 3559 6956 3608 6984
rect 3559 6953 3571 6956
rect 3513 6947 3571 6953
rect 3602 6944 3608 6956
rect 3660 6944 3666 6996
rect 3878 6944 3884 6996
rect 3936 6984 3942 6996
rect 3936 6956 4108 6984
rect 3936 6944 3942 6956
rect 1486 6876 1492 6928
rect 1544 6876 1550 6928
rect 3620 6916 3648 6944
rect 3970 6916 3976 6928
rect 3620 6888 3976 6916
rect 3970 6876 3976 6888
rect 4028 6876 4034 6928
rect 4080 6916 4108 6956
rect 5350 6944 5356 6996
rect 5408 6984 5414 6996
rect 5813 6987 5871 6993
rect 5813 6984 5825 6987
rect 5408 6956 5825 6984
rect 5408 6944 5414 6956
rect 5813 6953 5825 6956
rect 5859 6953 5871 6987
rect 5813 6947 5871 6953
rect 5994 6944 6000 6996
rect 6052 6984 6058 6996
rect 6273 6987 6331 6993
rect 6273 6984 6285 6987
rect 6052 6956 6285 6984
rect 6052 6944 6058 6956
rect 6273 6953 6285 6956
rect 6319 6953 6331 6987
rect 6273 6947 6331 6953
rect 6362 6944 6368 6996
rect 6420 6984 6426 6996
rect 6546 6984 6552 6996
rect 6420 6956 6552 6984
rect 6420 6944 6426 6956
rect 6546 6944 6552 6956
rect 6604 6984 6610 6996
rect 6641 6987 6699 6993
rect 6641 6984 6653 6987
rect 6604 6956 6653 6984
rect 6604 6944 6610 6956
rect 6641 6953 6653 6956
rect 6687 6953 6699 6987
rect 6641 6947 6699 6953
rect 8478 6944 8484 6996
rect 8536 6984 8542 6996
rect 8595 6987 8653 6993
rect 8595 6984 8607 6987
rect 8536 6956 8607 6984
rect 8536 6944 8542 6956
rect 8595 6953 8607 6956
rect 8641 6953 8653 6987
rect 8595 6947 8653 6953
rect 9585 6987 9643 6993
rect 9585 6953 9597 6987
rect 9631 6984 9643 6987
rect 9766 6984 9772 6996
rect 9631 6956 9772 6984
rect 9631 6953 9643 6956
rect 9585 6947 9643 6953
rect 9766 6944 9772 6956
rect 9824 6944 9830 6996
rect 9858 6944 9864 6996
rect 9916 6944 9922 6996
rect 6089 6919 6147 6925
rect 6089 6916 6101 6919
rect 4080 6888 6101 6916
rect 6089 6885 6101 6888
rect 6135 6885 6147 6919
rect 9490 6916 9496 6928
rect 6089 6879 6147 6885
rect 8680 6888 9496 6916
rect 3418 6808 3424 6860
rect 3476 6848 3482 6860
rect 3789 6851 3847 6857
rect 3789 6848 3801 6851
rect 3476 6820 3801 6848
rect 3476 6808 3482 6820
rect 3789 6817 3801 6820
rect 3835 6817 3847 6851
rect 3789 6811 3847 6817
rect 3878 6808 3884 6860
rect 3936 6808 3942 6860
rect 3988 6848 4016 6876
rect 8680 6860 8708 6888
rect 9490 6876 9496 6888
rect 9548 6876 9554 6928
rect 4249 6851 4307 6857
rect 4249 6848 4261 6851
rect 3988 6820 4261 6848
rect 4249 6817 4261 6820
rect 4295 6817 4307 6851
rect 4709 6851 4767 6857
rect 4709 6848 4721 6851
rect 4249 6811 4307 6817
rect 4356 6820 4721 6848
rect 1673 6783 1731 6789
rect 1673 6749 1685 6783
rect 1719 6749 1731 6783
rect 1673 6743 1731 6749
rect 1688 6712 1716 6743
rect 1762 6740 1768 6792
rect 1820 6740 1826 6792
rect 3510 6740 3516 6792
rect 3568 6740 3574 6792
rect 3896 6780 3924 6808
rect 3973 6783 4031 6789
rect 3973 6780 3985 6783
rect 3896 6752 3985 6780
rect 3973 6749 3985 6752
rect 4019 6749 4031 6783
rect 3973 6743 4031 6749
rect 4065 6783 4123 6789
rect 4065 6749 4077 6783
rect 4111 6749 4123 6783
rect 4065 6743 4123 6749
rect 2038 6712 2044 6724
rect 1688 6684 2044 6712
rect 2038 6672 2044 6684
rect 2096 6672 2102 6724
rect 3050 6672 3056 6724
rect 3108 6672 3114 6724
rect 3326 6672 3332 6724
rect 3384 6712 3390 6724
rect 3528 6712 3556 6740
rect 4080 6712 4108 6743
rect 4154 6740 4160 6792
rect 4212 6740 4218 6792
rect 3384 6684 4108 6712
rect 3384 6672 3390 6684
rect 3418 6604 3424 6656
rect 3476 6644 3482 6656
rect 4356 6644 4384 6820
rect 4709 6817 4721 6820
rect 4755 6817 4767 6851
rect 4709 6811 4767 6817
rect 5074 6808 5080 6860
rect 5132 6848 5138 6860
rect 5169 6851 5227 6857
rect 5169 6848 5181 6851
rect 5132 6820 5181 6848
rect 5132 6808 5138 6820
rect 5169 6817 5181 6820
rect 5215 6817 5227 6851
rect 5169 6811 5227 6817
rect 5258 6808 5264 6860
rect 5316 6848 5322 6860
rect 5316 6820 6500 6848
rect 5316 6808 5322 6820
rect 4430 6740 4436 6792
rect 4488 6780 4494 6792
rect 4801 6783 4859 6789
rect 4801 6780 4813 6783
rect 4488 6752 4813 6780
rect 4488 6740 4494 6752
rect 4801 6749 4813 6752
rect 4847 6749 4859 6783
rect 4801 6743 4859 6749
rect 5350 6740 5356 6792
rect 5408 6780 5414 6792
rect 6362 6780 6368 6792
rect 5408 6752 6368 6780
rect 5408 6740 5414 6752
rect 5767 6749 5840 6752
rect 5445 6715 5503 6721
rect 5445 6681 5457 6715
rect 5491 6712 5503 6715
rect 5534 6712 5540 6724
rect 5491 6684 5540 6712
rect 5491 6681 5503 6684
rect 5445 6675 5503 6681
rect 5534 6672 5540 6684
rect 5592 6672 5598 6724
rect 5767 6715 5779 6749
rect 5813 6718 5840 6749
rect 6362 6740 6368 6752
rect 6420 6740 6426 6792
rect 5994 6721 6000 6724
rect 5813 6715 5825 6718
rect 5767 6709 5825 6715
rect 5971 6715 6000 6721
rect 5971 6681 5983 6715
rect 5971 6675 6000 6681
rect 5994 6672 6000 6675
rect 6052 6672 6058 6724
rect 6472 6721 6500 6820
rect 6546 6808 6552 6860
rect 6604 6848 6610 6860
rect 8662 6848 8668 6860
rect 6604 6820 7144 6848
rect 6604 6808 6610 6820
rect 6914 6740 6920 6792
rect 6972 6740 6978 6792
rect 7116 6789 7144 6820
rect 8404 6820 8668 6848
rect 7101 6783 7159 6789
rect 7101 6749 7113 6783
rect 7147 6749 7159 6783
rect 7101 6743 7159 6749
rect 6457 6715 6515 6721
rect 6457 6681 6469 6715
rect 6503 6681 6515 6715
rect 6457 6675 6515 6681
rect 6638 6672 6644 6724
rect 6696 6712 6702 6724
rect 8404 6721 8432 6820
rect 8662 6808 8668 6820
rect 8720 6808 8726 6860
rect 9876 6848 9904 6944
rect 8772 6820 9904 6848
rect 8772 6780 8800 6820
rect 8938 6780 8944 6792
rect 8496 6752 8800 6780
rect 8864 6752 8944 6780
rect 6733 6715 6791 6721
rect 6733 6712 6745 6715
rect 6696 6684 6745 6712
rect 6696 6672 6702 6684
rect 6733 6681 6745 6684
rect 6779 6681 6791 6715
rect 6733 6675 6791 6681
rect 8389 6715 8447 6721
rect 8389 6681 8401 6715
rect 8435 6681 8447 6715
rect 8389 6675 8447 6681
rect 3476 6616 4384 6644
rect 4433 6647 4491 6653
rect 3476 6604 3482 6616
rect 4433 6613 4445 6647
rect 4479 6644 4491 6647
rect 4706 6644 4712 6656
rect 4479 6616 4712 6644
rect 4479 6613 4491 6616
rect 4433 6607 4491 6613
rect 4706 6604 4712 6616
rect 4764 6604 4770 6656
rect 5626 6604 5632 6656
rect 5684 6604 5690 6656
rect 6257 6647 6315 6653
rect 6257 6613 6269 6647
rect 6303 6644 6315 6647
rect 6362 6644 6368 6656
rect 6303 6616 6368 6644
rect 6303 6613 6315 6616
rect 6257 6607 6315 6613
rect 6362 6604 6368 6616
rect 6420 6604 6426 6656
rect 7006 6604 7012 6656
rect 7064 6604 7070 6656
rect 8496 6644 8524 6752
rect 8605 6715 8663 6721
rect 8605 6681 8617 6715
rect 8651 6712 8663 6715
rect 8864 6712 8892 6752
rect 8938 6740 8944 6752
rect 8996 6780 9002 6792
rect 9125 6783 9183 6789
rect 9125 6780 9137 6783
rect 8996 6752 9137 6780
rect 8996 6740 9002 6752
rect 9125 6749 9137 6752
rect 9171 6749 9183 6783
rect 9125 6743 9183 6749
rect 9306 6740 9312 6792
rect 9364 6740 9370 6792
rect 9582 6740 9588 6792
rect 9640 6740 9646 6792
rect 9861 6783 9919 6789
rect 9861 6749 9873 6783
rect 9907 6749 9919 6783
rect 9861 6743 9919 6749
rect 8651 6684 8892 6712
rect 8651 6681 8663 6684
rect 8605 6675 8663 6681
rect 8757 6647 8815 6653
rect 8757 6644 8769 6647
rect 8496 6616 8769 6644
rect 8757 6613 8769 6616
rect 8803 6613 8815 6647
rect 8757 6607 8815 6613
rect 8938 6604 8944 6656
rect 8996 6604 9002 6656
rect 9214 6604 9220 6656
rect 9272 6604 9278 6656
rect 9324 6644 9352 6740
rect 9490 6672 9496 6724
rect 9548 6712 9554 6724
rect 9769 6715 9827 6721
rect 9769 6712 9781 6715
rect 9548 6684 9781 6712
rect 9548 6672 9554 6684
rect 9769 6681 9781 6684
rect 9815 6681 9827 6715
rect 9769 6675 9827 6681
rect 9876 6644 9904 6743
rect 9324 6616 9904 6644
rect 1104 6554 10396 6576
rect 1104 6502 4874 6554
rect 4926 6502 4938 6554
rect 4990 6502 5002 6554
rect 5054 6502 5066 6554
rect 5118 6502 5130 6554
rect 5182 6502 10396 6554
rect 1104 6480 10396 6502
rect 3697 6443 3755 6449
rect 3697 6409 3709 6443
rect 3743 6440 3755 6443
rect 4338 6440 4344 6452
rect 3743 6412 4344 6440
rect 3743 6409 3755 6412
rect 3697 6403 3755 6409
rect 4338 6400 4344 6412
rect 4396 6400 4402 6452
rect 4430 6400 4436 6452
rect 4488 6400 4494 6452
rect 4614 6400 4620 6452
rect 4672 6440 4678 6452
rect 4709 6443 4767 6449
rect 4709 6440 4721 6443
rect 4672 6412 4721 6440
rect 4672 6400 4678 6412
rect 4709 6409 4721 6412
rect 4755 6409 4767 6443
rect 4709 6403 4767 6409
rect 4890 6400 4896 6452
rect 4948 6400 4954 6452
rect 5718 6400 5724 6452
rect 5776 6440 5782 6452
rect 5813 6443 5871 6449
rect 5813 6440 5825 6443
rect 5776 6412 5825 6440
rect 5776 6400 5782 6412
rect 5813 6409 5825 6412
rect 5859 6409 5871 6443
rect 5813 6403 5871 6409
rect 6365 6443 6423 6449
rect 6365 6409 6377 6443
rect 6411 6440 6423 6443
rect 6638 6440 6644 6452
rect 6411 6412 6644 6440
rect 6411 6409 6423 6412
rect 6365 6403 6423 6409
rect 6638 6400 6644 6412
rect 6696 6400 6702 6452
rect 8938 6400 8944 6452
rect 8996 6400 9002 6452
rect 9309 6443 9367 6449
rect 9309 6409 9321 6443
rect 9355 6440 9367 6443
rect 9674 6440 9680 6452
rect 9355 6412 9680 6440
rect 9355 6409 9367 6412
rect 9309 6403 9367 6409
rect 9674 6400 9680 6412
rect 9732 6400 9738 6452
rect 9950 6400 9956 6452
rect 10008 6400 10014 6452
rect 2130 6332 2136 6384
rect 2188 6332 2194 6384
rect 3605 6375 3663 6381
rect 3605 6341 3617 6375
rect 3651 6372 3663 6375
rect 4798 6372 4804 6384
rect 3651 6344 4804 6372
rect 3651 6341 3663 6344
rect 3605 6335 3663 6341
rect 3421 6307 3479 6313
rect 3421 6273 3433 6307
rect 3467 6304 3479 6307
rect 3510 6304 3516 6316
rect 3467 6276 3516 6304
rect 3467 6273 3479 6276
rect 3421 6267 3479 6273
rect 3510 6264 3516 6276
rect 3568 6264 3574 6316
rect 3896 6313 3924 6344
rect 4798 6332 4804 6344
rect 4856 6372 4862 6384
rect 5353 6375 5411 6381
rect 5353 6372 5365 6375
rect 4856 6344 5365 6372
rect 4856 6332 4862 6344
rect 5353 6341 5365 6344
rect 5399 6341 5411 6375
rect 5353 6335 5411 6341
rect 5534 6338 5540 6384
rect 5460 6332 5540 6338
rect 5592 6332 5598 6384
rect 7098 6372 7104 6384
rect 5920 6344 6776 6372
rect 3697 6307 3755 6313
rect 3697 6302 3709 6307
rect 3620 6274 3709 6302
rect 1397 6239 1455 6245
rect 1397 6205 1409 6239
rect 1443 6205 1455 6239
rect 1397 6199 1455 6205
rect 1673 6239 1731 6245
rect 1673 6205 1685 6239
rect 1719 6236 1731 6239
rect 2222 6236 2228 6248
rect 1719 6208 2228 6236
rect 1719 6205 1731 6208
rect 1673 6199 1731 6205
rect 1412 6100 1440 6199
rect 2222 6196 2228 6208
rect 2280 6196 2286 6248
rect 1762 6100 1768 6112
rect 1412 6072 1768 6100
rect 1762 6060 1768 6072
rect 1820 6100 1826 6112
rect 2222 6100 2228 6112
rect 1820 6072 2228 6100
rect 1820 6060 1826 6072
rect 2222 6060 2228 6072
rect 2280 6060 2286 6112
rect 3142 6060 3148 6112
rect 3200 6060 3206 6112
rect 3620 6100 3648 6274
rect 3697 6273 3709 6274
rect 3743 6273 3755 6307
rect 3697 6267 3755 6273
rect 3881 6307 3939 6313
rect 3881 6273 3893 6307
rect 3927 6273 3939 6307
rect 3881 6267 3939 6273
rect 3970 6264 3976 6316
rect 4028 6264 4034 6316
rect 4154 6264 4160 6316
rect 4212 6304 4218 6316
rect 4525 6307 4583 6313
rect 4525 6304 4537 6307
rect 4212 6276 4537 6304
rect 4212 6264 4218 6276
rect 4525 6273 4537 6276
rect 4571 6273 4583 6307
rect 4525 6267 4583 6273
rect 4617 6307 4675 6313
rect 4617 6273 4629 6307
rect 4663 6273 4675 6307
rect 4617 6267 4675 6273
rect 4893 6307 4951 6313
rect 4893 6273 4905 6307
rect 4939 6304 4951 6307
rect 5074 6304 5080 6316
rect 4939 6276 5080 6304
rect 4939 6273 4951 6276
rect 4893 6267 4951 6273
rect 3988 6236 4016 6264
rect 4632 6236 4660 6267
rect 5074 6264 5080 6276
rect 5132 6264 5138 6316
rect 5460 6313 5580 6332
rect 5920 6316 5948 6344
rect 5261 6310 5319 6313
rect 5184 6307 5319 6310
rect 5184 6282 5273 6307
rect 5184 6236 5212 6282
rect 5261 6273 5273 6282
rect 5307 6273 5319 6307
rect 5261 6267 5319 6273
rect 5445 6310 5580 6313
rect 5813 6310 5871 6313
rect 5902 6310 5908 6316
rect 5445 6307 5503 6310
rect 5445 6273 5457 6307
rect 5491 6273 5503 6307
rect 5445 6267 5503 6273
rect 5813 6307 5908 6310
rect 5813 6273 5825 6307
rect 5859 6282 5908 6307
rect 5859 6273 5871 6282
rect 5813 6267 5871 6273
rect 5902 6264 5908 6282
rect 5960 6264 5966 6316
rect 5994 6264 6000 6316
rect 6052 6264 6058 6316
rect 6089 6307 6147 6313
rect 6089 6273 6101 6307
rect 6135 6304 6147 6307
rect 6178 6304 6184 6316
rect 6135 6276 6184 6304
rect 6135 6273 6147 6276
rect 6089 6267 6147 6273
rect 6178 6264 6184 6276
rect 6236 6304 6242 6316
rect 6546 6304 6552 6316
rect 6236 6276 6552 6304
rect 6236 6264 6242 6276
rect 6546 6264 6552 6276
rect 6604 6264 6610 6316
rect 6748 6313 6776 6344
rect 6840 6344 7104 6372
rect 6840 6313 6868 6344
rect 7098 6332 7104 6344
rect 7156 6372 7162 6384
rect 8956 6372 8984 6400
rect 7156 6344 8984 6372
rect 9692 6372 9720 6400
rect 9692 6344 9812 6372
rect 7156 6332 7162 6344
rect 6641 6307 6699 6313
rect 6641 6273 6653 6307
rect 6687 6273 6699 6307
rect 6641 6267 6699 6273
rect 6733 6307 6791 6313
rect 6733 6273 6745 6307
rect 6779 6273 6791 6307
rect 6733 6267 6791 6273
rect 6825 6307 6883 6313
rect 6825 6273 6837 6307
rect 6871 6273 6883 6307
rect 6825 6267 6883 6273
rect 7009 6307 7067 6313
rect 7009 6273 7021 6307
rect 7055 6273 7067 6307
rect 7009 6267 7067 6273
rect 3988 6208 4660 6236
rect 4816 6208 5212 6236
rect 4816 6100 4844 6208
rect 5184 6180 5212 6208
rect 5721 6239 5779 6245
rect 5721 6205 5733 6239
rect 5767 6236 5779 6239
rect 6012 6236 6040 6264
rect 6656 6236 6684 6267
rect 6914 6236 6920 6248
rect 5767 6208 6040 6236
rect 6104 6208 6920 6236
rect 5767 6205 5779 6208
rect 5721 6199 5779 6205
rect 5166 6128 5172 6180
rect 5224 6128 5230 6180
rect 5902 6128 5908 6180
rect 5960 6168 5966 6180
rect 6104 6168 6132 6208
rect 6914 6196 6920 6208
rect 6972 6196 6978 6248
rect 7024 6236 7052 6267
rect 7190 6264 7196 6316
rect 7248 6304 7254 6316
rect 7929 6307 7987 6313
rect 7929 6304 7941 6307
rect 7248 6276 7941 6304
rect 7248 6264 7254 6276
rect 7929 6273 7941 6276
rect 7975 6273 7987 6307
rect 8956 6304 8984 6344
rect 9784 6313 9812 6344
rect 9125 6307 9183 6313
rect 9125 6304 9137 6307
rect 8956 6276 9137 6304
rect 7929 6267 7987 6273
rect 9125 6273 9137 6276
rect 9171 6273 9183 6307
rect 9125 6267 9183 6273
rect 9677 6307 9735 6313
rect 9677 6273 9689 6307
rect 9723 6273 9735 6307
rect 9677 6267 9735 6273
rect 9769 6307 9827 6313
rect 9769 6273 9781 6307
rect 9815 6273 9827 6307
rect 9769 6267 9827 6273
rect 7653 6239 7711 6245
rect 7653 6236 7665 6239
rect 7024 6208 7665 6236
rect 7653 6205 7665 6208
rect 7699 6236 7711 6239
rect 8662 6236 8668 6248
rect 7699 6208 8668 6236
rect 7699 6205 7711 6208
rect 7653 6199 7711 6205
rect 8662 6196 8668 6208
rect 8720 6236 8726 6248
rect 8941 6239 8999 6245
rect 8941 6236 8953 6239
rect 8720 6208 8953 6236
rect 8720 6196 8726 6208
rect 8941 6205 8953 6208
rect 8987 6205 8999 6239
rect 9692 6236 9720 6267
rect 10318 6264 10324 6316
rect 10376 6264 10382 6316
rect 10336 6236 10364 6264
rect 9692 6208 10364 6236
rect 8941 6199 8999 6205
rect 5960 6140 6132 6168
rect 5960 6128 5966 6140
rect 7006 6128 7012 6180
rect 7064 6128 7070 6180
rect 7745 6171 7803 6177
rect 7745 6137 7757 6171
rect 7791 6168 7803 6171
rect 7791 6140 8340 6168
rect 7791 6137 7803 6140
rect 7745 6131 7803 6137
rect 3620 6072 4844 6100
rect 4982 6060 4988 6112
rect 5040 6060 5046 6112
rect 5074 6060 5080 6112
rect 5132 6100 5138 6112
rect 5629 6103 5687 6109
rect 5629 6100 5641 6103
rect 5132 6072 5641 6100
rect 5132 6060 5138 6072
rect 5629 6069 5641 6072
rect 5675 6100 5687 6103
rect 7024 6100 7052 6128
rect 8312 6112 8340 6140
rect 5675 6072 7052 6100
rect 5675 6069 5687 6072
rect 5629 6063 5687 6069
rect 8110 6060 8116 6112
rect 8168 6060 8174 6112
rect 8294 6060 8300 6112
rect 8352 6060 8358 6112
rect 9398 6060 9404 6112
rect 9456 6100 9462 6112
rect 9493 6103 9551 6109
rect 9493 6100 9505 6103
rect 9456 6072 9505 6100
rect 9456 6060 9462 6072
rect 9493 6069 9505 6072
rect 9539 6100 9551 6103
rect 9582 6100 9588 6112
rect 9539 6072 9588 6100
rect 9539 6069 9551 6072
rect 9493 6063 9551 6069
rect 9582 6060 9588 6072
rect 9640 6060 9646 6112
rect 1104 6010 10396 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 10396 6010
rect 1104 5936 10396 5958
rect 1397 5899 1455 5905
rect 1397 5865 1409 5899
rect 1443 5896 1455 5899
rect 1578 5896 1584 5908
rect 1443 5868 1584 5896
rect 1443 5865 1455 5868
rect 1397 5859 1455 5865
rect 1578 5856 1584 5868
rect 1636 5856 1642 5908
rect 3326 5856 3332 5908
rect 3384 5856 3390 5908
rect 3418 5856 3424 5908
rect 3476 5856 3482 5908
rect 3513 5899 3571 5905
rect 3513 5865 3525 5899
rect 3559 5896 3571 5899
rect 4154 5896 4160 5908
rect 3559 5868 4160 5896
rect 3559 5865 3571 5868
rect 3513 5859 3571 5865
rect 4154 5856 4160 5868
rect 4212 5896 4218 5908
rect 5074 5896 5080 5908
rect 4212 5868 5080 5896
rect 4212 5856 4218 5868
rect 5074 5856 5080 5868
rect 5132 5856 5138 5908
rect 7098 5856 7104 5908
rect 7156 5856 7162 5908
rect 7190 5856 7196 5908
rect 7248 5896 7254 5908
rect 9033 5899 9091 5905
rect 9033 5896 9045 5899
rect 7248 5868 9045 5896
rect 7248 5856 7254 5868
rect 9033 5865 9045 5868
rect 9079 5865 9091 5899
rect 9033 5859 9091 5865
rect 3344 5769 3372 5856
rect 3896 5800 5304 5828
rect 3329 5763 3387 5769
rect 3329 5729 3341 5763
rect 3375 5729 3387 5763
rect 3896 5760 3924 5800
rect 3329 5723 3387 5729
rect 3528 5732 3924 5760
rect 4448 5732 4844 5760
rect 3142 5652 3148 5704
rect 3200 5692 3206 5704
rect 3528 5692 3556 5732
rect 4448 5704 4476 5732
rect 4816 5704 4844 5732
rect 3200 5664 3556 5692
rect 3605 5695 3663 5701
rect 3200 5652 3206 5664
rect 3605 5661 3617 5695
rect 3651 5692 3663 5695
rect 3694 5692 3700 5704
rect 3651 5664 3700 5692
rect 3651 5661 3663 5664
rect 3605 5655 3663 5661
rect 3694 5652 3700 5664
rect 3752 5692 3758 5704
rect 4065 5695 4123 5701
rect 4065 5692 4077 5695
rect 3752 5664 4077 5692
rect 3752 5652 3758 5664
rect 4065 5661 4077 5664
rect 4111 5661 4123 5695
rect 4065 5655 4123 5661
rect 4154 5652 4160 5704
rect 4212 5652 4218 5704
rect 4249 5695 4307 5701
rect 4249 5661 4261 5695
rect 4295 5661 4307 5695
rect 4249 5655 4307 5661
rect 2130 5584 2136 5636
rect 2188 5584 2194 5636
rect 2869 5627 2927 5633
rect 2869 5593 2881 5627
rect 2915 5624 2927 5627
rect 2958 5624 2964 5636
rect 2915 5596 2964 5624
rect 2915 5593 2927 5596
rect 2869 5587 2927 5593
rect 2958 5584 2964 5596
rect 3016 5584 3022 5636
rect 3326 5584 3332 5636
rect 3384 5624 3390 5636
rect 4264 5624 4292 5655
rect 4338 5652 4344 5704
rect 4396 5652 4402 5704
rect 4430 5652 4436 5704
rect 4488 5652 4494 5704
rect 4525 5695 4583 5701
rect 4525 5661 4537 5695
rect 4571 5661 4583 5695
rect 4525 5655 4583 5661
rect 3384 5596 4292 5624
rect 4356 5624 4384 5652
rect 4540 5624 4568 5655
rect 4798 5652 4804 5704
rect 4856 5652 4862 5704
rect 5276 5701 5304 5800
rect 5534 5720 5540 5772
rect 5592 5760 5598 5772
rect 6730 5760 6736 5772
rect 5592 5732 6736 5760
rect 5592 5720 5598 5732
rect 6730 5720 6736 5732
rect 6788 5760 6794 5772
rect 7009 5763 7067 5769
rect 7009 5760 7021 5763
rect 6788 5732 7021 5760
rect 6788 5720 6794 5732
rect 7009 5729 7021 5732
rect 7055 5729 7067 5763
rect 7009 5723 7067 5729
rect 7116 5701 7144 5856
rect 8110 5788 8116 5840
rect 8168 5788 8174 5840
rect 8021 5763 8079 5769
rect 8021 5729 8033 5763
rect 8067 5760 8079 5763
rect 8128 5760 8156 5788
rect 8067 5732 8156 5760
rect 8067 5729 8079 5732
rect 8021 5723 8079 5729
rect 8662 5720 8668 5772
rect 8720 5720 8726 5772
rect 5261 5695 5319 5701
rect 5261 5661 5273 5695
rect 5307 5661 5319 5695
rect 5261 5655 5319 5661
rect 7101 5695 7159 5701
rect 7101 5661 7113 5695
rect 7147 5661 7159 5695
rect 7101 5655 7159 5661
rect 7561 5695 7619 5701
rect 7561 5661 7573 5695
rect 7607 5661 7619 5695
rect 7561 5655 7619 5661
rect 7653 5695 7711 5701
rect 7653 5661 7665 5695
rect 7699 5692 7711 5695
rect 8941 5695 8999 5701
rect 7699 5664 8156 5692
rect 7699 5661 7711 5664
rect 7653 5655 7711 5661
rect 4356 5596 4568 5624
rect 5276 5624 5304 5655
rect 5442 5624 5448 5636
rect 5276 5596 5448 5624
rect 3384 5584 3390 5596
rect 5442 5584 5448 5596
rect 5500 5584 5506 5636
rect 5534 5584 5540 5636
rect 5592 5584 5598 5636
rect 6822 5624 6828 5636
rect 6762 5596 6828 5624
rect 6822 5584 6828 5596
rect 6880 5584 6886 5636
rect 3786 5516 3792 5568
rect 3844 5516 3850 5568
rect 5169 5559 5227 5565
rect 5169 5525 5181 5559
rect 5215 5556 5227 5559
rect 5626 5556 5632 5568
rect 5215 5528 5632 5556
rect 5215 5525 5227 5528
rect 5169 5519 5227 5525
rect 5626 5516 5632 5528
rect 5684 5556 5690 5568
rect 6454 5556 6460 5568
rect 5684 5528 6460 5556
rect 5684 5516 5690 5528
rect 6454 5516 6460 5528
rect 6512 5516 6518 5568
rect 7374 5516 7380 5568
rect 7432 5516 7438 5568
rect 7576 5556 7604 5655
rect 8128 5633 8156 5664
rect 8941 5661 8953 5695
rect 8987 5661 8999 5695
rect 8941 5655 8999 5661
rect 9217 5695 9275 5701
rect 9217 5661 9229 5695
rect 9263 5692 9275 5695
rect 9493 5695 9551 5701
rect 9493 5692 9505 5695
rect 9263 5664 9505 5692
rect 9263 5661 9275 5664
rect 9217 5655 9275 5661
rect 9493 5661 9505 5664
rect 9539 5661 9551 5695
rect 9493 5655 9551 5661
rect 9677 5695 9735 5701
rect 9677 5661 9689 5695
rect 9723 5692 9735 5695
rect 9858 5692 9864 5704
rect 9723 5664 9864 5692
rect 9723 5661 9735 5664
rect 9677 5655 9735 5661
rect 8113 5627 8171 5633
rect 8113 5593 8125 5627
rect 8159 5624 8171 5627
rect 8956 5624 8984 5655
rect 9858 5652 9864 5664
rect 9916 5652 9922 5704
rect 9950 5652 9956 5704
rect 10008 5652 10014 5704
rect 8159 5596 8984 5624
rect 9048 5596 9536 5624
rect 8159 5593 8171 5596
rect 8113 5587 8171 5593
rect 8294 5556 8300 5568
rect 7576 5528 8300 5556
rect 8294 5516 8300 5528
rect 8352 5556 8358 5568
rect 9048 5556 9076 5596
rect 9508 5568 9536 5596
rect 8352 5528 9076 5556
rect 8352 5516 8358 5528
rect 9398 5516 9404 5568
rect 9456 5516 9462 5568
rect 9490 5516 9496 5568
rect 9548 5556 9554 5568
rect 9861 5559 9919 5565
rect 9861 5556 9873 5559
rect 9548 5528 9873 5556
rect 9548 5516 9554 5528
rect 9861 5525 9873 5528
rect 9907 5525 9919 5559
rect 9861 5519 9919 5525
rect 1104 5466 10396 5488
rect 1104 5414 4874 5466
rect 4926 5414 4938 5466
rect 4990 5414 5002 5466
rect 5054 5414 5066 5466
rect 5118 5414 5130 5466
rect 5182 5414 10396 5466
rect 1104 5392 10396 5414
rect 2130 5312 2136 5364
rect 2188 5312 2194 5364
rect 2222 5312 2228 5364
rect 2280 5352 2286 5364
rect 3142 5352 3148 5364
rect 2280 5324 3148 5352
rect 2280 5312 2286 5324
rect 3142 5312 3148 5324
rect 3200 5312 3206 5364
rect 3973 5355 4031 5361
rect 3973 5321 3985 5355
rect 4019 5352 4031 5355
rect 4430 5352 4436 5364
rect 4019 5324 4436 5352
rect 4019 5321 4031 5324
rect 3973 5315 4031 5321
rect 4430 5312 4436 5324
rect 4488 5312 4494 5364
rect 7374 5312 7380 5364
rect 7432 5312 7438 5364
rect 8481 5355 8539 5361
rect 8481 5321 8493 5355
rect 8527 5352 8539 5355
rect 8662 5352 8668 5364
rect 8527 5324 8668 5352
rect 8527 5321 8539 5324
rect 8481 5315 8539 5321
rect 8662 5312 8668 5324
rect 8720 5312 8726 5364
rect 8757 5355 8815 5361
rect 8757 5321 8769 5355
rect 8803 5352 8815 5355
rect 9490 5352 9496 5364
rect 8803 5324 9496 5352
rect 8803 5321 8815 5324
rect 8757 5315 8815 5321
rect 9490 5312 9496 5324
rect 9548 5312 9554 5364
rect 9861 5355 9919 5361
rect 9861 5321 9873 5355
rect 9907 5352 9919 5355
rect 9950 5352 9956 5364
rect 9907 5324 9956 5352
rect 9907 5321 9919 5324
rect 9861 5315 9919 5321
rect 9950 5312 9956 5324
rect 10008 5312 10014 5364
rect 1670 5176 1676 5228
rect 1728 5216 1734 5228
rect 2148 5225 2176 5312
rect 2240 5225 2268 5312
rect 3050 5244 3056 5296
rect 3108 5244 3114 5296
rect 5810 5244 5816 5296
rect 5868 5244 5874 5296
rect 7009 5287 7067 5293
rect 7009 5253 7021 5287
rect 7055 5284 7067 5287
rect 7392 5284 7420 5312
rect 8386 5284 8392 5296
rect 7055 5256 7420 5284
rect 8234 5256 8392 5284
rect 7055 5253 7067 5256
rect 7009 5247 7067 5253
rect 8386 5244 8392 5256
rect 8444 5244 8450 5296
rect 9214 5244 9220 5296
rect 9272 5284 9278 5296
rect 9677 5287 9735 5293
rect 9677 5284 9689 5287
rect 9272 5256 9689 5284
rect 9272 5244 9278 5256
rect 9677 5253 9689 5256
rect 9723 5253 9735 5287
rect 9677 5247 9735 5253
rect 1765 5219 1823 5225
rect 1765 5216 1777 5219
rect 1728 5188 1777 5216
rect 1728 5176 1734 5188
rect 1765 5185 1777 5188
rect 1811 5185 1823 5219
rect 1765 5179 1823 5185
rect 2133 5219 2191 5225
rect 2133 5185 2145 5219
rect 2179 5185 2191 5219
rect 2133 5179 2191 5185
rect 2225 5219 2283 5225
rect 2225 5185 2237 5219
rect 2271 5185 2283 5219
rect 2225 5179 2283 5185
rect 8573 5219 8631 5225
rect 8573 5185 8585 5219
rect 8619 5185 8631 5219
rect 8573 5179 8631 5185
rect 2501 5151 2559 5157
rect 2501 5117 2513 5151
rect 2547 5148 2559 5151
rect 4706 5148 4712 5160
rect 2547 5120 4712 5148
rect 2547 5117 2559 5120
rect 2501 5111 2559 5117
rect 4706 5108 4712 5120
rect 4764 5108 4770 5160
rect 5442 5108 5448 5160
rect 5500 5148 5506 5160
rect 6733 5151 6791 5157
rect 6733 5148 6745 5151
rect 5500 5120 6745 5148
rect 5500 5108 5506 5120
rect 6733 5117 6745 5120
rect 6779 5148 6791 5151
rect 7006 5148 7012 5160
rect 6779 5120 7012 5148
rect 6779 5117 6791 5120
rect 6733 5111 6791 5117
rect 7006 5108 7012 5120
rect 7064 5108 7070 5160
rect 7466 5108 7472 5160
rect 7524 5148 7530 5160
rect 8588 5148 8616 5179
rect 8754 5176 8760 5228
rect 8812 5216 8818 5228
rect 9232 5216 9260 5244
rect 8812 5188 9260 5216
rect 9493 5219 9551 5225
rect 8812 5176 8818 5188
rect 9493 5185 9505 5219
rect 9539 5216 9551 5219
rect 9582 5216 9588 5228
rect 9539 5188 9588 5216
rect 9539 5185 9551 5188
rect 9493 5179 9551 5185
rect 9508 5148 9536 5179
rect 9582 5176 9588 5188
rect 9640 5176 9646 5228
rect 7524 5120 9536 5148
rect 7524 5108 7530 5120
rect 4525 5083 4583 5089
rect 4525 5049 4537 5083
rect 4571 5080 4583 5083
rect 4614 5080 4620 5092
rect 4571 5052 4620 5080
rect 4571 5049 4583 5052
rect 4525 5043 4583 5049
rect 4614 5040 4620 5052
rect 4672 5080 4678 5092
rect 5460 5080 5488 5108
rect 4672 5052 5488 5080
rect 4672 5040 4678 5052
rect 1578 4972 1584 5024
rect 1636 4972 1642 5024
rect 2038 4972 2044 5024
rect 2096 4972 2102 5024
rect 1104 4922 10396 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 10396 4922
rect 1104 4848 10396 4870
rect 1578 4768 1584 4820
rect 1636 4768 1642 4820
rect 2130 4768 2136 4820
rect 2188 4808 2194 4820
rect 2225 4811 2283 4817
rect 2225 4808 2237 4811
rect 2188 4780 2237 4808
rect 2188 4768 2194 4780
rect 2225 4777 2237 4780
rect 2271 4777 2283 4811
rect 2225 4771 2283 4777
rect 5258 4768 5264 4820
rect 5316 4808 5322 4820
rect 5718 4808 5724 4820
rect 5316 4780 5724 4808
rect 5316 4768 5322 4780
rect 5718 4768 5724 4780
rect 5776 4808 5782 4820
rect 5997 4811 6055 4817
rect 5997 4808 6009 4811
rect 5776 4780 6009 4808
rect 5776 4768 5782 4780
rect 5997 4777 6009 4780
rect 6043 4777 6055 4811
rect 5997 4771 6055 4777
rect 6822 4768 6828 4820
rect 6880 4808 6886 4820
rect 8386 4808 8392 4820
rect 6880 4780 8392 4808
rect 6880 4768 6886 4780
rect 8386 4768 8392 4780
rect 8444 4768 8450 4820
rect 8754 4768 8760 4820
rect 8812 4768 8818 4820
rect 9398 4768 9404 4820
rect 9456 4768 9462 4820
rect 1596 4604 1624 4768
rect 4249 4675 4307 4681
rect 4249 4641 4261 4675
rect 4295 4672 4307 4675
rect 4614 4672 4620 4684
rect 4295 4644 4620 4672
rect 4295 4641 4307 4644
rect 4249 4635 4307 4641
rect 4614 4632 4620 4644
rect 4672 4632 4678 4684
rect 6730 4632 6736 4684
rect 6788 4632 6794 4684
rect 1795 4607 1853 4613
rect 1795 4604 1807 4607
rect 1596 4576 1807 4604
rect 1795 4573 1807 4576
rect 1841 4573 1853 4607
rect 1795 4567 1853 4573
rect 1946 4564 1952 4616
rect 2004 4564 2010 4616
rect 2041 4607 2099 4613
rect 2041 4573 2053 4607
rect 2087 4573 2099 4607
rect 6840 4604 6868 4768
rect 7006 4632 7012 4684
rect 7064 4632 7070 4684
rect 7285 4675 7343 4681
rect 7285 4641 7297 4675
rect 7331 4672 7343 4675
rect 9416 4672 9444 4768
rect 7331 4644 9444 4672
rect 7331 4641 7343 4644
rect 7285 4635 7343 4641
rect 5658 4576 6868 4604
rect 2041 4567 2099 4573
rect 1026 4496 1032 4548
rect 1084 4536 1090 4548
rect 2056 4536 2084 4567
rect 8386 4564 8392 4616
rect 8444 4564 8450 4616
rect 1084 4508 2084 4536
rect 1084 4496 1090 4508
rect 4522 4496 4528 4548
rect 4580 4496 4586 4548
rect 1578 4428 1584 4480
rect 1636 4428 1642 4480
rect 6086 4428 6092 4480
rect 6144 4428 6150 4480
rect 1104 4378 10396 4400
rect 1104 4326 4874 4378
rect 4926 4326 4938 4378
rect 4990 4326 5002 4378
rect 5054 4326 5066 4378
rect 5118 4326 5130 4378
rect 5182 4326 10396 4378
rect 1104 4304 10396 4326
rect 1486 4224 1492 4276
rect 1544 4224 1550 4276
rect 1765 4267 1823 4273
rect 1765 4233 1777 4267
rect 1811 4264 1823 4267
rect 1946 4264 1952 4276
rect 1811 4236 1952 4264
rect 1811 4233 1823 4236
rect 1765 4227 1823 4233
rect 1946 4224 1952 4236
rect 2004 4224 2010 4276
rect 6454 4156 6460 4208
rect 6512 4156 6518 4208
rect 1578 4088 1584 4140
rect 1636 4128 1642 4140
rect 1673 4131 1731 4137
rect 1673 4128 1685 4131
rect 1636 4100 1685 4128
rect 1636 4088 1642 4100
rect 1673 4097 1685 4100
rect 1719 4097 1731 4131
rect 1673 4091 1731 4097
rect 1946 4088 1952 4140
rect 2004 4088 2010 4140
rect 4065 4131 4123 4137
rect 4065 4097 4077 4131
rect 4111 4097 4123 4131
rect 4065 4091 4123 4097
rect 4709 4131 4767 4137
rect 4709 4097 4721 4131
rect 4755 4128 4767 4131
rect 6086 4128 6092 4140
rect 4755 4100 6092 4128
rect 4755 4097 4767 4100
rect 4709 4091 4767 4097
rect 3786 4020 3792 4072
rect 3844 4060 3850 4072
rect 3973 4063 4031 4069
rect 3973 4060 3985 4063
rect 3844 4032 3985 4060
rect 3844 4020 3850 4032
rect 3973 4029 3985 4032
rect 4019 4029 4031 4063
rect 3973 4023 4031 4029
rect 4080 3992 4108 4091
rect 6086 4088 6092 4100
rect 6144 4088 6150 4140
rect 4433 4063 4491 4069
rect 4433 4029 4445 4063
rect 4479 4060 4491 4063
rect 4522 4060 4528 4072
rect 4479 4032 4528 4060
rect 4479 4029 4491 4032
rect 4433 4023 4491 4029
rect 4522 4020 4528 4032
rect 4580 4020 4586 4072
rect 4798 4020 4804 4072
rect 4856 4020 4862 4072
rect 5077 4063 5135 4069
rect 5077 4029 5089 4063
rect 5123 4060 5135 4063
rect 5534 4060 5540 4072
rect 5123 4032 5540 4060
rect 5123 4029 5135 4032
rect 5077 4023 5135 4029
rect 5534 4020 5540 4032
rect 5592 4020 5598 4072
rect 5718 4020 5724 4072
rect 5776 4020 5782 4072
rect 6641 4063 6699 4069
rect 6641 4029 6653 4063
rect 6687 4060 6699 4063
rect 6822 4060 6828 4072
rect 6687 4032 6828 4060
rect 6687 4029 6699 4032
rect 6641 4023 6699 4029
rect 6822 4020 6828 4032
rect 6880 4020 6886 4072
rect 5169 3995 5227 4001
rect 5169 3992 5181 3995
rect 4080 3964 5181 3992
rect 5169 3961 5181 3964
rect 5215 3961 5227 3995
rect 5169 3955 5227 3961
rect 1104 3834 10396 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 10396 3834
rect 1104 3760 10396 3782
rect 5534 3612 5540 3664
rect 5592 3652 5598 3664
rect 5813 3655 5871 3661
rect 5813 3652 5825 3655
rect 5592 3624 5825 3652
rect 5592 3612 5598 3624
rect 5813 3621 5825 3624
rect 5859 3621 5871 3655
rect 5813 3615 5871 3621
rect 5905 3655 5963 3661
rect 5905 3621 5917 3655
rect 5951 3652 5963 3655
rect 8478 3652 8484 3664
rect 5951 3624 8484 3652
rect 5951 3621 5963 3624
rect 5905 3615 5963 3621
rect 8478 3612 8484 3624
rect 8536 3612 8542 3664
rect 6086 3584 6092 3596
rect 5000 3556 6092 3584
rect 1670 3476 1676 3528
rect 1728 3476 1734 3528
rect 4062 3476 4068 3528
rect 4120 3516 4126 3528
rect 5000 3525 5028 3556
rect 5920 3525 5948 3556
rect 6086 3544 6092 3556
rect 6144 3544 6150 3596
rect 4985 3519 5043 3525
rect 4985 3516 4997 3519
rect 4120 3488 4997 3516
rect 4120 3476 4126 3488
rect 4985 3485 4997 3488
rect 5031 3485 5043 3519
rect 4985 3479 5043 3485
rect 5077 3519 5135 3525
rect 5077 3485 5089 3519
rect 5123 3485 5135 3519
rect 5077 3479 5135 3485
rect 5169 3519 5227 3525
rect 5169 3485 5181 3519
rect 5215 3516 5227 3519
rect 5629 3519 5687 3525
rect 5629 3516 5641 3519
rect 5215 3488 5641 3516
rect 5215 3485 5227 3488
rect 5169 3479 5227 3485
rect 5629 3485 5641 3488
rect 5675 3485 5687 3519
rect 5629 3479 5687 3485
rect 5905 3519 5963 3525
rect 5905 3485 5917 3519
rect 5951 3485 5963 3519
rect 5905 3479 5963 3485
rect 5997 3519 6055 3525
rect 5997 3485 6009 3519
rect 6043 3485 6055 3519
rect 5997 3479 6055 3485
rect 5092 3448 5120 3479
rect 5092 3420 5580 3448
rect 5552 3392 5580 3420
rect 5644 3392 5672 3479
rect 5718 3408 5724 3460
rect 5776 3448 5782 3460
rect 6012 3448 6040 3479
rect 5776 3420 6040 3448
rect 5776 3408 5782 3420
rect 1210 3340 1216 3392
rect 1268 3380 1274 3392
rect 1489 3383 1547 3389
rect 1489 3380 1501 3383
rect 1268 3352 1501 3380
rect 1268 3340 1274 3352
rect 1489 3349 1501 3352
rect 1535 3349 1547 3383
rect 1489 3343 1547 3349
rect 4798 3340 4804 3392
rect 4856 3340 4862 3392
rect 5534 3340 5540 3392
rect 5592 3340 5598 3392
rect 5626 3340 5632 3392
rect 5684 3340 5690 3392
rect 5994 3340 6000 3392
rect 6052 3380 6058 3392
rect 6181 3383 6239 3389
rect 6181 3380 6193 3383
rect 6052 3352 6193 3380
rect 6052 3340 6058 3352
rect 6181 3349 6193 3352
rect 6227 3349 6239 3383
rect 6181 3343 6239 3349
rect 1104 3290 10396 3312
rect 1104 3238 4874 3290
rect 4926 3238 4938 3290
rect 4990 3238 5002 3290
rect 5054 3238 5066 3290
rect 5118 3238 5130 3290
rect 5182 3238 10396 3290
rect 1104 3216 10396 3238
rect 1670 3136 1676 3188
rect 1728 3176 1734 3188
rect 1857 3179 1915 3185
rect 1857 3176 1869 3179
rect 1728 3148 1869 3176
rect 1728 3136 1734 3148
rect 1857 3145 1869 3148
rect 1903 3145 1915 3179
rect 3878 3176 3884 3188
rect 1857 3139 1915 3145
rect 3252 3148 3884 3176
rect 1394 3000 1400 3052
rect 1452 3000 1458 3052
rect 1765 3043 1823 3049
rect 1765 3040 1777 3043
rect 1596 3012 1777 3040
rect 1596 2913 1624 3012
rect 1765 3009 1777 3012
rect 1811 3009 1823 3043
rect 1765 3003 1823 3009
rect 2958 3000 2964 3052
rect 3016 3000 3022 3052
rect 3252 2984 3280 3148
rect 3878 3136 3884 3148
rect 3936 3176 3942 3188
rect 4203 3179 4261 3185
rect 4203 3176 4215 3179
rect 3936 3148 4215 3176
rect 3936 3136 3942 3148
rect 4203 3145 4215 3148
rect 4249 3145 4261 3179
rect 4203 3139 4261 3145
rect 5537 3179 5595 3185
rect 5537 3145 5549 3179
rect 5583 3176 5595 3179
rect 5718 3176 5724 3188
rect 5583 3148 5724 3176
rect 5583 3145 5595 3148
rect 5537 3139 5595 3145
rect 5718 3136 5724 3148
rect 5776 3136 5782 3188
rect 6181 3179 6239 3185
rect 5828 3148 6132 3176
rect 5353 3111 5411 3117
rect 5353 3108 5365 3111
rect 3344 3080 5365 3108
rect 3234 2932 3240 2984
rect 3292 2932 3298 2984
rect 3344 2981 3372 3080
rect 5353 3077 5365 3080
rect 5399 3077 5411 3111
rect 5828 3108 5856 3148
rect 5353 3071 5411 3077
rect 5644 3080 5856 3108
rect 4062 3040 4068 3052
rect 3528 3012 4068 3040
rect 3528 2984 3556 3012
rect 4062 3000 4068 3012
rect 4120 3040 4126 3052
rect 4985 3043 5043 3049
rect 4985 3040 4997 3043
rect 4120 3012 4997 3040
rect 4120 3000 4126 3012
rect 4985 3009 4997 3012
rect 5031 3009 5043 3043
rect 5368 3040 5396 3071
rect 5644 3052 5672 3080
rect 5994 3068 6000 3120
rect 6052 3068 6058 3120
rect 6104 3108 6132 3148
rect 6181 3145 6193 3179
rect 6227 3176 6239 3179
rect 7834 3176 7840 3188
rect 6227 3148 7840 3176
rect 6227 3145 6239 3148
rect 6181 3139 6239 3145
rect 7834 3136 7840 3148
rect 7892 3136 7898 3188
rect 6549 3111 6607 3117
rect 6549 3108 6561 3111
rect 6104 3080 6561 3108
rect 6549 3077 6561 3080
rect 6595 3077 6607 3111
rect 6549 3071 6607 3077
rect 5626 3040 5632 3052
rect 5368 3012 5632 3040
rect 4985 3003 5043 3009
rect 5626 3000 5632 3012
rect 5684 3000 5690 3052
rect 3329 2975 3387 2981
rect 3329 2941 3341 2975
rect 3375 2941 3387 2975
rect 3329 2935 3387 2941
rect 3421 2975 3479 2981
rect 3421 2941 3433 2975
rect 3467 2972 3479 2975
rect 3510 2972 3516 2984
rect 3467 2944 3516 2972
rect 3467 2941 3479 2944
rect 3421 2935 3479 2941
rect 1581 2907 1639 2913
rect 1581 2873 1593 2907
rect 1627 2873 1639 2907
rect 3344 2904 3372 2935
rect 3510 2932 3516 2944
rect 3568 2932 3574 2984
rect 3970 2932 3976 2984
rect 4028 2932 4034 2984
rect 6012 2904 6040 3068
rect 6086 2932 6092 2984
rect 6144 2972 6150 2984
rect 6917 2975 6975 2981
rect 6917 2972 6929 2975
rect 6144 2944 6929 2972
rect 6144 2932 6150 2944
rect 6917 2941 6929 2944
rect 6963 2941 6975 2975
rect 6917 2935 6975 2941
rect 3344 2876 3464 2904
rect 6012 2876 6592 2904
rect 1581 2867 1639 2873
rect 3436 2848 3464 2876
rect 2590 2796 2596 2848
rect 2648 2836 2654 2848
rect 2777 2839 2835 2845
rect 2777 2836 2789 2839
rect 2648 2808 2789 2836
rect 2648 2796 2654 2808
rect 2777 2805 2789 2808
rect 2823 2805 2835 2839
rect 2777 2799 2835 2805
rect 3418 2796 3424 2848
rect 3476 2796 3482 2848
rect 3602 2796 3608 2848
rect 3660 2796 3666 2848
rect 3878 2796 3884 2848
rect 3936 2836 3942 2848
rect 5353 2839 5411 2845
rect 5353 2836 5365 2839
rect 3936 2808 5365 2836
rect 3936 2796 3942 2808
rect 5353 2805 5365 2808
rect 5399 2836 5411 2839
rect 5534 2836 5540 2848
rect 5399 2808 5540 2836
rect 5399 2805 5411 2808
rect 5353 2799 5411 2805
rect 5534 2796 5540 2808
rect 5592 2836 5598 2848
rect 5994 2836 6000 2848
rect 5592 2808 6000 2836
rect 5592 2796 5598 2808
rect 5994 2796 6000 2808
rect 6052 2796 6058 2848
rect 6362 2796 6368 2848
rect 6420 2796 6426 2848
rect 6564 2845 6592 2876
rect 6549 2839 6607 2845
rect 6549 2805 6561 2839
rect 6595 2805 6607 2839
rect 6549 2799 6607 2805
rect 1104 2746 10396 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 10396 2746
rect 1104 2672 10396 2694
rect 2958 2592 2964 2644
rect 3016 2632 3022 2644
rect 3145 2635 3203 2641
rect 3145 2632 3157 2635
rect 3016 2604 3157 2632
rect 3016 2592 3022 2604
rect 3145 2601 3157 2604
rect 3191 2601 3203 2635
rect 3145 2595 3203 2601
rect 5994 2592 6000 2644
rect 6052 2592 6058 2644
rect 3436 2536 4936 2564
rect 3436 2508 3464 2536
rect 3234 2456 3240 2508
rect 3292 2496 3298 2508
rect 3329 2499 3387 2505
rect 3329 2496 3341 2499
rect 3292 2468 3341 2496
rect 3292 2456 3298 2468
rect 3329 2465 3341 2468
rect 3375 2465 3387 2499
rect 3329 2459 3387 2465
rect 3418 2456 3424 2508
rect 3476 2456 3482 2508
rect 4908 2505 4936 2536
rect 4893 2499 4951 2505
rect 4540 2468 4844 2496
rect 2038 2388 2044 2440
rect 2096 2388 2102 2440
rect 2317 2431 2375 2437
rect 2317 2397 2329 2431
rect 2363 2428 2375 2431
rect 3510 2428 3516 2440
rect 2363 2400 3516 2428
rect 2363 2397 2375 2400
rect 2317 2391 2375 2397
rect 3510 2388 3516 2400
rect 3568 2388 3574 2440
rect 3602 2388 3608 2440
rect 3660 2428 3666 2440
rect 4540 2437 4568 2468
rect 4816 2440 4844 2468
rect 4893 2465 4905 2499
rect 4939 2465 4951 2499
rect 4893 2459 4951 2465
rect 3789 2431 3847 2437
rect 3789 2428 3801 2431
rect 3660 2400 3801 2428
rect 3660 2388 3666 2400
rect 3789 2397 3801 2400
rect 3835 2397 3847 2431
rect 3789 2391 3847 2397
rect 4525 2431 4583 2437
rect 4525 2397 4537 2431
rect 4571 2397 4583 2431
rect 4525 2391 4583 2397
rect 4614 2388 4620 2440
rect 4672 2388 4678 2440
rect 4798 2388 4804 2440
rect 4856 2388 4862 2440
rect 4908 2360 4936 2459
rect 5902 2388 5908 2440
rect 5960 2388 5966 2440
rect 6362 2388 6368 2440
rect 6420 2428 6426 2440
rect 6549 2431 6607 2437
rect 6549 2428 6561 2431
rect 6420 2400 6561 2428
rect 6420 2388 6426 2400
rect 6549 2397 6561 2400
rect 6595 2397 6607 2431
rect 7193 2431 7251 2437
rect 7193 2428 7205 2431
rect 6549 2391 6607 2397
rect 6886 2400 7205 2428
rect 5813 2363 5871 2369
rect 5813 2360 5825 2363
rect 4908 2332 5825 2360
rect 5813 2329 5825 2332
rect 5859 2329 5871 2363
rect 5920 2360 5948 2388
rect 6013 2363 6071 2369
rect 6013 2360 6025 2363
rect 5920 2332 6025 2360
rect 5813 2323 5871 2329
rect 6013 2329 6025 2332
rect 6059 2329 6071 2363
rect 6886 2360 6914 2400
rect 7193 2397 7205 2400
rect 7239 2397 7251 2431
rect 7193 2391 7251 2397
rect 7834 2388 7840 2440
rect 7892 2388 7898 2440
rect 8478 2388 8484 2440
rect 8536 2388 8542 2440
rect 6013 2323 6071 2329
rect 6196 2332 6914 2360
rect 3234 2252 3240 2304
rect 3292 2292 3298 2304
rect 3973 2295 4031 2301
rect 3973 2292 3985 2295
rect 3292 2264 3985 2292
rect 3292 2252 3298 2264
rect 3973 2261 3985 2264
rect 4019 2261 4031 2295
rect 3973 2255 4031 2261
rect 4341 2295 4399 2301
rect 4341 2261 4353 2295
rect 4387 2292 4399 2295
rect 4798 2292 4804 2304
rect 4387 2264 4804 2292
rect 4387 2261 4399 2264
rect 4341 2255 4399 2261
rect 4798 2252 4804 2264
rect 4856 2252 4862 2304
rect 6196 2301 6224 2332
rect 6181 2295 6239 2301
rect 6181 2261 6193 2295
rect 6227 2261 6239 2295
rect 6181 2255 6239 2261
rect 6454 2252 6460 2304
rect 6512 2292 6518 2304
rect 6733 2295 6791 2301
rect 6733 2292 6745 2295
rect 6512 2264 6745 2292
rect 6512 2252 6518 2264
rect 6733 2261 6745 2264
rect 6779 2261 6791 2295
rect 6733 2255 6791 2261
rect 7098 2252 7104 2304
rect 7156 2292 7162 2304
rect 7377 2295 7435 2301
rect 7377 2292 7389 2295
rect 7156 2264 7389 2292
rect 7156 2252 7162 2264
rect 7377 2261 7389 2264
rect 7423 2261 7435 2295
rect 7377 2255 7435 2261
rect 7742 2252 7748 2304
rect 7800 2292 7806 2304
rect 8021 2295 8079 2301
rect 8021 2292 8033 2295
rect 7800 2264 8033 2292
rect 7800 2252 7806 2264
rect 8021 2261 8033 2264
rect 8067 2261 8079 2295
rect 8021 2255 8079 2261
rect 8386 2252 8392 2304
rect 8444 2292 8450 2304
rect 8665 2295 8723 2301
rect 8665 2292 8677 2295
rect 8444 2264 8677 2292
rect 8444 2252 8450 2264
rect 8665 2261 8677 2264
rect 8711 2261 8723 2295
rect 8665 2255 8723 2261
rect 1104 2202 10396 2224
rect 1104 2150 4874 2202
rect 4926 2150 4938 2202
rect 4990 2150 5002 2202
rect 5054 2150 5066 2202
rect 5118 2150 5130 2202
rect 5182 2150 10396 2202
rect 1104 2128 10396 2150
<< via1 >>
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 5816 11296 5868 11348
rect 6092 11271 6144 11280
rect 6092 11237 6101 11271
rect 6101 11237 6135 11271
rect 6135 11237 6144 11271
rect 6092 11228 6144 11237
rect 4804 11160 4856 11212
rect 5816 11135 5868 11144
rect 5816 11101 5825 11135
rect 5825 11101 5859 11135
rect 5859 11101 5868 11135
rect 5816 11092 5868 11101
rect 6736 11092 6788 11144
rect 5264 11024 5316 11076
rect 5632 11024 5684 11076
rect 4712 10956 4764 11008
rect 5908 10999 5960 11008
rect 5908 10965 5917 10999
rect 5917 10965 5951 10999
rect 5951 10965 5960 10999
rect 5908 10956 5960 10965
rect 4874 10854 4926 10906
rect 4938 10854 4990 10906
rect 5002 10854 5054 10906
rect 5066 10854 5118 10906
rect 5130 10854 5182 10906
rect 5816 10795 5868 10804
rect 4160 10616 4212 10668
rect 5816 10761 5841 10795
rect 5841 10761 5868 10795
rect 5816 10752 5868 10761
rect 6000 10752 6052 10804
rect 6092 10752 6144 10804
rect 5632 10727 5684 10736
rect 5632 10693 5641 10727
rect 5641 10693 5675 10727
rect 5675 10693 5684 10727
rect 5632 10684 5684 10693
rect 5080 10659 5132 10668
rect 5080 10625 5090 10659
rect 5090 10625 5124 10659
rect 5124 10625 5132 10659
rect 5080 10616 5132 10625
rect 2780 10591 2832 10600
rect 2780 10557 2789 10591
rect 2789 10557 2823 10591
rect 2823 10557 2832 10591
rect 2780 10548 2832 10557
rect 3056 10591 3108 10600
rect 3056 10557 3065 10591
rect 3065 10557 3099 10591
rect 3099 10557 3108 10591
rect 3056 10548 3108 10557
rect 3516 10412 3568 10464
rect 5632 10548 5684 10600
rect 6644 10591 6696 10600
rect 6644 10557 6653 10591
rect 6653 10557 6687 10591
rect 6687 10557 6696 10591
rect 6644 10548 6696 10557
rect 4528 10455 4580 10464
rect 4528 10421 4537 10455
rect 4537 10421 4571 10455
rect 4571 10421 4580 10455
rect 4528 10412 4580 10421
rect 5080 10412 5132 10464
rect 5908 10412 5960 10464
rect 6552 10455 6604 10464
rect 6552 10421 6561 10455
rect 6561 10421 6595 10455
rect 6595 10421 6604 10455
rect 6552 10412 6604 10421
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 3056 10208 3108 10260
rect 4344 10208 4396 10260
rect 4804 10208 4856 10260
rect 6184 10208 6236 10260
rect 2780 10140 2832 10192
rect 5540 10140 5592 10192
rect 3516 10072 3568 10124
rect 4712 10072 4764 10124
rect 2872 9936 2924 9988
rect 4252 10004 4304 10056
rect 4344 10004 4396 10056
rect 4620 10047 4672 10056
rect 4620 10013 4629 10047
rect 4629 10013 4663 10047
rect 4663 10013 4672 10047
rect 4620 10004 4672 10013
rect 5356 10072 5408 10124
rect 5908 10072 5960 10124
rect 2964 9911 3016 9920
rect 2964 9877 2973 9911
rect 2973 9877 3007 9911
rect 3007 9877 3016 9911
rect 2964 9868 3016 9877
rect 3148 9911 3200 9920
rect 3148 9877 3157 9911
rect 3157 9877 3191 9911
rect 3191 9877 3200 9911
rect 3148 9868 3200 9877
rect 4344 9911 4396 9920
rect 4344 9877 4353 9911
rect 4353 9877 4387 9911
rect 4387 9877 4396 9911
rect 4344 9868 4396 9877
rect 4436 9911 4488 9920
rect 4436 9877 4445 9911
rect 4445 9877 4479 9911
rect 4479 9877 4488 9911
rect 4436 9868 4488 9877
rect 4528 9868 4580 9920
rect 5540 10047 5592 10056
rect 5540 10013 5549 10047
rect 5549 10013 5583 10047
rect 5583 10013 5592 10047
rect 5540 10004 5592 10013
rect 6920 10004 6972 10056
rect 5816 9979 5868 9988
rect 5816 9945 5825 9979
rect 5825 9945 5859 9979
rect 5859 9945 5868 9979
rect 5816 9936 5868 9945
rect 5908 9936 5960 9988
rect 5632 9868 5684 9920
rect 4874 9766 4926 9818
rect 4938 9766 4990 9818
rect 5002 9766 5054 9818
rect 5066 9766 5118 9818
rect 5130 9766 5182 9818
rect 4528 9707 4580 9716
rect 4528 9673 4537 9707
rect 4537 9673 4571 9707
rect 4571 9673 4580 9707
rect 4528 9664 4580 9673
rect 5356 9664 5408 9716
rect 5816 9664 5868 9716
rect 7012 9664 7064 9716
rect 3148 9596 3200 9648
rect 4620 9596 4672 9648
rect 5264 9639 5316 9648
rect 5264 9605 5273 9639
rect 5273 9605 5307 9639
rect 5307 9605 5316 9639
rect 5264 9596 5316 9605
rect 2780 9571 2832 9580
rect 2780 9537 2789 9571
rect 2789 9537 2823 9571
rect 2823 9537 2832 9571
rect 2780 9528 2832 9537
rect 4160 9528 4212 9580
rect 4344 9528 4396 9580
rect 5540 9596 5592 9648
rect 6552 9596 6604 9648
rect 6000 9528 6052 9580
rect 6368 9571 6420 9580
rect 6368 9537 6377 9571
rect 6377 9537 6411 9571
rect 6411 9537 6420 9571
rect 6368 9528 6420 9537
rect 5632 9460 5684 9512
rect 5724 9503 5776 9512
rect 5724 9469 5733 9503
rect 5733 9469 5767 9503
rect 5767 9469 5776 9503
rect 5724 9460 5776 9469
rect 5908 9460 5960 9512
rect 4252 9392 4304 9444
rect 5448 9324 5500 9376
rect 7012 9324 7064 9376
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 2964 9120 3016 9172
rect 5724 9120 5776 9172
rect 4160 8984 4212 9036
rect 5356 8984 5408 9036
rect 6000 8916 6052 8968
rect 9404 8916 9456 8968
rect 4620 8780 4672 8832
rect 5816 8848 5868 8900
rect 5632 8780 5684 8832
rect 6368 8780 6420 8832
rect 6828 8823 6880 8832
rect 6828 8789 6837 8823
rect 6837 8789 6871 8823
rect 6871 8789 6880 8823
rect 6828 8780 6880 8789
rect 8944 8823 8996 8832
rect 8944 8789 8953 8823
rect 8953 8789 8987 8823
rect 8987 8789 8996 8823
rect 8944 8780 8996 8789
rect 4874 8678 4926 8730
rect 4938 8678 4990 8730
rect 5002 8678 5054 8730
rect 5066 8678 5118 8730
rect 5130 8678 5182 8730
rect 3976 8619 4028 8628
rect 1400 8483 1452 8492
rect 1400 8449 1409 8483
rect 1409 8449 1443 8483
rect 1443 8449 1452 8483
rect 1400 8440 1452 8449
rect 2872 8440 2924 8492
rect 3976 8585 3985 8619
rect 3985 8585 4019 8619
rect 4019 8585 4028 8619
rect 3976 8576 4028 8585
rect 3424 8508 3476 8560
rect 5540 8619 5592 8628
rect 5540 8585 5549 8619
rect 5549 8585 5583 8619
rect 5583 8585 5592 8619
rect 5540 8576 5592 8585
rect 6644 8576 6696 8628
rect 8944 8576 8996 8628
rect 3240 8483 3292 8492
rect 3240 8449 3249 8483
rect 3249 8449 3283 8483
rect 3283 8449 3292 8483
rect 3240 8440 3292 8449
rect 1676 8304 1728 8356
rect 2964 8304 3016 8356
rect 2872 8236 2924 8288
rect 3516 8483 3568 8492
rect 3516 8449 3525 8483
rect 3525 8449 3559 8483
rect 3559 8449 3568 8483
rect 3516 8440 3568 8449
rect 3608 8415 3660 8424
rect 3608 8381 3617 8415
rect 3617 8381 3651 8415
rect 3651 8381 3660 8415
rect 3608 8372 3660 8381
rect 3884 8440 3936 8492
rect 4896 8440 4948 8492
rect 5632 8440 5684 8492
rect 4068 8304 4120 8356
rect 3884 8236 3936 8288
rect 6000 8440 6052 8492
rect 6092 8483 6144 8492
rect 6092 8449 6101 8483
rect 6101 8449 6135 8483
rect 6135 8449 6144 8483
rect 6092 8440 6144 8449
rect 8392 8508 8444 8560
rect 6828 8440 6880 8492
rect 9036 8508 9088 8560
rect 9404 8508 9456 8560
rect 9220 8483 9272 8492
rect 9220 8449 9221 8483
rect 9221 8449 9255 8483
rect 9255 8449 9272 8483
rect 9220 8440 9272 8449
rect 9496 8483 9548 8492
rect 9496 8449 9505 8483
rect 9505 8449 9539 8483
rect 9539 8449 9548 8483
rect 9496 8440 9548 8449
rect 9680 8483 9732 8492
rect 9680 8449 9689 8483
rect 9689 8449 9723 8483
rect 9723 8449 9732 8483
rect 9680 8440 9732 8449
rect 8484 8304 8536 8356
rect 4804 8279 4856 8288
rect 4804 8245 4813 8279
rect 4813 8245 4847 8279
rect 4847 8245 4856 8279
rect 4804 8236 4856 8245
rect 5264 8279 5316 8288
rect 5264 8245 5273 8279
rect 5273 8245 5307 8279
rect 5307 8245 5316 8279
rect 5264 8236 5316 8245
rect 5724 8279 5776 8288
rect 5724 8245 5733 8279
rect 5733 8245 5767 8279
rect 5767 8245 5776 8279
rect 5724 8236 5776 8245
rect 9312 8279 9364 8288
rect 9312 8245 9321 8279
rect 9321 8245 9355 8279
rect 9355 8245 9364 8279
rect 9312 8236 9364 8245
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 3240 8032 3292 8084
rect 2780 7896 2832 7948
rect 3884 7896 3936 7948
rect 4804 8032 4856 8084
rect 5540 8032 5592 8084
rect 4620 7964 4672 8016
rect 3516 7828 3568 7880
rect 3608 7871 3660 7880
rect 3608 7837 3617 7871
rect 3617 7837 3651 7871
rect 3651 7837 3660 7871
rect 3608 7828 3660 7837
rect 3792 7871 3844 7880
rect 3792 7837 3801 7871
rect 3801 7837 3835 7871
rect 3835 7837 3844 7871
rect 3792 7828 3844 7837
rect 3976 7871 4028 7880
rect 3976 7837 3985 7871
rect 3985 7837 4019 7871
rect 4019 7837 4028 7871
rect 3976 7828 4028 7837
rect 4160 7871 4212 7880
rect 4160 7837 4169 7871
rect 4169 7837 4203 7871
rect 4203 7837 4212 7871
rect 4160 7828 4212 7837
rect 4804 7939 4856 7948
rect 4804 7905 4813 7939
rect 4813 7905 4847 7939
rect 4847 7905 4856 7939
rect 4804 7896 4856 7905
rect 5172 7896 5224 7948
rect 5356 7896 5408 7948
rect 6828 7939 6880 7948
rect 6828 7905 6837 7939
rect 6837 7905 6871 7939
rect 6871 7905 6880 7939
rect 6828 7896 6880 7905
rect 8392 7896 8444 7948
rect 9128 7896 9180 7948
rect 5264 7828 5316 7880
rect 5448 7828 5500 7880
rect 8944 7871 8996 7880
rect 8944 7837 8953 7871
rect 8953 7837 8987 7871
rect 8987 7837 8996 7871
rect 8944 7828 8996 7837
rect 9404 7828 9456 7880
rect 2780 7760 2832 7812
rect 4068 7692 4120 7744
rect 4896 7692 4948 7744
rect 5264 7692 5316 7744
rect 7196 7803 7248 7812
rect 7196 7769 7205 7803
rect 7205 7769 7239 7803
rect 7239 7769 7248 7803
rect 7196 7760 7248 7769
rect 9220 7760 9272 7812
rect 8668 7735 8720 7744
rect 8668 7701 8677 7735
rect 8677 7701 8711 7735
rect 8711 7701 8720 7735
rect 8668 7692 8720 7701
rect 9588 7735 9640 7744
rect 9588 7701 9597 7735
rect 9597 7701 9631 7735
rect 9631 7701 9640 7735
rect 9588 7692 9640 7701
rect 4874 7590 4926 7642
rect 4938 7590 4990 7642
rect 5002 7590 5054 7642
rect 5066 7590 5118 7642
rect 5130 7590 5182 7642
rect 3792 7488 3844 7540
rect 6000 7488 6052 7540
rect 6552 7488 6604 7540
rect 3056 7420 3108 7472
rect 4712 7420 4764 7472
rect 5356 7420 5408 7472
rect 4620 7352 4672 7404
rect 6000 7352 6052 7404
rect 6460 7352 6512 7404
rect 7012 7488 7064 7540
rect 7196 7488 7248 7540
rect 6828 7352 6880 7404
rect 9128 7488 9180 7540
rect 9312 7352 9364 7404
rect 9680 7488 9732 7540
rect 9496 7395 9548 7404
rect 9496 7361 9505 7395
rect 9505 7361 9539 7395
rect 9539 7361 9548 7395
rect 9496 7352 9548 7361
rect 9864 7395 9916 7404
rect 9864 7361 9873 7395
rect 9873 7361 9907 7395
rect 9907 7361 9916 7395
rect 9864 7352 9916 7361
rect 1584 7327 1636 7336
rect 1584 7293 1593 7327
rect 1593 7293 1627 7327
rect 1627 7293 1636 7327
rect 1584 7284 1636 7293
rect 1768 7284 1820 7336
rect 2780 7284 2832 7336
rect 3148 7284 3200 7336
rect 5080 7284 5132 7336
rect 5724 7284 5776 7336
rect 9036 7284 9088 7336
rect 2228 7191 2280 7200
rect 2228 7157 2237 7191
rect 2237 7157 2271 7191
rect 2271 7157 2280 7191
rect 2228 7148 2280 7157
rect 4804 7148 4856 7200
rect 5264 7148 5316 7200
rect 5816 7191 5868 7200
rect 5816 7157 5825 7191
rect 5825 7157 5859 7191
rect 5859 7157 5868 7191
rect 5816 7148 5868 7157
rect 8944 7148 8996 7200
rect 9772 7191 9824 7200
rect 9772 7157 9781 7191
rect 9781 7157 9815 7191
rect 9815 7157 9824 7191
rect 9772 7148 9824 7157
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 2780 6944 2832 6996
rect 3608 6944 3660 6996
rect 3884 6944 3936 6996
rect 1492 6919 1544 6928
rect 1492 6885 1501 6919
rect 1501 6885 1535 6919
rect 1535 6885 1544 6919
rect 1492 6876 1544 6885
rect 3976 6876 4028 6928
rect 5356 6944 5408 6996
rect 6000 6944 6052 6996
rect 6368 6944 6420 6996
rect 6552 6944 6604 6996
rect 8484 6944 8536 6996
rect 9772 6944 9824 6996
rect 9864 6944 9916 6996
rect 9496 6919 9548 6928
rect 3424 6808 3476 6860
rect 3884 6808 3936 6860
rect 9496 6885 9505 6919
rect 9505 6885 9539 6919
rect 9539 6885 9548 6919
rect 9496 6876 9548 6885
rect 1768 6783 1820 6792
rect 1768 6749 1777 6783
rect 1777 6749 1811 6783
rect 1811 6749 1820 6783
rect 1768 6740 1820 6749
rect 3516 6740 3568 6792
rect 2044 6672 2096 6724
rect 3056 6672 3108 6724
rect 3332 6672 3384 6724
rect 4160 6783 4212 6792
rect 4160 6749 4169 6783
rect 4169 6749 4203 6783
rect 4203 6749 4212 6783
rect 4160 6740 4212 6749
rect 3424 6604 3476 6656
rect 5080 6808 5132 6860
rect 5264 6808 5316 6860
rect 4436 6740 4488 6792
rect 5356 6740 5408 6792
rect 5540 6672 5592 6724
rect 6368 6740 6420 6792
rect 6000 6715 6052 6724
rect 6000 6681 6017 6715
rect 6017 6681 6052 6715
rect 6000 6672 6052 6681
rect 6552 6808 6604 6860
rect 6920 6783 6972 6792
rect 6920 6749 6929 6783
rect 6929 6749 6963 6783
rect 6963 6749 6972 6783
rect 6920 6740 6972 6749
rect 6644 6672 6696 6724
rect 8668 6808 8720 6860
rect 4712 6604 4764 6656
rect 5632 6647 5684 6656
rect 5632 6613 5641 6647
rect 5641 6613 5675 6647
rect 5675 6613 5684 6647
rect 5632 6604 5684 6613
rect 6368 6604 6420 6656
rect 7012 6647 7064 6656
rect 7012 6613 7021 6647
rect 7021 6613 7055 6647
rect 7055 6613 7064 6647
rect 7012 6604 7064 6613
rect 8944 6740 8996 6792
rect 9312 6783 9364 6792
rect 9312 6749 9321 6783
rect 9321 6749 9355 6783
rect 9355 6749 9364 6783
rect 9312 6740 9364 6749
rect 9588 6783 9640 6792
rect 9588 6749 9597 6783
rect 9597 6749 9631 6783
rect 9631 6749 9640 6783
rect 9588 6740 9640 6749
rect 8944 6647 8996 6656
rect 8944 6613 8953 6647
rect 8953 6613 8987 6647
rect 8987 6613 8996 6647
rect 8944 6604 8996 6613
rect 9220 6647 9272 6656
rect 9220 6613 9229 6647
rect 9229 6613 9263 6647
rect 9263 6613 9272 6647
rect 9220 6604 9272 6613
rect 9496 6672 9548 6724
rect 4874 6502 4926 6554
rect 4938 6502 4990 6554
rect 5002 6502 5054 6554
rect 5066 6502 5118 6554
rect 5130 6502 5182 6554
rect 4344 6400 4396 6452
rect 4436 6443 4488 6452
rect 4436 6409 4445 6443
rect 4445 6409 4479 6443
rect 4479 6409 4488 6443
rect 4436 6400 4488 6409
rect 4620 6400 4672 6452
rect 4896 6443 4948 6452
rect 4896 6409 4905 6443
rect 4905 6409 4939 6443
rect 4939 6409 4948 6443
rect 4896 6400 4948 6409
rect 5724 6400 5776 6452
rect 6644 6400 6696 6452
rect 8944 6400 8996 6452
rect 9680 6400 9732 6452
rect 9956 6443 10008 6452
rect 9956 6409 9965 6443
rect 9965 6409 9999 6443
rect 9999 6409 10008 6443
rect 9956 6400 10008 6409
rect 2136 6332 2188 6384
rect 3516 6264 3568 6316
rect 4804 6332 4856 6384
rect 5540 6332 5592 6384
rect 2228 6196 2280 6248
rect 1768 6060 1820 6112
rect 2228 6060 2280 6112
rect 3148 6103 3200 6112
rect 3148 6069 3157 6103
rect 3157 6069 3191 6103
rect 3191 6069 3200 6103
rect 3148 6060 3200 6069
rect 3976 6264 4028 6316
rect 4160 6264 4212 6316
rect 5080 6264 5132 6316
rect 5908 6264 5960 6316
rect 6000 6264 6052 6316
rect 6184 6264 6236 6316
rect 6552 6307 6604 6316
rect 6552 6273 6561 6307
rect 6561 6273 6595 6307
rect 6595 6273 6604 6307
rect 6552 6264 6604 6273
rect 7104 6332 7156 6384
rect 5172 6128 5224 6180
rect 5908 6171 5960 6180
rect 5908 6137 5917 6171
rect 5917 6137 5951 6171
rect 5951 6137 5960 6171
rect 6920 6196 6972 6248
rect 7196 6264 7248 6316
rect 8668 6196 8720 6248
rect 10324 6264 10376 6316
rect 5908 6128 5960 6137
rect 7012 6128 7064 6180
rect 4988 6103 5040 6112
rect 4988 6069 4997 6103
rect 4997 6069 5031 6103
rect 5031 6069 5040 6103
rect 4988 6060 5040 6069
rect 5080 6060 5132 6112
rect 8116 6103 8168 6112
rect 8116 6069 8125 6103
rect 8125 6069 8159 6103
rect 8159 6069 8168 6103
rect 8116 6060 8168 6069
rect 8300 6060 8352 6112
rect 9404 6060 9456 6112
rect 9588 6060 9640 6112
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 1584 5856 1636 5908
rect 3332 5856 3384 5908
rect 3424 5899 3476 5908
rect 3424 5865 3433 5899
rect 3433 5865 3467 5899
rect 3467 5865 3476 5899
rect 3424 5856 3476 5865
rect 4160 5856 4212 5908
rect 5080 5856 5132 5908
rect 7104 5856 7156 5908
rect 7196 5899 7248 5908
rect 7196 5865 7205 5899
rect 7205 5865 7239 5899
rect 7239 5865 7248 5899
rect 7196 5856 7248 5865
rect 3148 5695 3200 5704
rect 3148 5661 3157 5695
rect 3157 5661 3191 5695
rect 3191 5661 3200 5695
rect 3148 5652 3200 5661
rect 3700 5652 3752 5704
rect 4160 5695 4212 5704
rect 4160 5661 4169 5695
rect 4169 5661 4203 5695
rect 4203 5661 4212 5695
rect 4160 5652 4212 5661
rect 2136 5584 2188 5636
rect 2964 5584 3016 5636
rect 3332 5584 3384 5636
rect 4344 5652 4396 5704
rect 4436 5695 4488 5704
rect 4436 5661 4445 5695
rect 4445 5661 4479 5695
rect 4479 5661 4488 5695
rect 4436 5652 4488 5661
rect 4804 5652 4856 5704
rect 5540 5720 5592 5772
rect 6736 5720 6788 5772
rect 8116 5788 8168 5840
rect 8668 5763 8720 5772
rect 8668 5729 8677 5763
rect 8677 5729 8711 5763
rect 8711 5729 8720 5763
rect 8668 5720 8720 5729
rect 5448 5584 5500 5636
rect 5540 5627 5592 5636
rect 5540 5593 5549 5627
rect 5549 5593 5583 5627
rect 5583 5593 5592 5627
rect 5540 5584 5592 5593
rect 6828 5584 6880 5636
rect 3792 5559 3844 5568
rect 3792 5525 3801 5559
rect 3801 5525 3835 5559
rect 3835 5525 3844 5559
rect 3792 5516 3844 5525
rect 5632 5516 5684 5568
rect 6460 5516 6512 5568
rect 7380 5559 7432 5568
rect 7380 5525 7389 5559
rect 7389 5525 7423 5559
rect 7423 5525 7432 5559
rect 7380 5516 7432 5525
rect 9864 5652 9916 5704
rect 9956 5695 10008 5704
rect 9956 5661 9965 5695
rect 9965 5661 9999 5695
rect 9999 5661 10008 5695
rect 9956 5652 10008 5661
rect 8300 5516 8352 5568
rect 9404 5559 9456 5568
rect 9404 5525 9413 5559
rect 9413 5525 9447 5559
rect 9447 5525 9456 5559
rect 9404 5516 9456 5525
rect 9496 5516 9548 5568
rect 4874 5414 4926 5466
rect 4938 5414 4990 5466
rect 5002 5414 5054 5466
rect 5066 5414 5118 5466
rect 5130 5414 5182 5466
rect 2136 5312 2188 5364
rect 2228 5312 2280 5364
rect 3148 5312 3200 5364
rect 4436 5312 4488 5364
rect 7380 5312 7432 5364
rect 8668 5312 8720 5364
rect 9496 5312 9548 5364
rect 9956 5312 10008 5364
rect 1676 5176 1728 5228
rect 3056 5244 3108 5296
rect 5816 5287 5868 5296
rect 5816 5253 5825 5287
rect 5825 5253 5859 5287
rect 5859 5253 5868 5287
rect 5816 5244 5868 5253
rect 8392 5244 8444 5296
rect 9220 5244 9272 5296
rect 4712 5108 4764 5160
rect 5448 5108 5500 5160
rect 7012 5108 7064 5160
rect 7472 5108 7524 5160
rect 8760 5219 8812 5228
rect 8760 5185 8769 5219
rect 8769 5185 8803 5219
rect 8803 5185 8812 5219
rect 8760 5176 8812 5185
rect 9588 5176 9640 5228
rect 4620 5040 4672 5092
rect 1584 5015 1636 5024
rect 1584 4981 1593 5015
rect 1593 4981 1627 5015
rect 1627 4981 1636 5015
rect 1584 4972 1636 4981
rect 2044 5015 2096 5024
rect 2044 4981 2053 5015
rect 2053 4981 2087 5015
rect 2087 4981 2096 5015
rect 2044 4972 2096 4981
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 1584 4768 1636 4820
rect 2136 4768 2188 4820
rect 5264 4768 5316 4820
rect 5724 4768 5776 4820
rect 6828 4768 6880 4820
rect 8392 4768 8444 4820
rect 8760 4811 8812 4820
rect 8760 4777 8769 4811
rect 8769 4777 8803 4811
rect 8803 4777 8812 4811
rect 8760 4768 8812 4777
rect 9404 4768 9456 4820
rect 4620 4632 4672 4684
rect 6736 4675 6788 4684
rect 6736 4641 6745 4675
rect 6745 4641 6779 4675
rect 6779 4641 6788 4675
rect 6736 4632 6788 4641
rect 1952 4607 2004 4616
rect 1952 4573 1961 4607
rect 1961 4573 1995 4607
rect 1995 4573 2004 4607
rect 1952 4564 2004 4573
rect 7012 4675 7064 4684
rect 7012 4641 7021 4675
rect 7021 4641 7055 4675
rect 7055 4641 7064 4675
rect 7012 4632 7064 4641
rect 1032 4496 1084 4548
rect 8392 4564 8444 4616
rect 4528 4539 4580 4548
rect 4528 4505 4537 4539
rect 4537 4505 4571 4539
rect 4571 4505 4580 4539
rect 4528 4496 4580 4505
rect 1584 4471 1636 4480
rect 1584 4437 1593 4471
rect 1593 4437 1627 4471
rect 1627 4437 1636 4471
rect 1584 4428 1636 4437
rect 6092 4471 6144 4480
rect 6092 4437 6101 4471
rect 6101 4437 6135 4471
rect 6135 4437 6144 4471
rect 6092 4428 6144 4437
rect 4874 4326 4926 4378
rect 4938 4326 4990 4378
rect 5002 4326 5054 4378
rect 5066 4326 5118 4378
rect 5130 4326 5182 4378
rect 1492 4267 1544 4276
rect 1492 4233 1501 4267
rect 1501 4233 1535 4267
rect 1535 4233 1544 4267
rect 1492 4224 1544 4233
rect 1952 4224 2004 4276
rect 6460 4199 6512 4208
rect 6460 4165 6469 4199
rect 6469 4165 6503 4199
rect 6503 4165 6512 4199
rect 6460 4156 6512 4165
rect 1584 4088 1636 4140
rect 1952 4131 2004 4140
rect 1952 4097 1961 4131
rect 1961 4097 1995 4131
rect 1995 4097 2004 4131
rect 1952 4088 2004 4097
rect 3792 4020 3844 4072
rect 6092 4088 6144 4140
rect 4528 4020 4580 4072
rect 4804 4063 4856 4072
rect 4804 4029 4813 4063
rect 4813 4029 4847 4063
rect 4847 4029 4856 4063
rect 4804 4020 4856 4029
rect 5540 4020 5592 4072
rect 5724 4063 5776 4072
rect 5724 4029 5733 4063
rect 5733 4029 5767 4063
rect 5767 4029 5776 4063
rect 5724 4020 5776 4029
rect 6828 4020 6880 4072
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 5540 3612 5592 3664
rect 8484 3612 8536 3664
rect 1676 3519 1728 3528
rect 1676 3485 1685 3519
rect 1685 3485 1719 3519
rect 1719 3485 1728 3519
rect 1676 3476 1728 3485
rect 4068 3476 4120 3528
rect 6092 3544 6144 3596
rect 5724 3408 5776 3460
rect 1216 3340 1268 3392
rect 4804 3383 4856 3392
rect 4804 3349 4813 3383
rect 4813 3349 4847 3383
rect 4847 3349 4856 3383
rect 4804 3340 4856 3349
rect 5540 3340 5592 3392
rect 5632 3340 5684 3392
rect 6000 3340 6052 3392
rect 4874 3238 4926 3290
rect 4938 3238 4990 3290
rect 5002 3238 5054 3290
rect 5066 3238 5118 3290
rect 5130 3238 5182 3290
rect 1676 3136 1728 3188
rect 1400 3043 1452 3052
rect 1400 3009 1409 3043
rect 1409 3009 1443 3043
rect 1443 3009 1452 3043
rect 1400 3000 1452 3009
rect 2964 3043 3016 3052
rect 2964 3009 2973 3043
rect 2973 3009 3007 3043
rect 3007 3009 3016 3043
rect 2964 3000 3016 3009
rect 3884 3136 3936 3188
rect 5724 3136 5776 3188
rect 3240 2975 3292 2984
rect 3240 2941 3249 2975
rect 3249 2941 3283 2975
rect 3283 2941 3292 2975
rect 3240 2932 3292 2941
rect 4068 3000 4120 3052
rect 6000 3111 6052 3120
rect 6000 3077 6009 3111
rect 6009 3077 6043 3111
rect 6043 3077 6052 3111
rect 6000 3068 6052 3077
rect 7840 3136 7892 3188
rect 5632 3043 5684 3052
rect 5632 3009 5641 3043
rect 5641 3009 5675 3043
rect 5675 3009 5684 3043
rect 5632 3000 5684 3009
rect 3516 2932 3568 2984
rect 3976 2975 4028 2984
rect 3976 2941 3985 2975
rect 3985 2941 4019 2975
rect 4019 2941 4028 2975
rect 3976 2932 4028 2941
rect 6092 2932 6144 2984
rect 2596 2796 2648 2848
rect 3424 2796 3476 2848
rect 3608 2839 3660 2848
rect 3608 2805 3617 2839
rect 3617 2805 3651 2839
rect 3651 2805 3660 2839
rect 3608 2796 3660 2805
rect 3884 2796 3936 2848
rect 5540 2796 5592 2848
rect 6000 2839 6052 2848
rect 6000 2805 6009 2839
rect 6009 2805 6043 2839
rect 6043 2805 6052 2839
rect 6000 2796 6052 2805
rect 6368 2839 6420 2848
rect 6368 2805 6377 2839
rect 6377 2805 6411 2839
rect 6411 2805 6420 2839
rect 6368 2796 6420 2805
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 2964 2592 3016 2644
rect 6000 2635 6052 2644
rect 6000 2601 6009 2635
rect 6009 2601 6043 2635
rect 6043 2601 6052 2635
rect 6000 2592 6052 2601
rect 3240 2456 3292 2508
rect 3424 2499 3476 2508
rect 3424 2465 3433 2499
rect 3433 2465 3467 2499
rect 3467 2465 3476 2499
rect 3424 2456 3476 2465
rect 2044 2431 2096 2440
rect 2044 2397 2053 2431
rect 2053 2397 2087 2431
rect 2087 2397 2096 2431
rect 2044 2388 2096 2397
rect 3516 2431 3568 2440
rect 3516 2397 3525 2431
rect 3525 2397 3559 2431
rect 3559 2397 3568 2431
rect 3516 2388 3568 2397
rect 3608 2388 3660 2440
rect 4620 2431 4672 2440
rect 4620 2397 4629 2431
rect 4629 2397 4663 2431
rect 4663 2397 4672 2431
rect 4620 2388 4672 2397
rect 4804 2388 4856 2440
rect 5908 2388 5960 2440
rect 6368 2388 6420 2440
rect 7840 2431 7892 2440
rect 7840 2397 7849 2431
rect 7849 2397 7883 2431
rect 7883 2397 7892 2431
rect 7840 2388 7892 2397
rect 8484 2431 8536 2440
rect 8484 2397 8493 2431
rect 8493 2397 8527 2431
rect 8527 2397 8536 2431
rect 8484 2388 8536 2397
rect 3240 2252 3292 2304
rect 4804 2252 4856 2304
rect 6460 2252 6512 2304
rect 7104 2252 7156 2304
rect 7748 2252 7800 2304
rect 8392 2252 8444 2304
rect 4874 2150 4926 2202
rect 4938 2150 4990 2202
rect 5002 2150 5054 2202
rect 5066 2150 5118 2202
rect 5130 2150 5182 2202
<< metal2 >>
rect 5814 12884 5870 13684
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 5828 11354 5856 12884
rect 5816 11348 5868 11354
rect 5816 11290 5868 11296
rect 6092 11280 6144 11286
rect 6092 11222 6144 11228
rect 4804 11212 4856 11218
rect 4804 11154 4856 11160
rect 4712 11008 4764 11014
rect 4712 10950 4764 10956
rect 4160 10668 4212 10674
rect 4160 10610 4212 10616
rect 2780 10600 2832 10606
rect 2780 10542 2832 10548
rect 3056 10600 3108 10606
rect 4172 10554 4200 10610
rect 3056 10542 3108 10548
rect 2792 10198 2820 10542
rect 3068 10266 3096 10542
rect 4080 10526 4200 10554
rect 3516 10464 3568 10470
rect 3516 10406 3568 10412
rect 3056 10260 3108 10266
rect 3056 10202 3108 10208
rect 2780 10192 2832 10198
rect 2780 10134 2832 10140
rect 2792 9586 2820 10134
rect 3528 10130 3556 10406
rect 4080 10146 4108 10526
rect 4528 10464 4580 10470
rect 4580 10424 4660 10452
rect 4528 10406 4580 10412
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 4344 10260 4396 10266
rect 4344 10202 4396 10208
rect 3516 10124 3568 10130
rect 4080 10118 4200 10146
rect 3516 10066 3568 10072
rect 2872 9988 2924 9994
rect 2872 9930 2924 9936
rect 2780 9580 2832 9586
rect 2780 9522 2832 9528
rect 1400 8492 1452 8498
rect 1400 8434 1452 8440
rect 1412 6361 1440 8434
rect 1676 8356 1728 8362
rect 1676 8298 1728 8304
rect 1584 7336 1636 7342
rect 1584 7278 1636 7284
rect 1492 6928 1544 6934
rect 1490 6896 1492 6905
rect 1544 6896 1546 6905
rect 1490 6831 1546 6840
rect 1398 6352 1454 6361
rect 1398 6287 1454 6296
rect 1596 5914 1624 7278
rect 1584 5908 1636 5914
rect 1584 5850 1636 5856
rect 1030 5536 1086 5545
rect 1030 5471 1086 5480
rect 1044 4554 1072 5471
rect 1688 5234 1716 8298
rect 2792 7954 2820 9522
rect 2884 8498 2912 9930
rect 2964 9920 3016 9926
rect 2964 9862 3016 9868
rect 3148 9920 3200 9926
rect 3148 9862 3200 9868
rect 2976 9178 3004 9862
rect 3160 9654 3188 9862
rect 3148 9648 3200 9654
rect 3148 9590 3200 9596
rect 4172 9586 4200 10118
rect 4356 10062 4384 10202
rect 4632 10062 4660 10424
rect 4724 10130 4752 10950
rect 4816 10266 4844 11154
rect 5816 11144 5868 11150
rect 5816 11086 5868 11092
rect 5264 11076 5316 11082
rect 5264 11018 5316 11024
rect 5632 11076 5684 11082
rect 5632 11018 5684 11024
rect 4874 10908 5182 10917
rect 4874 10906 4880 10908
rect 4936 10906 4960 10908
rect 5016 10906 5040 10908
rect 5096 10906 5120 10908
rect 5176 10906 5182 10908
rect 4936 10854 4938 10906
rect 5118 10854 5120 10906
rect 4874 10852 4880 10854
rect 4936 10852 4960 10854
rect 5016 10852 5040 10854
rect 5096 10852 5120 10854
rect 5176 10852 5182 10854
rect 4874 10843 5182 10852
rect 5080 10668 5132 10674
rect 5080 10610 5132 10616
rect 5092 10470 5120 10610
rect 5080 10464 5132 10470
rect 5080 10406 5132 10412
rect 4804 10260 4856 10266
rect 4804 10202 4856 10208
rect 4712 10124 4764 10130
rect 4712 10066 4764 10072
rect 4252 10056 4304 10062
rect 4252 9998 4304 10004
rect 4344 10056 4396 10062
rect 4620 10056 4672 10062
rect 4344 9998 4396 10004
rect 4448 10004 4620 10010
rect 4448 9998 4672 10004
rect 4160 9580 4212 9586
rect 4160 9522 4212 9528
rect 4264 9466 4292 9998
rect 4448 9982 4660 9998
rect 4448 9926 4476 9982
rect 4344 9920 4396 9926
rect 4344 9862 4396 9868
rect 4436 9920 4488 9926
rect 4436 9862 4488 9868
rect 4528 9920 4580 9926
rect 4528 9862 4580 9868
rect 4356 9586 4384 9862
rect 4540 9722 4568 9862
rect 4528 9716 4580 9722
rect 4528 9658 4580 9664
rect 4632 9654 4660 9982
rect 4874 9820 5182 9829
rect 4874 9818 4880 9820
rect 4936 9818 4960 9820
rect 5016 9818 5040 9820
rect 5096 9818 5120 9820
rect 5176 9818 5182 9820
rect 4936 9766 4938 9818
rect 5118 9766 5120 9818
rect 4874 9764 4880 9766
rect 4936 9764 4960 9766
rect 5016 9764 5040 9766
rect 5096 9764 5120 9766
rect 5176 9764 5182 9766
rect 4874 9755 5182 9764
rect 5276 9654 5304 11018
rect 5644 10742 5672 11018
rect 5828 10810 5856 11086
rect 5908 11008 5960 11014
rect 5908 10950 5960 10956
rect 5816 10804 5868 10810
rect 5816 10746 5868 10752
rect 5632 10736 5684 10742
rect 5632 10678 5684 10684
rect 5644 10606 5672 10678
rect 5632 10600 5684 10606
rect 5632 10542 5684 10548
rect 5540 10192 5592 10198
rect 5540 10134 5592 10140
rect 5356 10124 5408 10130
rect 5356 10066 5408 10072
rect 5368 9722 5396 10066
rect 5552 10062 5580 10134
rect 5540 10056 5592 10062
rect 5540 9998 5592 10004
rect 5356 9716 5408 9722
rect 5356 9658 5408 9664
rect 5552 9654 5580 9998
rect 5644 9926 5672 10542
rect 5920 10470 5948 10950
rect 6104 10810 6132 11222
rect 6736 11144 6788 11150
rect 6736 11086 6788 11092
rect 6000 10804 6052 10810
rect 6000 10746 6052 10752
rect 6092 10804 6144 10810
rect 6092 10746 6144 10752
rect 5908 10464 5960 10470
rect 5908 10406 5960 10412
rect 5920 10130 5948 10406
rect 5908 10124 5960 10130
rect 5908 10066 5960 10072
rect 5816 9988 5868 9994
rect 5816 9930 5868 9936
rect 5908 9988 5960 9994
rect 5908 9930 5960 9936
rect 5632 9920 5684 9926
rect 5632 9862 5684 9868
rect 5828 9722 5856 9930
rect 5816 9716 5868 9722
rect 5816 9658 5868 9664
rect 4620 9648 4672 9654
rect 5264 9648 5316 9654
rect 4620 9590 4672 9596
rect 4710 9616 4766 9625
rect 4344 9580 4396 9586
rect 4344 9522 4396 9528
rect 4080 9450 4292 9466
rect 4080 9444 4304 9450
rect 4080 9438 4252 9444
rect 2964 9172 3016 9178
rect 2964 9114 3016 9120
rect 4080 9058 4108 9438
rect 4252 9386 4304 9392
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 4080 9042 4200 9058
rect 4080 9036 4212 9042
rect 4080 9030 4160 9036
rect 4160 8978 4212 8984
rect 4632 8838 4660 9590
rect 5264 9590 5316 9596
rect 5540 9648 5592 9654
rect 5540 9590 5592 9596
rect 4710 9551 4766 9560
rect 4620 8832 4672 8838
rect 4620 8774 4672 8780
rect 3976 8628 4028 8634
rect 3976 8570 4028 8576
rect 3424 8560 3476 8566
rect 3424 8502 3476 8508
rect 3606 8528 3662 8537
rect 2872 8492 2924 8498
rect 2872 8434 2924 8440
rect 3240 8492 3292 8498
rect 3240 8434 3292 8440
rect 2964 8356 3016 8362
rect 2964 8298 3016 8304
rect 2872 8288 2924 8294
rect 2872 8230 2924 8236
rect 2780 7948 2832 7954
rect 2780 7890 2832 7896
rect 2780 7812 2832 7818
rect 2780 7754 2832 7760
rect 2792 7342 2820 7754
rect 1768 7336 1820 7342
rect 1768 7278 1820 7284
rect 2780 7336 2832 7342
rect 2780 7278 2832 7284
rect 1780 6798 1808 7278
rect 2228 7200 2280 7206
rect 2228 7142 2280 7148
rect 1768 6792 1820 6798
rect 1768 6734 1820 6740
rect 2042 6760 2098 6769
rect 1780 6118 1808 6734
rect 2042 6695 2044 6704
rect 2096 6695 2098 6704
rect 2044 6666 2096 6672
rect 1768 6112 1820 6118
rect 1768 6054 1820 6060
rect 1676 5228 1728 5234
rect 1676 5170 1728 5176
rect 2056 5030 2084 6666
rect 2136 6384 2188 6390
rect 2136 6326 2188 6332
rect 2148 5642 2176 6326
rect 2240 6254 2268 7142
rect 2884 7018 2912 8230
rect 2792 7002 2912 7018
rect 2780 6996 2912 7002
rect 2832 6990 2912 6996
rect 2780 6938 2832 6944
rect 2228 6248 2280 6254
rect 2228 6190 2280 6196
rect 2228 6112 2280 6118
rect 2228 6054 2280 6060
rect 2136 5636 2188 5642
rect 2136 5578 2188 5584
rect 2148 5370 2176 5578
rect 2240 5370 2268 6054
rect 2976 5642 3004 8298
rect 3252 8090 3280 8434
rect 3240 8084 3292 8090
rect 3240 8026 3292 8032
rect 3056 7472 3108 7478
rect 3056 7414 3108 7420
rect 3068 7324 3096 7414
rect 3148 7336 3200 7342
rect 3068 7296 3148 7324
rect 3068 6730 3096 7296
rect 3148 7278 3200 7284
rect 3436 6866 3464 8502
rect 3516 8492 3568 8498
rect 3606 8463 3662 8472
rect 3884 8492 3936 8498
rect 3516 8434 3568 8440
rect 3528 7886 3556 8434
rect 3620 8430 3648 8463
rect 3884 8434 3936 8440
rect 3608 8424 3660 8430
rect 3660 8384 3740 8412
rect 3608 8366 3660 8372
rect 3516 7880 3568 7886
rect 3516 7822 3568 7828
rect 3608 7880 3660 7886
rect 3608 7822 3660 7828
rect 3424 6860 3476 6866
rect 3424 6802 3476 6808
rect 3528 6798 3556 7822
rect 3620 7002 3648 7822
rect 3608 6996 3660 7002
rect 3608 6938 3660 6944
rect 3516 6792 3568 6798
rect 3516 6734 3568 6740
rect 3056 6724 3108 6730
rect 3056 6666 3108 6672
rect 3332 6724 3384 6730
rect 3332 6666 3384 6672
rect 2964 5636 3016 5642
rect 2964 5578 3016 5584
rect 2136 5364 2188 5370
rect 2136 5306 2188 5312
rect 2228 5364 2280 5370
rect 2228 5306 2280 5312
rect 1584 5024 1636 5030
rect 1584 4966 1636 4972
rect 2044 5024 2096 5030
rect 2044 4966 2096 4972
rect 1490 4856 1546 4865
rect 1596 4826 1624 4966
rect 2148 4826 2176 5306
rect 3068 5302 3096 6666
rect 3148 6112 3200 6118
rect 3148 6054 3200 6060
rect 3160 5817 3188 6054
rect 3344 5914 3372 6666
rect 3424 6656 3476 6662
rect 3424 6598 3476 6604
rect 3436 5914 3464 6598
rect 3516 6316 3568 6322
rect 3516 6258 3568 6264
rect 3528 6225 3556 6258
rect 3514 6216 3570 6225
rect 3514 6151 3570 6160
rect 3332 5908 3384 5914
rect 3332 5850 3384 5856
rect 3424 5908 3476 5914
rect 3424 5850 3476 5856
rect 3146 5808 3202 5817
rect 3146 5743 3202 5752
rect 3148 5704 3200 5710
rect 3148 5646 3200 5652
rect 3160 5370 3188 5646
rect 3344 5642 3372 5850
rect 3712 5710 3740 8384
rect 3896 8294 3924 8434
rect 3884 8288 3936 8294
rect 3884 8230 3936 8236
rect 3896 7954 3924 8230
rect 3884 7948 3936 7954
rect 3884 7890 3936 7896
rect 3792 7880 3844 7886
rect 3792 7822 3844 7828
rect 3804 7546 3832 7822
rect 3792 7540 3844 7546
rect 3792 7482 3844 7488
rect 3896 7002 3924 7890
rect 3988 7886 4016 8570
rect 4068 8356 4120 8362
rect 4068 8298 4120 8304
rect 4080 7970 4108 8298
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 4620 8016 4672 8022
rect 4080 7942 4200 7970
rect 4620 7958 4672 7964
rect 4172 7886 4200 7942
rect 3976 7880 4028 7886
rect 3976 7822 4028 7828
rect 4160 7880 4212 7886
rect 4160 7822 4212 7828
rect 4068 7744 4120 7750
rect 4068 7686 4120 7692
rect 3884 6996 3936 7002
rect 4080 6984 4108 7686
rect 4632 7410 4660 7958
rect 4724 7478 4752 9551
rect 4874 8732 5182 8741
rect 4874 8730 4880 8732
rect 4936 8730 4960 8732
rect 5016 8730 5040 8732
rect 5096 8730 5120 8732
rect 5176 8730 5182 8732
rect 4936 8678 4938 8730
rect 5118 8678 5120 8730
rect 4874 8676 4880 8678
rect 4936 8676 4960 8678
rect 5016 8676 5040 8678
rect 5096 8676 5120 8678
rect 5176 8676 5182 8678
rect 4874 8667 5182 8676
rect 4896 8492 4948 8498
rect 4896 8434 4948 8440
rect 4804 8288 4856 8294
rect 4804 8230 4856 8236
rect 4816 8090 4844 8230
rect 4804 8084 4856 8090
rect 4804 8026 4856 8032
rect 4804 7948 4856 7954
rect 4804 7890 4856 7896
rect 4712 7472 4764 7478
rect 4712 7414 4764 7420
rect 4620 7404 4672 7410
rect 4620 7346 4672 7352
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 4080 6956 4200 6984
rect 3884 6938 3936 6944
rect 3896 6866 3924 6938
rect 3976 6928 4028 6934
rect 3976 6870 4028 6876
rect 3884 6860 3936 6866
rect 3884 6802 3936 6808
rect 3988 6322 4016 6870
rect 4172 6798 4200 6956
rect 4160 6792 4212 6798
rect 4160 6734 4212 6740
rect 4436 6792 4488 6798
rect 4436 6734 4488 6740
rect 4172 6322 4200 6734
rect 4448 6458 4476 6734
rect 4632 6458 4660 7346
rect 4816 7206 4844 7890
rect 4908 7750 4936 8434
rect 5276 8378 5304 9590
rect 5920 9518 5948 9930
rect 6012 9586 6040 10746
rect 6644 10600 6696 10606
rect 6644 10542 6696 10548
rect 6552 10464 6604 10470
rect 6552 10406 6604 10412
rect 6184 10260 6236 10266
rect 6184 10202 6236 10208
rect 6000 9580 6052 9586
rect 6000 9522 6052 9528
rect 5632 9512 5684 9518
rect 5632 9454 5684 9460
rect 5724 9512 5776 9518
rect 5724 9454 5776 9460
rect 5908 9512 5960 9518
rect 5908 9454 5960 9460
rect 5448 9376 5500 9382
rect 5448 9318 5500 9324
rect 5356 9036 5408 9042
rect 5356 8978 5408 8984
rect 5368 8537 5396 8978
rect 5354 8528 5410 8537
rect 5354 8463 5410 8472
rect 5184 8350 5304 8378
rect 5184 7954 5212 8350
rect 5264 8288 5316 8294
rect 5264 8230 5316 8236
rect 5172 7948 5224 7954
rect 5172 7890 5224 7896
rect 5276 7886 5304 8230
rect 5356 7948 5408 7954
rect 5356 7890 5408 7896
rect 5264 7880 5316 7886
rect 5264 7822 5316 7828
rect 4896 7744 4948 7750
rect 4896 7686 4948 7692
rect 5264 7744 5316 7750
rect 5264 7686 5316 7692
rect 4874 7644 5182 7653
rect 4874 7642 4880 7644
rect 4936 7642 4960 7644
rect 5016 7642 5040 7644
rect 5096 7642 5120 7644
rect 5176 7642 5182 7644
rect 4936 7590 4938 7642
rect 5118 7590 5120 7642
rect 4874 7588 4880 7590
rect 4936 7588 4960 7590
rect 5016 7588 5040 7590
rect 5096 7588 5120 7590
rect 5176 7588 5182 7590
rect 4874 7579 5182 7588
rect 5080 7336 5132 7342
rect 5276 7324 5304 7686
rect 5368 7478 5396 7890
rect 5460 7886 5488 9318
rect 5644 8838 5672 9454
rect 5736 9178 5764 9454
rect 5724 9172 5776 9178
rect 5724 9114 5776 9120
rect 6012 8974 6040 9522
rect 6000 8968 6052 8974
rect 6000 8910 6052 8916
rect 5816 8900 5868 8906
rect 5816 8842 5868 8848
rect 5632 8832 5684 8838
rect 5632 8774 5684 8780
rect 5540 8628 5592 8634
rect 5540 8570 5592 8576
rect 5552 8090 5580 8570
rect 5632 8492 5684 8498
rect 5632 8434 5684 8440
rect 5540 8084 5592 8090
rect 5540 8026 5592 8032
rect 5448 7880 5500 7886
rect 5448 7822 5500 7828
rect 5356 7472 5408 7478
rect 5356 7414 5408 7420
rect 5132 7296 5304 7324
rect 5080 7278 5132 7284
rect 4804 7200 4856 7206
rect 4804 7142 4856 7148
rect 5092 6866 5120 7278
rect 5264 7200 5316 7206
rect 5264 7142 5316 7148
rect 5276 6866 5304 7142
rect 5368 7002 5396 7414
rect 5356 6996 5408 7002
rect 5356 6938 5408 6944
rect 5080 6860 5132 6866
rect 5080 6802 5132 6808
rect 5264 6860 5316 6866
rect 5264 6802 5316 6808
rect 4712 6656 4764 6662
rect 4712 6598 4764 6604
rect 4344 6452 4396 6458
rect 4344 6394 4396 6400
rect 4436 6452 4488 6458
rect 4436 6394 4488 6400
rect 4620 6452 4672 6458
rect 4620 6394 4672 6400
rect 4356 6361 4384 6394
rect 4342 6352 4398 6361
rect 3976 6316 4028 6322
rect 3976 6258 4028 6264
rect 4160 6316 4212 6322
rect 4342 6287 4398 6296
rect 4160 6258 4212 6264
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 4160 5908 4212 5914
rect 4160 5850 4212 5856
rect 4172 5710 4200 5850
rect 4250 5808 4306 5817
rect 4250 5743 4306 5752
rect 3700 5704 3752 5710
rect 3700 5646 3752 5652
rect 4160 5704 4212 5710
rect 4264 5692 4292 5743
rect 4344 5704 4396 5710
rect 4264 5664 4344 5692
rect 4160 5646 4212 5652
rect 4344 5646 4396 5652
rect 4436 5704 4488 5710
rect 4436 5646 4488 5652
rect 3332 5636 3384 5642
rect 3332 5578 3384 5584
rect 3792 5568 3844 5574
rect 3792 5510 3844 5516
rect 3148 5364 3200 5370
rect 3148 5306 3200 5312
rect 3056 5296 3108 5302
rect 3056 5238 3108 5244
rect 1490 4791 1546 4800
rect 1584 4820 1636 4826
rect 1032 4548 1084 4554
rect 1032 4490 1084 4496
rect 1504 4282 1532 4791
rect 1584 4762 1636 4768
rect 2136 4820 2188 4826
rect 2136 4762 2188 4768
rect 1952 4616 2004 4622
rect 1952 4558 2004 4564
rect 1584 4480 1636 4486
rect 1584 4422 1636 4428
rect 1492 4276 1544 4282
rect 1492 4218 1544 4224
rect 1596 4146 1624 4422
rect 1964 4282 1992 4558
rect 1952 4276 2004 4282
rect 1952 4218 2004 4224
rect 1950 4176 2006 4185
rect 1584 4140 1636 4146
rect 1950 4111 1952 4120
rect 1584 4082 1636 4088
rect 2004 4111 2006 4120
rect 1952 4082 2004 4088
rect 3804 4078 3832 5510
rect 4448 5370 4476 5646
rect 4436 5364 4488 5370
rect 4436 5306 4488 5312
rect 4724 5166 4752 6598
rect 4874 6556 5182 6565
rect 4874 6554 4880 6556
rect 4936 6554 4960 6556
rect 5016 6554 5040 6556
rect 5096 6554 5120 6556
rect 5176 6554 5182 6556
rect 4936 6502 4938 6554
rect 5118 6502 5120 6554
rect 4874 6500 4880 6502
rect 4936 6500 4960 6502
rect 5016 6500 5040 6502
rect 5096 6500 5120 6502
rect 5176 6500 5182 6502
rect 4874 6491 5182 6500
rect 4896 6452 4948 6458
rect 4896 6394 4948 6400
rect 4804 6384 4856 6390
rect 4804 6326 4856 6332
rect 4816 5710 4844 6326
rect 4908 6089 4936 6394
rect 5276 6338 5304 6802
rect 5356 6792 5408 6798
rect 5408 6752 5488 6780
rect 5356 6734 5408 6740
rect 5460 6372 5488 6752
rect 5540 6724 5592 6730
rect 5540 6666 5592 6672
rect 5552 6474 5580 6666
rect 5644 6662 5672 8434
rect 5724 8288 5776 8294
rect 5724 8230 5776 8236
rect 5736 7342 5764 8230
rect 5724 7336 5776 7342
rect 5724 7278 5776 7284
rect 5828 7206 5856 8842
rect 6012 8498 6040 8910
rect 6090 8528 6146 8537
rect 6000 8492 6052 8498
rect 6090 8463 6092 8472
rect 6000 8434 6052 8440
rect 6144 8463 6146 8472
rect 6092 8434 6144 8440
rect 6012 7546 6040 8434
rect 6000 7540 6052 7546
rect 6000 7482 6052 7488
rect 6000 7404 6052 7410
rect 6000 7346 6052 7352
rect 5816 7200 5868 7206
rect 5816 7142 5868 7148
rect 5722 6760 5778 6769
rect 5722 6695 5778 6704
rect 5632 6656 5684 6662
rect 5632 6598 5684 6604
rect 5552 6446 5672 6474
rect 5736 6458 5764 6695
rect 5540 6384 5592 6390
rect 5460 6344 5540 6372
rect 5092 6322 5304 6338
rect 5540 6326 5592 6332
rect 5080 6316 5304 6322
rect 5132 6310 5304 6316
rect 5080 6258 5132 6264
rect 5538 6216 5594 6225
rect 5172 6180 5224 6186
rect 5224 6140 5304 6168
rect 5538 6151 5594 6160
rect 5172 6122 5224 6128
rect 4988 6112 5040 6118
rect 4894 6080 4950 6089
rect 4988 6054 5040 6060
rect 5080 6112 5132 6118
rect 5080 6054 5132 6060
rect 4894 6015 4950 6024
rect 4804 5704 4856 5710
rect 4804 5646 4856 5652
rect 5000 5556 5028 6054
rect 5092 5914 5120 6054
rect 5080 5908 5132 5914
rect 5080 5850 5132 5856
rect 4816 5528 5028 5556
rect 4712 5160 4764 5166
rect 4712 5102 4764 5108
rect 4620 5092 4672 5098
rect 4620 5034 4672 5040
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 4632 4690 4660 5034
rect 4620 4684 4672 4690
rect 4620 4626 4672 4632
rect 4528 4548 4580 4554
rect 4528 4490 4580 4496
rect 4540 4078 4568 4490
rect 4816 4078 4844 5528
rect 4874 5468 5182 5477
rect 4874 5466 4880 5468
rect 4936 5466 4960 5468
rect 5016 5466 5040 5468
rect 5096 5466 5120 5468
rect 5176 5466 5182 5468
rect 4936 5414 4938 5466
rect 5118 5414 5120 5466
rect 4874 5412 4880 5414
rect 4936 5412 4960 5414
rect 5016 5412 5040 5414
rect 5096 5412 5120 5414
rect 5176 5412 5182 5414
rect 4874 5403 5182 5412
rect 5276 4826 5304 6140
rect 5552 5778 5580 6151
rect 5540 5772 5592 5778
rect 5540 5714 5592 5720
rect 5448 5636 5500 5642
rect 5448 5578 5500 5584
rect 5540 5636 5592 5642
rect 5540 5578 5592 5584
rect 5460 5166 5488 5578
rect 5448 5160 5500 5166
rect 5448 5102 5500 5108
rect 5264 4820 5316 4826
rect 5264 4762 5316 4768
rect 4874 4380 5182 4389
rect 4874 4378 4880 4380
rect 4936 4378 4960 4380
rect 5016 4378 5040 4380
rect 5096 4378 5120 4380
rect 5176 4378 5182 4380
rect 4936 4326 4938 4378
rect 5118 4326 5120 4378
rect 4874 4324 4880 4326
rect 4936 4324 4960 4326
rect 5016 4324 5040 4326
rect 5096 4324 5120 4326
rect 5176 4324 5182 4326
rect 4874 4315 5182 4324
rect 5552 4078 5580 5578
rect 5644 5574 5672 6446
rect 5724 6452 5776 6458
rect 5724 6394 5776 6400
rect 5632 5568 5684 5574
rect 5632 5510 5684 5516
rect 5828 5302 5856 7142
rect 6012 7002 6040 7346
rect 6000 6996 6052 7002
rect 6000 6938 6052 6944
rect 6012 6730 6040 6938
rect 6000 6724 6052 6730
rect 6000 6666 6052 6672
rect 5906 6352 5962 6361
rect 5906 6287 5908 6296
rect 5960 6287 5962 6296
rect 6000 6316 6052 6322
rect 5908 6258 5960 6264
rect 6104 6304 6132 8434
rect 6196 6322 6224 10202
rect 6564 9654 6592 10406
rect 6552 9648 6604 9654
rect 6552 9590 6604 9596
rect 6368 9580 6420 9586
rect 6368 9522 6420 9528
rect 6380 8838 6408 9522
rect 6368 8832 6420 8838
rect 6368 8774 6420 8780
rect 6656 8634 6684 10542
rect 6644 8628 6696 8634
rect 6644 8570 6696 8576
rect 6748 8514 6776 11086
rect 6920 10056 6972 10062
rect 6920 9998 6972 10004
rect 6932 9738 6960 9998
rect 6932 9722 7052 9738
rect 6932 9716 7064 9722
rect 6932 9710 7012 9716
rect 7012 9658 7064 9664
rect 7024 9382 7052 9658
rect 7012 9376 7064 9382
rect 7012 9318 7064 9324
rect 6828 8832 6880 8838
rect 6828 8774 6880 8780
rect 6656 8486 6776 8514
rect 6840 8498 6868 8774
rect 6828 8492 6880 8498
rect 6552 7540 6604 7546
rect 6552 7482 6604 7488
rect 6460 7404 6512 7410
rect 6460 7346 6512 7352
rect 6368 6996 6420 7002
rect 6368 6938 6420 6944
rect 6380 6798 6408 6938
rect 6368 6792 6420 6798
rect 6368 6734 6420 6740
rect 6368 6656 6420 6662
rect 6472 6610 6500 7346
rect 6564 7002 6592 7482
rect 6552 6996 6604 7002
rect 6552 6938 6604 6944
rect 6552 6860 6604 6866
rect 6552 6802 6604 6808
rect 6420 6604 6500 6610
rect 6368 6598 6500 6604
rect 6380 6582 6500 6598
rect 6564 6322 6592 6802
rect 6656 6730 6684 8486
rect 6828 8434 6880 8440
rect 6840 7954 6868 8434
rect 6828 7948 6880 7954
rect 6828 7890 6880 7896
rect 6840 7410 6868 7890
rect 7024 7546 7052 9318
rect 9404 8968 9456 8974
rect 9404 8910 9456 8916
rect 8944 8832 8996 8838
rect 8944 8774 8996 8780
rect 8956 8634 8984 8774
rect 8944 8628 8996 8634
rect 8944 8570 8996 8576
rect 9416 8566 9444 8910
rect 8392 8560 8444 8566
rect 8392 8502 8444 8508
rect 9036 8560 9088 8566
rect 9036 8502 9088 8508
rect 9404 8560 9456 8566
rect 9404 8502 9456 8508
rect 8404 7954 8432 8502
rect 8484 8356 8536 8362
rect 8484 8298 8536 8304
rect 8392 7948 8444 7954
rect 8392 7890 8444 7896
rect 7196 7812 7248 7818
rect 7196 7754 7248 7760
rect 7208 7546 7236 7754
rect 7012 7540 7064 7546
rect 7012 7482 7064 7488
rect 7196 7540 7248 7546
rect 7196 7482 7248 7488
rect 6828 7404 6880 7410
rect 6828 7346 6880 7352
rect 6920 6792 6972 6798
rect 6920 6734 6972 6740
rect 6644 6724 6696 6730
rect 6644 6666 6696 6672
rect 6656 6458 6684 6666
rect 6644 6452 6696 6458
rect 6644 6394 6696 6400
rect 6052 6276 6132 6304
rect 6000 6258 6052 6264
rect 6104 6225 6132 6276
rect 6184 6316 6236 6322
rect 6184 6258 6236 6264
rect 6552 6316 6604 6322
rect 6552 6258 6604 6264
rect 6932 6254 6960 6734
rect 7012 6656 7064 6662
rect 7012 6598 7064 6604
rect 6920 6248 6972 6254
rect 6090 6216 6146 6225
rect 5908 6180 5960 6186
rect 6920 6190 6972 6196
rect 7024 6186 7052 6598
rect 7104 6384 7156 6390
rect 7104 6326 7156 6332
rect 6090 6151 6146 6160
rect 7012 6180 7064 6186
rect 5908 6122 5960 6128
rect 7012 6122 7064 6128
rect 5920 6089 5948 6122
rect 5906 6080 5962 6089
rect 5906 6015 5962 6024
rect 7116 5914 7144 6326
rect 7196 6316 7248 6322
rect 7196 6258 7248 6264
rect 7208 5914 7236 6258
rect 7470 6216 7526 6225
rect 7470 6151 7526 6160
rect 7104 5908 7156 5914
rect 7104 5850 7156 5856
rect 7196 5908 7248 5914
rect 7196 5850 7248 5856
rect 6736 5772 6788 5778
rect 6736 5714 6788 5720
rect 6460 5568 6512 5574
rect 6460 5510 6512 5516
rect 5816 5296 5868 5302
rect 5816 5238 5868 5244
rect 5724 4820 5776 4826
rect 5724 4762 5776 4768
rect 5736 4078 5764 4762
rect 6092 4480 6144 4486
rect 6092 4422 6144 4428
rect 6104 4146 6132 4422
rect 6472 4214 6500 5510
rect 6748 4690 6776 5714
rect 6828 5636 6880 5642
rect 6828 5578 6880 5584
rect 6840 4826 6868 5578
rect 7380 5568 7432 5574
rect 7380 5510 7432 5516
rect 7392 5370 7420 5510
rect 7380 5364 7432 5370
rect 7380 5306 7432 5312
rect 7484 5166 7512 6151
rect 8116 6112 8168 6118
rect 8116 6054 8168 6060
rect 8300 6112 8352 6118
rect 8300 6054 8352 6060
rect 8128 5846 8156 6054
rect 8116 5840 8168 5846
rect 8116 5782 8168 5788
rect 8312 5574 8340 6054
rect 8300 5568 8352 5574
rect 8300 5510 8352 5516
rect 8404 5302 8432 7890
rect 8496 7002 8524 8298
rect 8944 7880 8996 7886
rect 8944 7822 8996 7828
rect 8668 7744 8720 7750
rect 8668 7686 8720 7692
rect 8484 6996 8536 7002
rect 8484 6938 8536 6944
rect 8680 6866 8708 7686
rect 8956 7206 8984 7822
rect 9048 7342 9076 8502
rect 9220 8492 9272 8498
rect 9220 8434 9272 8440
rect 9128 7948 9180 7954
rect 9128 7890 9180 7896
rect 9140 7546 9168 7890
rect 9232 7818 9260 8434
rect 9312 8288 9364 8294
rect 9312 8230 9364 8236
rect 9220 7812 9272 7818
rect 9220 7754 9272 7760
rect 9128 7540 9180 7546
rect 9128 7482 9180 7488
rect 9324 7410 9352 8230
rect 9416 7886 9444 8502
rect 9496 8492 9548 8498
rect 9496 8434 9548 8440
rect 9680 8492 9732 8498
rect 9680 8434 9732 8440
rect 9404 7880 9456 7886
rect 9404 7822 9456 7828
rect 9312 7404 9364 7410
rect 9312 7346 9364 7352
rect 9036 7336 9088 7342
rect 9416 7290 9444 7822
rect 9508 7410 9536 8434
rect 9588 7744 9640 7750
rect 9588 7686 9640 7692
rect 9496 7404 9548 7410
rect 9496 7346 9548 7352
rect 9036 7278 9088 7284
rect 9324 7262 9444 7290
rect 8944 7200 8996 7206
rect 8944 7142 8996 7148
rect 8668 6860 8720 6866
rect 8668 6802 8720 6808
rect 8956 6798 8984 7142
rect 9324 6798 9352 7262
rect 9508 7018 9536 7346
rect 9416 6990 9536 7018
rect 8944 6792 8996 6798
rect 8944 6734 8996 6740
rect 9312 6792 9364 6798
rect 9312 6734 9364 6740
rect 8944 6656 8996 6662
rect 8944 6598 8996 6604
rect 9220 6656 9272 6662
rect 9220 6598 9272 6604
rect 8956 6458 8984 6598
rect 8944 6452 8996 6458
rect 8944 6394 8996 6400
rect 8668 6248 8720 6254
rect 8668 6190 8720 6196
rect 8680 5778 8708 6190
rect 8668 5772 8720 5778
rect 8668 5714 8720 5720
rect 8680 5370 8708 5714
rect 8668 5364 8720 5370
rect 8668 5306 8720 5312
rect 9232 5302 9260 6598
rect 9416 6118 9444 6990
rect 9496 6928 9548 6934
rect 9496 6870 9548 6876
rect 9508 6730 9536 6870
rect 9600 6798 9628 7686
rect 9692 7546 9720 8434
rect 9954 7576 10010 7585
rect 9680 7540 9732 7546
rect 9954 7511 10010 7520
rect 9680 7482 9732 7488
rect 9588 6792 9640 6798
rect 9588 6734 9640 6740
rect 9496 6724 9548 6730
rect 9496 6666 9548 6672
rect 9692 6458 9720 7482
rect 9864 7404 9916 7410
rect 9864 7346 9916 7352
rect 9772 7200 9824 7206
rect 9772 7142 9824 7148
rect 9784 7002 9812 7142
rect 9876 7002 9904 7346
rect 9772 6996 9824 7002
rect 9772 6938 9824 6944
rect 9864 6996 9916 7002
rect 9864 6938 9916 6944
rect 9680 6452 9732 6458
rect 9680 6394 9732 6400
rect 9404 6112 9456 6118
rect 9404 6054 9456 6060
rect 9588 6112 9640 6118
rect 9588 6054 9640 6060
rect 9404 5568 9456 5574
rect 9404 5510 9456 5516
rect 9496 5568 9548 5574
rect 9496 5510 9548 5516
rect 8392 5296 8444 5302
rect 8392 5238 8444 5244
rect 9220 5296 9272 5302
rect 9220 5238 9272 5244
rect 7012 5160 7064 5166
rect 7012 5102 7064 5108
rect 7472 5160 7524 5166
rect 7472 5102 7524 5108
rect 6828 4820 6880 4826
rect 6828 4762 6880 4768
rect 6736 4684 6788 4690
rect 6736 4626 6788 4632
rect 6460 4208 6512 4214
rect 6460 4150 6512 4156
rect 6092 4140 6144 4146
rect 6092 4082 6144 4088
rect 6840 4078 6868 4762
rect 7024 4690 7052 5102
rect 8404 4826 8432 5238
rect 8760 5228 8812 5234
rect 8760 5170 8812 5176
rect 8772 4826 8800 5170
rect 9416 4826 9444 5510
rect 9508 5370 9536 5510
rect 9496 5364 9548 5370
rect 9496 5306 9548 5312
rect 9600 5234 9628 6054
rect 9876 5710 9904 6938
rect 9968 6458 9996 7511
rect 9956 6452 10008 6458
rect 9956 6394 10008 6400
rect 10324 6316 10376 6322
rect 10324 6258 10376 6264
rect 10336 6225 10364 6258
rect 10322 6216 10378 6225
rect 10322 6151 10378 6160
rect 9864 5704 9916 5710
rect 9864 5646 9916 5652
rect 9956 5704 10008 5710
rect 9956 5646 10008 5652
rect 9968 5370 9996 5646
rect 9956 5364 10008 5370
rect 9956 5306 10008 5312
rect 9588 5228 9640 5234
rect 9588 5170 9640 5176
rect 8392 4820 8444 4826
rect 8392 4762 8444 4768
rect 8760 4820 8812 4826
rect 8760 4762 8812 4768
rect 9404 4820 9456 4826
rect 9404 4762 9456 4768
rect 7012 4684 7064 4690
rect 7012 4626 7064 4632
rect 8404 4622 8432 4762
rect 8392 4616 8444 4622
rect 8392 4558 8444 4564
rect 3792 4072 3844 4078
rect 3792 4014 3844 4020
rect 4528 4072 4580 4078
rect 4528 4014 4580 4020
rect 4804 4072 4856 4078
rect 4804 4014 4856 4020
rect 5540 4072 5592 4078
rect 5540 4014 5592 4020
rect 5724 4072 5776 4078
rect 5724 4014 5776 4020
rect 6828 4072 6880 4078
rect 6828 4014 6880 4020
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 5540 3664 5592 3670
rect 5540 3606 5592 3612
rect 8484 3664 8536 3670
rect 8484 3606 8536 3612
rect 1676 3528 1728 3534
rect 1214 3496 1270 3505
rect 1676 3470 1728 3476
rect 4068 3528 4120 3534
rect 4068 3470 4120 3476
rect 1214 3431 1270 3440
rect 1228 3398 1256 3431
rect 1216 3392 1268 3398
rect 1216 3334 1268 3340
rect 1688 3194 1716 3470
rect 1676 3188 1728 3194
rect 1676 3130 1728 3136
rect 3884 3188 3936 3194
rect 3884 3130 3936 3136
rect 1400 3052 1452 3058
rect 1400 2994 1452 3000
rect 2964 3052 3016 3058
rect 2964 2994 3016 3000
rect 1412 2825 1440 2994
rect 2596 2848 2648 2854
rect 1398 2816 1454 2825
rect 2596 2790 2648 2796
rect 1398 2751 1454 2760
rect 2044 2440 2096 2446
rect 2044 2382 2096 2388
rect 2056 1306 2084 2382
rect 1964 1278 2084 1306
rect 1964 800 1992 1278
rect 2608 800 2636 2790
rect 2976 2650 3004 2994
rect 3240 2984 3292 2990
rect 3240 2926 3292 2932
rect 3516 2984 3568 2990
rect 3516 2926 3568 2932
rect 2964 2644 3016 2650
rect 2964 2586 3016 2592
rect 3252 2514 3280 2926
rect 3424 2848 3476 2854
rect 3424 2790 3476 2796
rect 3436 2514 3464 2790
rect 3240 2508 3292 2514
rect 3240 2450 3292 2456
rect 3424 2508 3476 2514
rect 3424 2450 3476 2456
rect 3528 2446 3556 2926
rect 3896 2854 3924 3130
rect 4080 3058 4108 3470
rect 5552 3398 5580 3606
rect 6092 3596 6144 3602
rect 6092 3538 6144 3544
rect 5724 3460 5776 3466
rect 5724 3402 5776 3408
rect 5828 3454 6040 3482
rect 4804 3392 4856 3398
rect 4804 3334 4856 3340
rect 5540 3392 5592 3398
rect 5540 3334 5592 3340
rect 5632 3392 5684 3398
rect 5632 3334 5684 3340
rect 4068 3052 4120 3058
rect 4068 2994 4120 3000
rect 3976 2984 4028 2990
rect 3976 2926 4028 2932
rect 3608 2848 3660 2854
rect 3608 2790 3660 2796
rect 3884 2848 3936 2854
rect 3884 2790 3936 2796
rect 3620 2446 3648 2790
rect 3516 2440 3568 2446
rect 3516 2382 3568 2388
rect 3608 2440 3660 2446
rect 3608 2382 3660 2388
rect 3240 2304 3292 2310
rect 3240 2246 3292 2252
rect 3252 800 3280 2246
rect 3988 1578 4016 2926
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 4816 2446 4844 3334
rect 4874 3292 5182 3301
rect 4874 3290 4880 3292
rect 4936 3290 4960 3292
rect 5016 3290 5040 3292
rect 5096 3290 5120 3292
rect 5176 3290 5182 3292
rect 4936 3238 4938 3290
rect 5118 3238 5120 3290
rect 4874 3236 4880 3238
rect 4936 3236 4960 3238
rect 5016 3236 5040 3238
rect 5096 3236 5120 3238
rect 5176 3236 5182 3238
rect 4874 3227 5182 3236
rect 5552 2854 5580 3334
rect 5644 3058 5672 3334
rect 5736 3194 5764 3402
rect 5724 3188 5776 3194
rect 5724 3130 5776 3136
rect 5632 3052 5684 3058
rect 5632 2994 5684 3000
rect 5540 2848 5592 2854
rect 5540 2790 5592 2796
rect 4620 2440 4672 2446
rect 3896 1550 4016 1578
rect 4540 2400 4620 2428
rect 3896 800 3924 1550
rect 4540 800 4568 2400
rect 4620 2382 4672 2388
rect 4804 2440 4856 2446
rect 4804 2382 4856 2388
rect 4804 2304 4856 2310
rect 4804 2246 4856 2252
rect 1950 0 2006 800
rect 2594 0 2650 800
rect 3238 0 3294 800
rect 3882 0 3938 800
rect 4526 0 4582 800
rect 4816 762 4844 2246
rect 4874 2204 5182 2213
rect 4874 2202 4880 2204
rect 4936 2202 4960 2204
rect 5016 2202 5040 2204
rect 5096 2202 5120 2204
rect 5176 2202 5182 2204
rect 4936 2150 4938 2202
rect 5118 2150 5120 2202
rect 4874 2148 4880 2150
rect 4936 2148 4960 2150
rect 5016 2148 5040 2150
rect 5096 2148 5120 2150
rect 5176 2148 5182 2150
rect 4874 2139 5182 2148
rect 5092 870 5212 898
rect 5092 762 5120 870
rect 5184 800 5212 870
rect 5828 800 5856 3454
rect 6012 3398 6040 3454
rect 6000 3392 6052 3398
rect 6000 3334 6052 3340
rect 6000 3120 6052 3126
rect 5920 3068 6000 3074
rect 6104 3074 6132 3538
rect 7840 3188 7892 3194
rect 7840 3130 7892 3136
rect 6052 3068 6132 3074
rect 5920 3046 6132 3068
rect 5920 2446 5948 3046
rect 6092 2984 6144 2990
rect 6012 2932 6092 2938
rect 6012 2926 6144 2932
rect 6012 2910 6132 2926
rect 6012 2854 6040 2910
rect 6000 2848 6052 2854
rect 6000 2790 6052 2796
rect 6368 2848 6420 2854
rect 6368 2790 6420 2796
rect 6012 2650 6040 2790
rect 6000 2644 6052 2650
rect 6000 2586 6052 2592
rect 6380 2446 6408 2790
rect 7852 2446 7880 3130
rect 8496 2446 8524 3606
rect 5908 2440 5960 2446
rect 5908 2382 5960 2388
rect 6368 2440 6420 2446
rect 6368 2382 6420 2388
rect 7840 2440 7892 2446
rect 7840 2382 7892 2388
rect 8484 2440 8536 2446
rect 8484 2382 8536 2388
rect 6460 2304 6512 2310
rect 6460 2246 6512 2252
rect 7104 2304 7156 2310
rect 7104 2246 7156 2252
rect 7748 2304 7800 2310
rect 7748 2246 7800 2252
rect 8392 2304 8444 2310
rect 8392 2246 8444 2252
rect 6472 800 6500 2246
rect 7116 800 7144 2246
rect 7760 800 7788 2246
rect 8404 800 8432 2246
rect 4816 734 5120 762
rect 5170 0 5226 800
rect 5814 0 5870 800
rect 6458 0 6514 800
rect 7102 0 7158 800
rect 7746 0 7802 800
rect 8390 0 8446 800
<< via2 >>
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 1490 6876 1492 6896
rect 1492 6876 1544 6896
rect 1544 6876 1546 6896
rect 1490 6840 1546 6876
rect 1398 6296 1454 6352
rect 1030 5480 1086 5536
rect 4880 10906 4936 10908
rect 4960 10906 5016 10908
rect 5040 10906 5096 10908
rect 5120 10906 5176 10908
rect 4880 10854 4926 10906
rect 4926 10854 4936 10906
rect 4960 10854 4990 10906
rect 4990 10854 5002 10906
rect 5002 10854 5016 10906
rect 5040 10854 5054 10906
rect 5054 10854 5066 10906
rect 5066 10854 5096 10906
rect 5120 10854 5130 10906
rect 5130 10854 5176 10906
rect 4880 10852 4936 10854
rect 4960 10852 5016 10854
rect 5040 10852 5096 10854
rect 5120 10852 5176 10854
rect 4880 9818 4936 9820
rect 4960 9818 5016 9820
rect 5040 9818 5096 9820
rect 5120 9818 5176 9820
rect 4880 9766 4926 9818
rect 4926 9766 4936 9818
rect 4960 9766 4990 9818
rect 4990 9766 5002 9818
rect 5002 9766 5016 9818
rect 5040 9766 5054 9818
rect 5054 9766 5066 9818
rect 5066 9766 5096 9818
rect 5120 9766 5130 9818
rect 5130 9766 5176 9818
rect 4880 9764 4936 9766
rect 4960 9764 5016 9766
rect 5040 9764 5096 9766
rect 5120 9764 5176 9766
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4710 9560 4766 9616
rect 2042 6724 2098 6760
rect 2042 6704 2044 6724
rect 2044 6704 2096 6724
rect 2096 6704 2098 6724
rect 3606 8472 3662 8528
rect 1490 4800 1546 4856
rect 3514 6160 3570 6216
rect 3146 5752 3202 5808
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4880 8730 4936 8732
rect 4960 8730 5016 8732
rect 5040 8730 5096 8732
rect 5120 8730 5176 8732
rect 4880 8678 4926 8730
rect 4926 8678 4936 8730
rect 4960 8678 4990 8730
rect 4990 8678 5002 8730
rect 5002 8678 5016 8730
rect 5040 8678 5054 8730
rect 5054 8678 5066 8730
rect 5066 8678 5096 8730
rect 5120 8678 5130 8730
rect 5130 8678 5176 8730
rect 4880 8676 4936 8678
rect 4960 8676 5016 8678
rect 5040 8676 5096 8678
rect 5120 8676 5176 8678
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 5354 8472 5410 8528
rect 4880 7642 4936 7644
rect 4960 7642 5016 7644
rect 5040 7642 5096 7644
rect 5120 7642 5176 7644
rect 4880 7590 4926 7642
rect 4926 7590 4936 7642
rect 4960 7590 4990 7642
rect 4990 7590 5002 7642
rect 5002 7590 5016 7642
rect 5040 7590 5054 7642
rect 5054 7590 5066 7642
rect 5066 7590 5096 7642
rect 5120 7590 5130 7642
rect 5130 7590 5176 7642
rect 4880 7588 4936 7590
rect 4960 7588 5016 7590
rect 5040 7588 5096 7590
rect 5120 7588 5176 7590
rect 4342 6296 4398 6352
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4250 5752 4306 5808
rect 1950 4140 2006 4176
rect 1950 4120 1952 4140
rect 1952 4120 2004 4140
rect 2004 4120 2006 4140
rect 4880 6554 4936 6556
rect 4960 6554 5016 6556
rect 5040 6554 5096 6556
rect 5120 6554 5176 6556
rect 4880 6502 4926 6554
rect 4926 6502 4936 6554
rect 4960 6502 4990 6554
rect 4990 6502 5002 6554
rect 5002 6502 5016 6554
rect 5040 6502 5054 6554
rect 5054 6502 5066 6554
rect 5066 6502 5096 6554
rect 5120 6502 5130 6554
rect 5130 6502 5176 6554
rect 4880 6500 4936 6502
rect 4960 6500 5016 6502
rect 5040 6500 5096 6502
rect 5120 6500 5176 6502
rect 6090 8492 6146 8528
rect 6090 8472 6092 8492
rect 6092 8472 6144 8492
rect 6144 8472 6146 8492
rect 5722 6704 5778 6760
rect 5538 6160 5594 6216
rect 4894 6024 4950 6080
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4880 5466 4936 5468
rect 4960 5466 5016 5468
rect 5040 5466 5096 5468
rect 5120 5466 5176 5468
rect 4880 5414 4926 5466
rect 4926 5414 4936 5466
rect 4960 5414 4990 5466
rect 4990 5414 5002 5466
rect 5002 5414 5016 5466
rect 5040 5414 5054 5466
rect 5054 5414 5066 5466
rect 5066 5414 5096 5466
rect 5120 5414 5130 5466
rect 5130 5414 5176 5466
rect 4880 5412 4936 5414
rect 4960 5412 5016 5414
rect 5040 5412 5096 5414
rect 5120 5412 5176 5414
rect 4880 4378 4936 4380
rect 4960 4378 5016 4380
rect 5040 4378 5096 4380
rect 5120 4378 5176 4380
rect 4880 4326 4926 4378
rect 4926 4326 4936 4378
rect 4960 4326 4990 4378
rect 4990 4326 5002 4378
rect 5002 4326 5016 4378
rect 5040 4326 5054 4378
rect 5054 4326 5066 4378
rect 5066 4326 5096 4378
rect 5120 4326 5130 4378
rect 5130 4326 5176 4378
rect 4880 4324 4936 4326
rect 4960 4324 5016 4326
rect 5040 4324 5096 4326
rect 5120 4324 5176 4326
rect 5906 6316 5962 6352
rect 5906 6296 5908 6316
rect 5908 6296 5960 6316
rect 5960 6296 5962 6316
rect 6090 6160 6146 6216
rect 5906 6024 5962 6080
rect 7470 6160 7526 6216
rect 9954 7520 10010 7576
rect 10322 6160 10378 6216
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 1214 3440 1270 3496
rect 1398 2760 1454 2816
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 4880 3290 4936 3292
rect 4960 3290 5016 3292
rect 5040 3290 5096 3292
rect 5120 3290 5176 3292
rect 4880 3238 4926 3290
rect 4926 3238 4936 3290
rect 4960 3238 4990 3290
rect 4990 3238 5002 3290
rect 5002 3238 5016 3290
rect 5040 3238 5054 3290
rect 5054 3238 5066 3290
rect 5066 3238 5096 3290
rect 5120 3238 5130 3290
rect 5130 3238 5176 3290
rect 4880 3236 4936 3238
rect 4960 3236 5016 3238
rect 5040 3236 5096 3238
rect 5120 3236 5176 3238
rect 4880 2202 4936 2204
rect 4960 2202 5016 2204
rect 5040 2202 5096 2204
rect 5120 2202 5176 2204
rect 4880 2150 4926 2202
rect 4926 2150 4936 2202
rect 4960 2150 4990 2202
rect 4990 2150 5002 2202
rect 5002 2150 5016 2202
rect 5040 2150 5054 2202
rect 5054 2150 5066 2202
rect 5066 2150 5096 2202
rect 5120 2150 5130 2202
rect 5130 2150 5176 2202
rect 4880 2148 4936 2150
rect 4960 2148 5016 2150
rect 5040 2148 5096 2150
rect 5120 2148 5176 2150
<< metal3 >>
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 4870 10912 5186 10913
rect 4870 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5186 10912
rect 4870 10847 5186 10848
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 4870 9824 5186 9825
rect 4870 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5186 9824
rect 4870 9759 5186 9760
rect 0 9618 800 9648
rect 4705 9618 4771 9621
rect 0 9616 4771 9618
rect 0 9560 4710 9616
rect 4766 9560 4771 9616
rect 0 9558 4771 9560
rect 0 9528 800 9558
rect 4705 9555 4771 9558
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 4870 8736 5186 8737
rect 4870 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5186 8736
rect 4870 8671 5186 8672
rect 3601 8530 3667 8533
rect 5349 8530 5415 8533
rect 6085 8530 6151 8533
rect 3601 8528 6151 8530
rect 3601 8472 3606 8528
rect 3662 8472 5354 8528
rect 5410 8472 6090 8528
rect 6146 8472 6151 8528
rect 3601 8470 6151 8472
rect 3601 8467 3667 8470
rect 5349 8467 5415 8470
rect 6085 8467 6151 8470
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 4870 7648 5186 7649
rect 4870 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5186 7648
rect 4870 7583 5186 7584
rect 9949 7578 10015 7581
rect 10740 7578 11540 7608
rect 9949 7576 11540 7578
rect 9949 7520 9954 7576
rect 10010 7520 11540 7576
rect 9949 7518 11540 7520
rect 9949 7515 10015 7518
rect 10740 7488 11540 7518
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 0 6898 800 6928
rect 1485 6898 1551 6901
rect 0 6896 1551 6898
rect 0 6840 1490 6896
rect 1546 6840 1551 6896
rect 0 6838 1551 6840
rect 0 6808 800 6838
rect 1485 6835 1551 6838
rect 2037 6762 2103 6765
rect 5717 6762 5783 6765
rect 2037 6760 5783 6762
rect 2037 6704 2042 6760
rect 2098 6704 5722 6760
rect 5778 6704 5783 6760
rect 2037 6702 5783 6704
rect 2037 6699 2103 6702
rect 5717 6699 5783 6702
rect 4870 6560 5186 6561
rect 4870 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5186 6560
rect 4870 6495 5186 6496
rect 1393 6354 1459 6357
rect 982 6352 1459 6354
rect 982 6296 1398 6352
rect 1454 6296 1459 6352
rect 982 6294 1459 6296
rect 0 6218 800 6248
rect 982 6218 1042 6294
rect 1393 6291 1459 6294
rect 4337 6354 4403 6357
rect 5901 6354 5967 6357
rect 4337 6352 5967 6354
rect 4337 6296 4342 6352
rect 4398 6296 5906 6352
rect 5962 6296 5967 6352
rect 4337 6294 5967 6296
rect 4337 6291 4403 6294
rect 5901 6291 5967 6294
rect 0 6158 1042 6218
rect 3509 6218 3575 6221
rect 5533 6218 5599 6221
rect 3509 6216 5599 6218
rect 3509 6160 3514 6216
rect 3570 6160 5538 6216
rect 5594 6160 5599 6216
rect 3509 6158 5599 6160
rect 0 6128 800 6158
rect 3509 6155 3575 6158
rect 5533 6155 5599 6158
rect 6085 6218 6151 6221
rect 7465 6218 7531 6221
rect 6085 6216 7531 6218
rect 6085 6160 6090 6216
rect 6146 6160 7470 6216
rect 7526 6160 7531 6216
rect 6085 6158 7531 6160
rect 6085 6155 6151 6158
rect 7465 6155 7531 6158
rect 10317 6218 10383 6221
rect 10740 6218 11540 6248
rect 10317 6216 11540 6218
rect 10317 6160 10322 6216
rect 10378 6160 11540 6216
rect 10317 6158 11540 6160
rect 10317 6155 10383 6158
rect 10740 6128 11540 6158
rect 4889 6082 4955 6085
rect 5901 6082 5967 6085
rect 4889 6080 5967 6082
rect 4889 6024 4894 6080
rect 4950 6024 5906 6080
rect 5962 6024 5967 6080
rect 4889 6022 5967 6024
rect 4889 6019 4955 6022
rect 5901 6019 5967 6022
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 3141 5810 3207 5813
rect 4245 5810 4311 5813
rect 3141 5808 4311 5810
rect 3141 5752 3146 5808
rect 3202 5752 4250 5808
rect 4306 5752 4311 5808
rect 3141 5750 4311 5752
rect 3141 5747 3207 5750
rect 4245 5747 4311 5750
rect 0 5538 800 5568
rect 1025 5538 1091 5541
rect 0 5536 1091 5538
rect 0 5480 1030 5536
rect 1086 5480 1091 5536
rect 0 5478 1091 5480
rect 0 5448 800 5478
rect 1025 5475 1091 5478
rect 4870 5472 5186 5473
rect 4870 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5186 5472
rect 4870 5407 5186 5408
rect 4210 4928 4526 4929
rect 0 4858 800 4888
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 1485 4858 1551 4861
rect 0 4856 1551 4858
rect 0 4800 1490 4856
rect 1546 4800 1551 4856
rect 0 4798 1551 4800
rect 0 4768 800 4798
rect 1485 4795 1551 4798
rect 4870 4384 5186 4385
rect 4870 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5186 4384
rect 4870 4319 5186 4320
rect 0 4178 800 4208
rect 1945 4178 2011 4181
rect 0 4176 2011 4178
rect 0 4120 1950 4176
rect 2006 4120 2011 4176
rect 0 4118 2011 4120
rect 0 4088 800 4118
rect 1945 4115 2011 4118
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 798 3574 1226 3634
rect 798 3528 858 3574
rect 0 3438 858 3528
rect 1166 3501 1226 3574
rect 1166 3496 1275 3501
rect 1166 3440 1214 3496
rect 1270 3440 1275 3496
rect 1166 3438 1275 3440
rect 0 3408 800 3438
rect 1209 3435 1275 3438
rect 4870 3296 5186 3297
rect 4870 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5186 3296
rect 4870 3231 5186 3232
rect 0 2818 800 2848
rect 1393 2818 1459 2821
rect 0 2816 1459 2818
rect 0 2760 1398 2816
rect 1454 2760 1459 2816
rect 0 2758 1459 2760
rect 0 2728 800 2758
rect 1393 2755 1459 2758
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 4870 2208 5186 2209
rect 4870 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5186 2208
rect 4870 2143 5186 2144
<< via3 >>
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 4876 10908 4940 10912
rect 4876 10852 4880 10908
rect 4880 10852 4936 10908
rect 4936 10852 4940 10908
rect 4876 10848 4940 10852
rect 4956 10908 5020 10912
rect 4956 10852 4960 10908
rect 4960 10852 5016 10908
rect 5016 10852 5020 10908
rect 4956 10848 5020 10852
rect 5036 10908 5100 10912
rect 5036 10852 5040 10908
rect 5040 10852 5096 10908
rect 5096 10852 5100 10908
rect 5036 10848 5100 10852
rect 5116 10908 5180 10912
rect 5116 10852 5120 10908
rect 5120 10852 5176 10908
rect 5176 10852 5180 10908
rect 5116 10848 5180 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 4876 9820 4940 9824
rect 4876 9764 4880 9820
rect 4880 9764 4936 9820
rect 4936 9764 4940 9820
rect 4876 9760 4940 9764
rect 4956 9820 5020 9824
rect 4956 9764 4960 9820
rect 4960 9764 5016 9820
rect 5016 9764 5020 9820
rect 4956 9760 5020 9764
rect 5036 9820 5100 9824
rect 5036 9764 5040 9820
rect 5040 9764 5096 9820
rect 5096 9764 5100 9820
rect 5036 9760 5100 9764
rect 5116 9820 5180 9824
rect 5116 9764 5120 9820
rect 5120 9764 5176 9820
rect 5176 9764 5180 9820
rect 5116 9760 5180 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 4876 8732 4940 8736
rect 4876 8676 4880 8732
rect 4880 8676 4936 8732
rect 4936 8676 4940 8732
rect 4876 8672 4940 8676
rect 4956 8732 5020 8736
rect 4956 8676 4960 8732
rect 4960 8676 5016 8732
rect 5016 8676 5020 8732
rect 4956 8672 5020 8676
rect 5036 8732 5100 8736
rect 5036 8676 5040 8732
rect 5040 8676 5096 8732
rect 5096 8676 5100 8732
rect 5036 8672 5100 8676
rect 5116 8732 5180 8736
rect 5116 8676 5120 8732
rect 5120 8676 5176 8732
rect 5176 8676 5180 8732
rect 5116 8672 5180 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 4876 7644 4940 7648
rect 4876 7588 4880 7644
rect 4880 7588 4936 7644
rect 4936 7588 4940 7644
rect 4876 7584 4940 7588
rect 4956 7644 5020 7648
rect 4956 7588 4960 7644
rect 4960 7588 5016 7644
rect 5016 7588 5020 7644
rect 4956 7584 5020 7588
rect 5036 7644 5100 7648
rect 5036 7588 5040 7644
rect 5040 7588 5096 7644
rect 5096 7588 5100 7644
rect 5036 7584 5100 7588
rect 5116 7644 5180 7648
rect 5116 7588 5120 7644
rect 5120 7588 5176 7644
rect 5176 7588 5180 7644
rect 5116 7584 5180 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 4876 6556 4940 6560
rect 4876 6500 4880 6556
rect 4880 6500 4936 6556
rect 4936 6500 4940 6556
rect 4876 6496 4940 6500
rect 4956 6556 5020 6560
rect 4956 6500 4960 6556
rect 4960 6500 5016 6556
rect 5016 6500 5020 6556
rect 4956 6496 5020 6500
rect 5036 6556 5100 6560
rect 5036 6500 5040 6556
rect 5040 6500 5096 6556
rect 5096 6500 5100 6556
rect 5036 6496 5100 6500
rect 5116 6556 5180 6560
rect 5116 6500 5120 6556
rect 5120 6500 5176 6556
rect 5176 6500 5180 6556
rect 5116 6496 5180 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 4876 5468 4940 5472
rect 4876 5412 4880 5468
rect 4880 5412 4936 5468
rect 4936 5412 4940 5468
rect 4876 5408 4940 5412
rect 4956 5468 5020 5472
rect 4956 5412 4960 5468
rect 4960 5412 5016 5468
rect 5016 5412 5020 5468
rect 4956 5408 5020 5412
rect 5036 5468 5100 5472
rect 5036 5412 5040 5468
rect 5040 5412 5096 5468
rect 5096 5412 5100 5468
rect 5036 5408 5100 5412
rect 5116 5468 5180 5472
rect 5116 5412 5120 5468
rect 5120 5412 5176 5468
rect 5176 5412 5180 5468
rect 5116 5408 5180 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 4876 4380 4940 4384
rect 4876 4324 4880 4380
rect 4880 4324 4936 4380
rect 4936 4324 4940 4380
rect 4876 4320 4940 4324
rect 4956 4380 5020 4384
rect 4956 4324 4960 4380
rect 4960 4324 5016 4380
rect 5016 4324 5020 4380
rect 4956 4320 5020 4324
rect 5036 4380 5100 4384
rect 5036 4324 5040 4380
rect 5040 4324 5096 4380
rect 5096 4324 5100 4380
rect 5036 4320 5100 4324
rect 5116 4380 5180 4384
rect 5116 4324 5120 4380
rect 5120 4324 5176 4380
rect 5176 4324 5180 4380
rect 5116 4320 5180 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 4876 3292 4940 3296
rect 4876 3236 4880 3292
rect 4880 3236 4936 3292
rect 4936 3236 4940 3292
rect 4876 3232 4940 3236
rect 4956 3292 5020 3296
rect 4956 3236 4960 3292
rect 4960 3236 5016 3292
rect 5016 3236 5020 3292
rect 4956 3232 5020 3236
rect 5036 3292 5100 3296
rect 5036 3236 5040 3292
rect 5040 3236 5096 3292
rect 5096 3236 5100 3292
rect 5036 3232 5100 3236
rect 5116 3292 5180 3296
rect 5116 3236 5120 3292
rect 5120 3236 5176 3292
rect 5176 3236 5180 3292
rect 5116 3232 5180 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 4876 2204 4940 2208
rect 4876 2148 4880 2204
rect 4880 2148 4936 2204
rect 4936 2148 4940 2204
rect 4876 2144 4940 2148
rect 4956 2204 5020 2208
rect 4956 2148 4960 2204
rect 4960 2148 5016 2204
rect 5016 2148 5020 2204
rect 4956 2144 5020 2148
rect 5036 2204 5100 2208
rect 5036 2148 5040 2204
rect 5040 2148 5096 2204
rect 5096 2148 5100 2204
rect 5036 2144 5100 2148
rect 5116 2204 5180 2208
rect 5116 2148 5120 2204
rect 5120 2148 5176 2204
rect 5176 2148 5180 2204
rect 5116 2144 5180 2148
<< metal4 >>
rect 4208 11456 4528 11472
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 4868 10912 5188 11472
rect 4868 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5188 10912
rect 4868 9824 5188 10848
rect 4868 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5188 9824
rect 4868 8736 5188 9760
rect 4868 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5188 8736
rect 4868 7648 5188 8672
rect 4868 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5188 7648
rect 4868 6560 5188 7584
rect 4868 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5188 6560
rect 4868 5472 5188 6496
rect 4868 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5188 5472
rect 4868 4384 5188 5408
rect 4868 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5188 4384
rect 4868 3296 5188 4320
rect 4868 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5188 3296
rect 4868 2208 5188 3232
rect 4868 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5188 2208
rect 4868 2128 5188 2144
use sky130_fd_sc_hd__inv_2  _054_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712980491
transform 1 0 1748 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _055_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712980491
transform -1 0 9476 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _056_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712980491
transform 1 0 8372 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _057_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712980491
transform -1 0 9568 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _058_
timestamp 1712980491
transform 1 0 7084 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _059_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712980491
transform 1 0 8924 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _060_
timestamp 1712980491
transform 1 0 4692 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__nand4_2  _061_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712980491
transform 1 0 4600 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__nand4_1  _062_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712980491
transform 1 0 4508 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _063_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712980491
transform 1 0 6900 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _064_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712980491
transform 1 0 3404 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_1  _065_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712980491
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_1  _066_
timestamp 1712980491
transform -1 0 5980 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__nor3b_1  _067_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712980491
transform 1 0 3128 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__nor3b_1  _068_
timestamp 1712980491
transform -1 0 3680 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _069_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712980491
transform 1 0 5612 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__nor3b_1  _070_
timestamp 1712980491
transform 1 0 4784 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _071_
timestamp 1712980491
transform -1 0 6992 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _072_
timestamp 1712980491
transform 1 0 4968 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _073_
timestamp 1712980491
transform 1 0 5796 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _074_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712980491
transform -1 0 2208 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_1  _075_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712980491
transform -1 0 2024 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__o311a_1  _076_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712980491
transform 1 0 6348 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _077_
timestamp 1712980491
transform -1 0 9752 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _078_
timestamp 1712980491
transform -1 0 9200 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _079_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712980491
transform -1 0 10120 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _080_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712980491
transform 1 0 8924 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _081_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712980491
transform 1 0 9568 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _082_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712980491
transform -1 0 9936 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _083_
timestamp 1712980491
transform 1 0 8556 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _084_
timestamp 1712980491
transform 1 0 9476 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _085_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712980491
transform 1 0 9476 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _086_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712980491
transform -1 0 9476 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _087_
timestamp 1712980491
transform -1 0 8188 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _088_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712980491
transform -1 0 8096 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__nand2b_1  _089_
timestamp 1712980491
transform 1 0 5060 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _090_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712980491
transform -1 0 6256 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _091_
timestamp 1712980491
transform 1 0 3588 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _092_
timestamp 1712980491
transform 1 0 5888 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _093_
timestamp 1712980491
transform -1 0 6164 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _094_
timestamp 1712980491
transform 1 0 5612 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _095_
timestamp 1712980491
transform 1 0 6348 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__nand4_1  _096_
timestamp 1712980491
transform -1 0 4692 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _097_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712980491
transform 1 0 4600 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _098_
timestamp 1712980491
transform 1 0 2576 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a41o_1  _099_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712980491
transform 1 0 3864 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _100_
timestamp 1712980491
transform -1 0 4416 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _101_
timestamp 1712980491
transform 1 0 3128 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _102_
timestamp 1712980491
transform -1 0 6072 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _103_
timestamp 1712980491
transform 1 0 6348 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _104_
timestamp 1712980491
transform -1 0 5888 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _105_
timestamp 1712980491
transform -1 0 6532 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _106_
timestamp 1712980491
transform 1 0 3312 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _107_
timestamp 1712980491
transform 1 0 4324 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _108_
timestamp 1712980491
transform 1 0 3772 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _109_
timestamp 1712980491
transform -1 0 4600 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _110_
timestamp 1712980491
transform 1 0 4600 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _111_
timestamp 1712980491
transform 1 0 5060 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _112_
timestamp 1712980491
transform 1 0 3772 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__nand4_1  _113_
timestamp 1712980491
transform 1 0 3220 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _114_
timestamp 1712980491
transform 1 0 2760 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _115_
timestamp 1712980491
transform -1 0 3680 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _116_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712980491
transform 1 0 3772 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _117_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712980491
transform -1 0 5060 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__o2111a_1  _118_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712980491
transform 1 0 4968 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_1  _119_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712980491
transform 1 0 3864 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _120_
timestamp 1712980491
transform 1 0 4508 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__dfrtp_1  _121_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712980491
transform 1 0 7084 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _122_
timestamp 1712980491
transform 1 0 6900 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _123_
timestamp 1712980491
transform 1 0 6900 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _124_
timestamp 1712980491
transform 1 0 6992 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _125_
timestamp 1712980491
transform 1 0 6716 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _126_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712980491
transform 1 0 5520 0 1 9792
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _127_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712980491
transform 1 0 6348 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _128_
timestamp 1712980491
transform 1 0 2760 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _129_
timestamp 1712980491
transform 1 0 2760 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _130_
timestamp 1712980491
transform -1 0 6900 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _131_
timestamp 1712980491
transform 1 0 2484 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _132_
timestamp 1712980491
transform -1 0 3220 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _133_
timestamp 1712980491
transform 1 0 1748 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _134_
timestamp 1712980491
transform 1 0 2208 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _135_
timestamp 1712980491
transform 1 0 4232 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _136_
timestamp 1712980491
transform 1 0 5244 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__conb_1  _137__26 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712980491
transform -1 0 2024 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _137_
timestamp 1712980491
transform -1 0 3220 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _138_
timestamp 1712980491
transform 1 0 1380 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_osc_ck $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712980491
transform 1 0 4324 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_osc_ck
timestamp 1712980491
transform -1 0 5888 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_osc_ck
timestamp 1712980491
transform 1 0 5520 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_2  fanout22 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712980491
transform -1 0 6716 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout23
timestamp 1712980491
transform -1 0 6900 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout24 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712980491
transform -1 0 5612 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout25
timestamp 1712980491
transform 1 0 6348 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712980491
transform 1 0 1380 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_9 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712980491
transform 1 0 1932 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_20 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712980491
transform 1 0 2944 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_33
timestamp 1712980491
transform 1 0 4140 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_48 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712980491
transform 1 0 5520 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_57
timestamp 1712980491
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_63
timestamp 1712980491
transform 1 0 6900 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_70
timestamp 1712980491
transform 1 0 7544 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_77
timestamp 1712980491
transform 1 0 8188 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_85 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712980491
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_97
timestamp 1712980491
transform 1 0 10028 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_6
timestamp 1712980491
transform 1 0 1656 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_10
timestamp 1712980491
transform 1 0 2024 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_16
timestamp 1712980491
transform 1 0 2576 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_21
timestamp 1712980491
transform 1 0 3036 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_28
timestamp 1712980491
transform 1 0 3680 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_41
timestamp 1712980491
transform 1 0 4876 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_64
timestamp 1712980491
transform 1 0 6992 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_76
timestamp 1712980491
transform 1 0 8096 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_88 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712980491
transform 1 0 9200 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_96
timestamp 1712980491
transform 1 0 9936 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_7
timestamp 1712980491
transform 1 0 1748 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_19
timestamp 1712980491
transform 1 0 2852 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1712980491
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_29
timestamp 1712980491
transform 1 0 3772 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_37
timestamp 1712980491
transform 1 0 4508 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_46
timestamp 1712980491
transform 1 0 5336 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_57
timestamp 1712980491
transform 1 0 6348 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_69
timestamp 1712980491
transform 1 0 7452 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_81
timestamp 1712980491
transform 1 0 8556 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_85
timestamp 1712980491
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_97
timestamp 1712980491
transform 1 0 10028 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_10
timestamp 1712980491
transform 1 0 2024 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_22
timestamp 1712980491
transform 1 0 3128 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_52 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712980491
transform 1 0 5888 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_61
timestamp 1712980491
transform 1 0 6716 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_73
timestamp 1712980491
transform 1 0 7820 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_85
timestamp 1712980491
transform 1 0 8924 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_97
timestamp 1712980491
transform 1 0 10028 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_3
timestamp 1712980491
transform 1 0 1380 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_13
timestamp 1712980491
transform 1 0 2300 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_25
timestamp 1712980491
transform 1 0 3404 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_29
timestamp 1712980491
transform 1 0 3772 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_33
timestamp 1712980491
transform 1 0 4140 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_62
timestamp 1712980491
transform 1 0 6808 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_85
timestamp 1712980491
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_97
timestamp 1712980491
transform 1 0 10028 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_3
timestamp 1712980491
transform 1 0 1380 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_52
timestamp 1712980491
transform 1 0 5888 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_57
timestamp 1712980491
transform 1 0 6348 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_84
timestamp 1712980491
transform 1 0 8832 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_90
timestamp 1712980491
transform 1 0 9384 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_96
timestamp 1712980491
transform 1 0 9936 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_23
timestamp 1712980491
transform 1 0 3220 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_97
timestamp 1712980491
transform 1 0 10028 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_23
timestamp 1712980491
transform 1 0 3220 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 1712980491
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_65
timestamp 1712980491
transform 1 0 7084 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_77
timestamp 1712980491
transform 1 0 8188 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1712980491
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_66
timestamp 1712980491
transform 1 0 7176 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_78
timestamp 1712980491
transform 1 0 8280 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_96
timestamp 1712980491
transform 1 0 9936 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_3
timestamp 1712980491
transform 1 0 1380 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_13
timestamp 1712980491
transform 1 0 2300 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp 1712980491
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_61
timestamp 1712980491
transform 1 0 6716 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_83
timestamp 1712980491
transform 1 0 8740 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_96
timestamp 1712980491
transform 1 0 9936 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_42
timestamp 1712980491
transform 1 0 4968 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_83
timestamp 1712980491
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_6
timestamp 1712980491
transform 1 0 1656 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_10
timestamp 1712980491
transform 1 0 2024 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_32
timestamp 1712980491
transform 1 0 4048 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_47
timestamp 1712980491
transform 1 0 5428 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_55
timestamp 1712980491
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_61
timestamp 1712980491
transform 1 0 6716 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_94
timestamp 1712980491
transform 1 0 9752 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_3
timestamp 1712980491
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_15
timestamp 1712980491
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 1712980491
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_29
timestamp 1712980491
transform 1 0 3772 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_33
timestamp 1712980491
transform 1 0 4140 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_39
timestamp 1712980491
transform 1 0 4692 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_68
timestamp 1712980491
transform 1 0 7360 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_80
timestamp 1712980491
transform 1 0 8464 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_93
timestamp 1712980491
transform 1 0 9660 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_97
timestamp 1712980491
transform 1 0 10028 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp 1712980491
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_15
timestamp 1712980491
transform 1 0 2484 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_38
timestamp 1712980491
transform 1 0 4600 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_46
timestamp 1712980491
transform 1 0 5336 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_78
timestamp 1712980491
transform 1 0 8280 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_90
timestamp 1712980491
transform 1 0 9384 0 -1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_3
timestamp 1712980491
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_15
timestamp 1712980491
transform 1 0 2484 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_29
timestamp 1712980491
transform 1 0 3772 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_71
timestamp 1712980491
transform 1 0 7636 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_83
timestamp 1712980491
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_85
timestamp 1712980491
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_97
timestamp 1712980491
transform 1 0 10028 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_3
timestamp 1712980491
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_15
timestamp 1712980491
transform 1 0 2484 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_45
timestamp 1712980491
transform 1 0 5244 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_54
timestamp 1712980491
transform 1 0 6072 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_61
timestamp 1712980491
transform 1 0 6716 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_73
timestamp 1712980491
transform 1 0 7820 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_85
timestamp 1712980491
transform 1 0 8924 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_97
timestamp 1712980491
transform 1 0 10028 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_3
timestamp 1712980491
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_15
timestamp 1712980491
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_27
timestamp 1712980491
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_29
timestamp 1712980491
transform 1 0 3772 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_36
timestamp 1712980491
transform 1 0 4416 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_48
timestamp 1712980491
transform 1 0 5520 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_55
timestamp 1712980491
transform 1 0 6164 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_61
timestamp 1712980491
transform 1 0 6716 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_73
timestamp 1712980491
transform 1 0 7820 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_81
timestamp 1712980491
transform 1 0 8556 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_85
timestamp 1712980491
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_97
timestamp 1712980491
transform 1 0 10028 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712980491
transform 1 0 4508 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1712980491
transform 1 0 1564 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1712980491
transform -1 0 6808 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1712980491
transform -1 0 5888 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1712980491
transform -1 0 9660 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1712980491
transform 1 0 3772 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1712980491
transform 1 0 8924 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 1712980491
transform -1 0 8832 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712980491
transform -1 0 1656 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1712980491
transform 1 0 1748 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1712980491
transform -1 0 1656 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input4 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712980491
transform -1 0 9752 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input5 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712980491
transform 1 0 2024 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input6
timestamp 1712980491
transform 1 0 3956 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input7
timestamp 1712980491
transform 1 0 4600 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input8 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712980491
transform 1 0 2024 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output9
timestamp 1712980491
transform -1 0 1748 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output10
timestamp 1712980491
transform -1 0 1748 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output11
timestamp 1712980491
transform 1 0 8464 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output12
timestamp 1712980491
transform -1 0 3036 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output13
timestamp 1712980491
transform 1 0 3772 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output14
timestamp 1712980491
transform 1 0 7820 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output15
timestamp 1712980491
transform -1 0 4600 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output16
timestamp 1712980491
transform 1 0 6532 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output17
timestamp 1712980491
transform 1 0 5980 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output18
timestamp 1712980491
transform 1 0 7176 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output19
timestamp 1712980491
transform -1 0 1748 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output20
timestamp 1712980491
transform -1 0 6716 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output21
timestamp 1712980491
transform 1 0 9752 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_17
timestamp 1712980491
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1712980491
transform -1 0 10396 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_18
timestamp 1712980491
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1712980491
transform -1 0 10396 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_19
timestamp 1712980491
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1712980491
transform -1 0 10396 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_20
timestamp 1712980491
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1712980491
transform -1 0 10396 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_21
timestamp 1712980491
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1712980491
transform -1 0 10396 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_22
timestamp 1712980491
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1712980491
transform -1 0 10396 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_23
timestamp 1712980491
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1712980491
transform -1 0 10396 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_24
timestamp 1712980491
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1712980491
transform -1 0 10396 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_25
timestamp 1712980491
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1712980491
transform -1 0 10396 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_26
timestamp 1712980491
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1712980491
transform -1 0 10396 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_27
timestamp 1712980491
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 1712980491
transform -1 0 10396 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_28
timestamp 1712980491
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 1712980491
transform -1 0 10396 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_29
timestamp 1712980491
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 1712980491
transform -1 0 10396 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_30
timestamp 1712980491
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 1712980491
transform -1 0 10396 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_31
timestamp 1712980491
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 1712980491
transform -1 0 10396 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_32
timestamp 1712980491
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 1712980491
transform -1 0 10396 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_33
timestamp 1712980491
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 1712980491
transform -1 0 10396 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_34 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712980491
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_35
timestamp 1712980491
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_36
timestamp 1712980491
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_37
timestamp 1712980491
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_38
timestamp 1712980491
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_39
timestamp 1712980491
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_40
timestamp 1712980491
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_41
timestamp 1712980491
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_42
timestamp 1712980491
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_43
timestamp 1712980491
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_44
timestamp 1712980491
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_45
timestamp 1712980491
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_46
timestamp 1712980491
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_47
timestamp 1712980491
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_48
timestamp 1712980491
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_49
timestamp 1712980491
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_50
timestamp 1712980491
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_51
timestamp 1712980491
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_52
timestamp 1712980491
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_53
timestamp 1712980491
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_54
timestamp 1712980491
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_55
timestamp 1712980491
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_56
timestamp 1712980491
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_57
timestamp 1712980491
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_58
timestamp 1712980491
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_59
timestamp 1712980491
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_60
timestamp 1712980491
transform 1 0 6256 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_61
timestamp 1712980491
transform 1 0 8832 0 1 10880
box -38 -48 130 592
<< labels >>
flabel metal4 s 4868 2128 5188 11472 0 FreeSans 1920 90 0 0 VGND
port 3 nsew ground bidirectional
flabel metal4 s 4208 2128 4528 11472 0 FreeSans 1920 90 0 0 VPWR
port 2 nsew power bidirectional
flabel metal3 s 0 6128 800 6248 0 FreeSans 480 0 0 0 force_dis_rc_osc
port 17 nsew signal input
flabel metal3 s 0 4088 800 4208 0 FreeSans 480 0 0 0 force_ena_rc_osc
port 18 nsew signal input
flabel metal3 s 0 2728 800 2848 0 FreeSans 480 0 0 0 force_pdn
port 21 nsew signal input
flabel metal3 s 0 3408 800 3528 0 FreeSans 480 0 0 0 force_pdnb
port 4 nsew signal output
flabel metal3 s 10740 6128 11540 6248 0 FreeSans 480 0 0 0 force_short_oneshot
port 23 nsew signal input
flabel metal3 s 0 9528 800 9648 0 FreeSans 480 0 0 0 osc_ck
port 24 nsew signal input
flabel metal3 s 0 4768 800 4888 0 FreeSans 480 0 0 0 osc_ena
port 5 nsew signal output
flabel metal2 s 1950 0 2006 800 0 FreeSans 224 90 0 0 otrip[0]
port 8 nsew signal input
flabel metal2 s 3882 0 3938 800 0 FreeSans 224 90 0 0 otrip[1]
port 7 nsew signal input
flabel metal2 s 4526 0 4582 800 0 FreeSans 224 90 0 0 otrip[2]
port 6 nsew signal input
flabel metal2 s 8390 0 8446 800 0 FreeSans 224 90 0 0 otrip_decoded[0]
port 16 nsew signal output
flabel metal2 s 2594 0 2650 800 0 FreeSans 224 90 0 0 otrip_decoded[1]
port 15 nsew signal output
flabel metal2 s 3238 0 3294 800 0 FreeSans 224 90 0 0 otrip_decoded[2]
port 14 nsew signal output
flabel metal2 s 7746 0 7802 800 0 FreeSans 224 90 0 0 otrip_decoded[3]
port 13 nsew signal output
flabel metal2 s 5170 0 5226 800 0 FreeSans 224 90 0 0 otrip_decoded[4]
port 12 nsew signal output
flabel metal2 s 6458 0 6514 800 0 FreeSans 224 90 0 0 otrip_decoded[5]
port 11 nsew signal output
flabel metal2 s 5814 0 5870 800 0 FreeSans 224 90 0 0 otrip_decoded[6]
port 10 nsew signal output
flabel metal2 s 7102 0 7158 800 0 FreeSans 224 90 0 0 otrip_decoded[7]
port 9 nsew signal output
flabel metal3 s 0 6808 800 6928 0 FreeSans 480 0 0 0 por_timed_out
port 20 nsew signal output
flabel metal2 s 5814 12884 5870 13684 0 FreeSans 224 90 0 0 por_unbuf
port 1 nsew signal output
flabel metal3 s 0 5448 800 5568 0 FreeSans 480 0 0 0 pwup_filt
port 22 nsew signal input
flabel metal3 s 10740 7488 11540 7608 0 FreeSans 480 0 0 0 startup_timed_out
port 19 nsew signal output
rlabel metal1 5750 10880 5750 10880 0 VGND
rlabel metal1 5750 11424 5750 11424 0 VPWR
rlabel metal1 8234 8398 8234 8398 0 _000_
rlabel metal1 8096 7514 8096 7514 0 _001_
rlabel metal1 9108 7242 9108 7242 0 _002_
rlabel metal1 8372 4658 8372 4658 0 _003_
rlabel metal1 7222 5270 7222 5270 0 _004_
rlabel metal1 6026 9690 6026 9690 0 _005_
rlabel metal1 6624 9622 6624 9622 0 _006_
rlabel metal2 3082 10404 3082 10404 0 _007_
rlabel metal1 3128 9622 3128 9622 0 _008_
rlabel metal1 6072 7922 6072 7922 0 _009_
rlabel metal1 2806 7480 2806 7480 0 _010_
rlabel metal1 4094 7786 4094 7786 0 _011_
rlabel via1 2806 6987 2806 6987 0 _012_
rlabel metal2 4738 5882 4738 5882 0 _013_
rlabel metal1 4508 4046 4508 4046 0 _014_
rlabel metal1 5336 4046 5336 4046 0 _015_
rlabel metal1 3634 10064 3634 10064 0 _016_
rlabel metal2 5658 7548 5658 7548 0 _017_
rlabel metal1 6072 7242 6072 7242 0 _018_
rlabel metal1 3956 6766 3956 6766 0 _019_
rlabel metal2 4186 7905 4186 7905 0 _020_
rlabel metal1 4324 7854 4324 7854 0 _021_
rlabel metal1 5106 8432 5106 8432 0 _022_
rlabel metal1 5198 8500 5198 8500 0 _023_
rlabel metal1 3634 6834 3634 6834 0 _024_
rlabel metal2 3266 8262 3266 8262 0 _025_
rlabel metal2 3450 6256 3450 6256 0 _026_
rlabel metal1 3910 4046 3910 4046 0 _027_
rlabel metal2 4830 4794 4830 4794 0 _028_
rlabel metal1 9292 7378 9292 7378 0 _029_
rlabel metal1 8648 6630 8648 6630 0 _030_
rlabel metal1 9062 6290 9062 6290 0 _031_
rlabel metal1 7590 6290 7590 6290 0 _032_
rlabel metal2 5290 10336 5290 10336 0 _033_
rlabel metal1 6164 6290 6164 6290 0 _034_
rlabel metal2 5934 6103 5934 6103 0 _035_
rlabel metal1 6348 6086 6348 6086 0 _036_
rlabel metal1 6762 6324 6762 6324 0 _037_
rlabel metal1 1717 4590 1717 4590 0 _038_
rlabel metal1 9338 8602 9338 8602 0 _039_
rlabel metal1 9108 7378 9108 7378 0 _040_
rlabel metal1 9706 6970 9706 6970 0 _041_
rlabel metal1 9154 5338 9154 5338 0 _042_
rlabel metal1 9936 5338 9936 5338 0 _043_
rlabel metal1 9384 5678 9384 5678 0 _044_
rlabel metal1 8096 5746 8096 5746 0 _045_
rlabel metal1 5520 9146 5520 9146 0 _046_
rlabel metal1 3358 9996 3358 9996 0 _047_
rlabel metal1 6394 8602 6394 8602 0 _048_
rlabel metal1 6256 10642 6256 10642 0 _049_
rlabel metal1 6256 10438 6256 10438 0 _050_
rlabel metal1 3680 9146 3680 9146 0 _051_
rlabel metal1 3082 10064 3082 10064 0 _052_
rlabel metal1 3726 9894 3726 9894 0 _053_
rlabel metal2 5842 6222 5842 6222 0 clknet_0_osc_ck
rlabel metal1 6900 5134 6900 5134 0 clknet_1_0__leaf_osc_ck
rlabel metal2 2806 10064 2806 10064 0 clknet_1_1__leaf_osc_ck
rlabel metal1 5152 9554 5152 9554 0 cnt_por\[0\]
rlabel metal1 6302 5746 6302 5746 0 cnt_por\[10\]
rlabel metal1 5474 9962 5474 9962 0 cnt_por\[1\]
rlabel metal1 4600 8806 4600 8806 0 cnt_por\[2\]
rlabel metal1 4830 9996 4830 9996 0 cnt_por\[3\]
rlabel metal1 4738 7956 4738 7956 0 cnt_por\[4\]
rlabel metal1 5014 6290 5014 6290 0 cnt_por\[5\]
rlabel metal1 2438 7718 2438 7718 0 cnt_por\[6\]
rlabel metal1 3588 6970 3588 6970 0 cnt_por\[7\]
rlabel metal1 3910 6324 3910 6324 0 cnt_por\[8\]
rlabel viali 5290 6293 5290 6293 0 cnt_por\[9\]
rlabel metal1 4554 5644 4554 5644 0 cnt_rsb
rlabel metal1 1518 5882 1518 5882 0 cnt_rsb_stg1
rlabel metal1 9890 6698 9890 6698 0 cnt_st\[0\]
rlabel metal1 9108 6902 9108 6902 0 cnt_st\[1\]
rlabel metal1 8832 7174 8832 7174 0 cnt_st\[2\]
rlabel metal1 9476 5270 9476 5270 0 cnt_st\[3\]
rlabel metal1 7360 6222 7360 6222 0 cnt_st\[4\]
rlabel metal3 843 6188 843 6188 0 force_dis_rc_osc
rlabel metal3 1326 4148 1326 4148 0 force_ena_rc_osc
rlabel metal3 1050 2788 1050 2788 0 force_pdn
rlabel metal3 751 3468 751 3468 0 force_pdnb
rlabel metal1 9706 6256 9706 6256 0 force_short_oneshot
rlabel metal1 1748 5202 1748 5202 0 net1
rlabel metal1 1656 4114 1656 4114 0 net10
rlabel metal1 7222 3638 7222 3638 0 net11
rlabel metal1 3082 2618 3082 2618 0 net12
rlabel metal1 3726 2414 3726 2414 0 net13
rlabel metal1 7038 3162 7038 3162 0 net14
rlabel metal1 4554 2448 4554 2448 0 net15
rlabel metal1 6486 2414 6486 2414 0 net16
rlabel metal1 5658 3162 5658 3162 0 net17
rlabel metal1 6210 2312 6210 2312 0 net18
rlabel metal1 1702 6732 1702 6732 0 net19
rlabel metal1 1886 4250 1886 4250 0 net2
rlabel metal1 6716 6698 6716 6698 0 net20
rlabel metal1 9430 7446 9430 7446 0 net21
rlabel metal1 5934 8398 5934 8398 0 net22
rlabel metal1 5344 10778 5344 10778 0 net23
rlabel metal2 3082 5984 3082 5984 0 net24
rlabel metal1 8379 7854 8379 7854 0 net25
rlabel metal1 2369 8398 2369 8398 0 net26
rlabel metal1 5842 5542 5842 5542 0 net27
rlabel metal1 1978 6222 1978 6222 0 net28
rlabel metal1 5428 4114 5428 4114 0 net29
rlabel metal1 1702 3026 1702 3026 0 net3
rlabel metal1 4094 4046 4094 4046 0 net30
rlabel metal1 8970 8534 8970 8534 0 net31
rlabel metal2 4462 6596 4462 6596 0 net32
rlabel metal2 9614 7242 9614 7242 0 net33
rlabel metal1 8556 5610 8556 5610 0 net34
rlabel via2 6118 8483 6118 8483 0 net4
rlabel metal1 5988 2346 5988 2346 0 net5
rlabel metal1 3312 2482 3312 2482 0 net6
rlabel metal1 4922 2516 4922 2516 0 net7
rlabel metal2 2162 5984 2162 5984 0 net8
rlabel metal1 1794 3162 1794 3162 0 net9
rlabel metal2 4738 8517 4738 8517 0 osc_ck
rlabel metal2 1518 4539 1518 4539 0 osc_ena
rlabel metal2 1978 1027 1978 1027 0 otrip[0]
rlabel metal2 3910 1163 3910 1163 0 otrip[1]
rlabel metal2 4554 1588 4554 1588 0 otrip[2]
rlabel metal2 8418 1520 8418 1520 0 otrip_decoded[0]
rlabel metal2 2622 1792 2622 1792 0 otrip_decoded[1]
rlabel metal2 3266 1520 3266 1520 0 otrip_decoded[2]
rlabel metal2 7774 1520 7774 1520 0 otrip_decoded[3]
rlabel metal2 5198 823 5198 823 0 otrip_decoded[4]
rlabel metal2 6486 1520 6486 1520 0 otrip_decoded[5]
rlabel metal2 5934 3468 5934 3468 0 otrip_decoded[6]
rlabel metal2 7130 1520 7130 1520 0 otrip_decoded[7]
rlabel metal3 1096 6868 1096 6868 0 por_timed_out
rlabel metal1 6164 11322 6164 11322 0 por_unbuf
rlabel metal3 866 5508 866 5508 0 pwup_filt
rlabel metal2 9982 6987 9982 6987 0 startup_timed_out
<< properties >>
string FIXED_BBOX 0 0 11540 13684
<< end >>
