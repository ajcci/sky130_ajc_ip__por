magic
tech sky130A
magscale 1 2
timestamp 1714586768
<< error_s >>
rect 10454 -2676 10455 -2622
rect 10514 -2726 10515 -2676
rect 10514 -2996 10515 -2912
<< dnwell >>
rect -28958 13452 -6352 13820
rect -28958 499 -6351 13452
rect -5033 10587 -2433 13187
rect -28958 -5451 -10341 499
rect -5033 -184 -950 5889
rect -28958 -19950 12219 -5451
rect -28958 -24330 -16201 -19950
<< nwell >>
rect -29038 13614 -6271 13900
rect -29038 -24124 -28752 13614
rect -6558 705 -6271 13614
rect -5113 12981 -2353 13267
rect -5113 10793 -4827 12981
rect -2639 10793 -2353 12981
rect -5113 10507 -2353 10793
rect -10547 419 -6271 705
rect -5113 5683 -870 5969
rect -10547 -5371 -10261 419
rect -5113 22 -4827 5683
rect -4388 5340 -2380 5389
rect -4324 5319 -4293 5340
rect -2487 5319 -2456 5340
rect -4388 4513 -2380 4562
rect -4324 4492 -4293 4513
rect -2487 4492 -2456 4513
rect -4388 2364 -2380 2418
rect -4388 1615 -1920 1655
rect -1156 22 -870 5683
rect -5113 -264 -870 22
rect -10547 -5657 12299 -5371
rect 12013 -15596 12299 -5657
rect 12012 -19551 12299 -15596
rect 12012 -19721 12300 -19551
rect -16408 -20030 12300 -19721
rect -16408 -23396 -16121 -20030
rect -16407 -24124 -16121 -23396
rect -29038 -24410 -16121 -24124
<< pwell >>
rect -4339 4686 -2430 4779
rect -4339 3859 -2430 3952
rect -4380 1695 -2381 1803
rect -4339 936 -1970 1054
<< psubdiff >>
rect -4324 4740 -2456 4749
rect -4324 4706 -4279 4740
rect -2497 4706 -2456 4740
rect -4324 4696 -2456 4706
rect -4324 3913 -2456 3922
rect -4324 3879 -4279 3913
rect -2497 3879 -2456 3913
rect -4324 3869 -2456 3879
rect -4350 1726 -4272 1765
rect -2513 1726 -2418 1765
rect -4324 986 -4252 1020
rect -2051 986 -1996 1020
<< nsubdiff >>
rect -29001 13843 -6309 13863
rect -29001 13809 -28921 13843
rect -6415 13809 -6309 13843
rect -29001 13789 -6309 13809
rect -29001 13783 -28927 13789
rect -29001 -24293 -28981 13783
rect -28947 -24293 -28927 13783
rect -6383 13757 -6309 13789
rect -6383 536 -6363 13757
rect -6329 536 -6309 13757
rect -5076 13210 -2390 13230
rect -5076 13176 -4996 13210
rect -2470 13176 -2390 13210
rect -5076 13156 -2390 13176
rect -5076 13150 -5002 13156
rect -5076 10624 -5056 13150
rect -5022 10624 -5002 13150
rect -5076 10618 -5002 10624
rect -2464 13150 -2390 13156
rect -2464 10624 -2444 13150
rect -2410 10624 -2390 13150
rect -2464 10618 -2390 10624
rect -5076 10598 -2390 10618
rect -5076 10564 -4996 10598
rect -2470 10564 -2390 10598
rect -5076 10544 -2390 10564
rect -6383 530 -6309 536
rect -10372 510 -6309 530
rect -10372 476 -9897 510
rect -6389 476 -6309 510
rect -10372 456 -6309 476
rect -5076 5912 -907 5932
rect -5076 5878 -4996 5912
rect -987 5878 -907 5912
rect -5076 5858 -907 5878
rect -5076 5852 -5002 5858
rect -10372 189 -10298 456
rect -10372 -5328 -10352 189
rect -10318 -5328 -10298 189
rect -5076 -147 -5056 5852
rect -5022 -147 -5002 5852
rect -981 5852 -907 5858
rect -4324 5319 -4293 5353
rect -2487 5319 -2456 5353
rect -4324 4492 -4293 4526
rect -2487 4492 -2456 4526
rect -4350 2343 -4291 2382
rect -2491 2343 -2418 2382
rect -4350 1585 -4268 1619
rect -2004 1585 -1958 1619
rect -5076 -153 -5002 -147
rect -981 -147 -961 5852
rect -927 -147 -907 5852
rect -981 -153 -907 -147
rect -5076 -173 -907 -153
rect -5076 -207 -4996 -173
rect -987 -207 -907 -173
rect -5076 -227 -907 -207
rect -10372 -5408 -10298 -5328
rect -10372 -5428 12262 -5408
rect -10372 -5462 -10214 -5428
rect 12182 -5462 12262 -5428
rect -10372 -5482 12262 -5462
rect 12188 -5488 12262 -5482
rect 12188 -19839 12208 -5488
rect 12242 -19839 12262 -5488
rect -29001 -24299 -28927 -24293
rect -16232 -19915 -15757 -19895
rect 12188 -19896 12262 -19839
rect 11650 -19915 12262 -19896
rect -16232 -19949 -16152 -19915
rect 12182 -19949 12262 -19915
rect -16232 -19969 -15757 -19949
rect -16232 -19976 -16158 -19969
rect 11650 -19970 12262 -19949
rect -16232 -24270 -16212 -19976
rect -16178 -24270 -16158 -19976
rect -16232 -24299 -16158 -24270
rect -29001 -24319 -16158 -24299
rect -29001 -24353 -28921 -24319
rect -16232 -24353 -16158 -24319
rect -29001 -24373 -16158 -24353
<< psubdiffcont >>
rect -4279 4706 -2497 4740
rect -4279 3879 -2497 3913
rect -4272 1726 -2513 1765
rect -4252 986 -2051 1020
<< nsubdiffcont >>
rect -28921 13809 -6415 13843
rect -28981 -24293 -28947 13783
rect -6363 536 -6329 13757
rect -4996 13176 -2470 13210
rect -5056 10624 -5022 13150
rect -2444 10624 -2410 13150
rect -4996 10564 -2470 10598
rect -9897 476 -6389 510
rect -4996 5878 -987 5912
rect -10352 -5328 -10318 189
rect -5056 -147 -5022 5852
rect -4293 5319 -2487 5353
rect -4293 4492 -2487 4526
rect -4291 2343 -2491 2382
rect -4268 1585 -2004 1619
rect -961 -147 -927 5852
rect -4996 -207 -987 -173
rect -10214 -5462 12182 -5428
rect 12208 -19839 12242 -5488
rect -16152 -19949 12182 -19915
rect -16212 -24270 -16178 -19976
rect -28921 -24353 -16232 -24319
<< locali >>
rect -11148 11324 -11104 11358
rect -14959 9923 -14938 9957
rect -5056 13176 -4996 13210
rect -2470 13176 -2410 13210
rect -5056 13150 -5022 13176
rect -2444 13150 -2410 13176
rect -5056 10598 -5022 10624
rect -2444 10598 -2410 10624
rect -5056 10564 -4996 10598
rect -2470 10564 -2410 10598
rect -10352 476 -9897 510
rect -5056 5878 -4996 5912
rect -987 5878 -927 5912
rect -5056 5852 -5022 5878
rect -10352 189 -10318 476
rect -961 5852 -927 5878
rect -4350 5353 -2418 5359
rect -4350 5319 -4293 5353
rect -2487 5319 -2418 5353
rect -4350 5315 -2418 5319
rect -3916 4973 -3873 5021
rect -4324 4740 -2418 4741
rect -4324 4706 -4279 4740
rect -2497 4706 -2418 4740
rect -4324 4703 -2418 4706
rect -4350 4526 -2418 4532
rect -4350 4492 -4293 4526
rect -2487 4492 -2418 4526
rect -4350 4488 -2418 4492
rect -3916 4146 -3873 4194
rect -4324 3913 -2418 3914
rect -4324 3879 -4279 3913
rect -2497 3879 -2418 3913
rect -4324 3876 -2418 3879
rect -4350 2343 -4291 2382
rect -2491 2343 -2418 2382
rect -3916 1997 -3873 2045
rect -2588 1891 -2544 1915
rect -4350 1726 -4272 1765
rect -2513 1726 -2418 1765
rect -4350 1619 -1958 1625
rect -4350 1585 -4268 1619
rect -2004 1585 -1958 1619
rect -3916 1248 -3869 1298
rect -3456 1248 -3413 1296
rect -4314 986 -4252 1016
rect -2051 986 -1996 1016
rect -4314 970 -1996 986
rect -5056 -173 -5022 -147
rect -961 -173 -927 -147
rect -5056 -207 -4996 -173
rect -987 -207 -927 -173
rect -6515 -1210 -6451 -1195
rect -6515 -1308 -6500 -1210
rect -6466 -1308 -6451 -1210
rect -6515 -1323 -6451 -1308
rect -4403 -1210 -4339 -1195
rect -4403 -1308 -4388 -1210
rect -4354 -1308 -4339 -1210
rect -4403 -1323 -4339 -1308
rect -2291 -1210 -2227 -1195
rect -2291 -1308 -2276 -1210
rect -2242 -1308 -2227 -1210
rect -2291 -1323 -2227 -1308
rect -179 -1210 -115 -1195
rect -179 -1308 -164 -1210
rect -130 -1308 -115 -1210
rect -179 -1323 -115 -1308
rect 1933 -1210 1997 -1195
rect 1933 -1308 1948 -1210
rect 1982 -1308 1997 -1210
rect 1933 -1323 1997 -1308
rect 4045 -1210 4109 -1195
rect 4045 -1308 4060 -1210
rect 4094 -1308 4109 -1210
rect 4045 -1323 4109 -1308
rect 6157 -1210 6221 -1195
rect 6157 -1308 6172 -1210
rect 6206 -1308 6221 -1210
rect 6157 -1323 6221 -1308
rect 8269 -1210 8333 -1195
rect 8269 -1308 8284 -1210
rect 8318 -1308 8333 -1210
rect 8269 -1323 8333 -1308
rect 10381 -1210 10445 -1195
rect 10381 -1308 10396 -1210
rect 10430 -1308 10445 -1210
rect 10381 -1323 10445 -1308
rect 11174 -1843 11250 -1831
rect 11174 -1895 11186 -1843
rect 11238 -1895 11250 -1843
rect 11174 -1907 11250 -1895
rect -8047 -1942 -7983 -1927
rect -8047 -2040 -8032 -1942
rect -7998 -2040 -7983 -1942
rect -8047 -2055 -7983 -2040
rect -5935 -1942 -5871 -1927
rect -5935 -2040 -5920 -1942
rect -5886 -2040 -5871 -1942
rect -5935 -2055 -5871 -2040
rect -3823 -1942 -3759 -1927
rect -3823 -2040 -3808 -1942
rect -3774 -2040 -3759 -1942
rect -3823 -2055 -3759 -2040
rect -1711 -1942 -1647 -1927
rect -1711 -2040 -1696 -1942
rect -1662 -2040 -1647 -1942
rect -1711 -2055 -1647 -2040
rect 401 -1942 465 -1927
rect 401 -2040 416 -1942
rect 450 -2040 465 -1942
rect 401 -2055 465 -2040
rect 2513 -1942 2577 -1927
rect 2513 -2040 2528 -1942
rect 2562 -2040 2577 -1942
rect 2513 -2055 2577 -2040
rect 4625 -1942 4689 -1927
rect 4625 -2040 4640 -1942
rect 4674 -2040 4689 -1942
rect 4625 -2055 4689 -2040
rect 6737 -1942 6801 -1927
rect 6737 -2040 6752 -1942
rect 6786 -2040 6801 -1942
rect 6737 -2055 6801 -2040
rect 8849 -1942 8913 -1927
rect 8849 -2040 8864 -1942
rect 8898 -2040 8913 -1942
rect 8849 -2055 8913 -2040
rect -6515 -2944 -6451 -2929
rect -6515 -3042 -6500 -2944
rect -6466 -3042 -6451 -2944
rect -6515 -3057 -6451 -3042
rect -4403 -2944 -4339 -2929
rect -4403 -3042 -4388 -2944
rect -4354 -3042 -4339 -2944
rect -4403 -3057 -4339 -3042
rect -2291 -2944 -2227 -2929
rect -2291 -3042 -2276 -2944
rect -2242 -3042 -2227 -2944
rect -2291 -3057 -2227 -3042
rect -179 -2944 -115 -2929
rect -179 -3042 -164 -2944
rect -130 -3042 -115 -2944
rect -179 -3057 -115 -3042
rect 1933 -2944 1997 -2929
rect 1933 -3042 1948 -2944
rect 1982 -3042 1997 -2944
rect 1933 -3057 1997 -3042
rect 4045 -2944 4109 -2929
rect 4045 -3042 4060 -2944
rect 4094 -3042 4109 -2944
rect 4045 -3057 4109 -3042
rect 6157 -2944 6221 -2929
rect 6157 -3042 6172 -2944
rect 6206 -3042 6221 -2944
rect 6157 -3057 6221 -3042
rect 8269 -2944 8333 -2929
rect 8269 -3042 8284 -2944
rect 8318 -3042 8333 -2944
rect 8269 -3057 8333 -3042
rect 10381 -2944 10445 -2929
rect 10381 -3042 10396 -2944
rect 10430 -3042 10445 -2944
rect 10381 -3057 10445 -3042
rect -8047 -3676 -7983 -3661
rect -8047 -3774 -8032 -3676
rect -7998 -3774 -7983 -3676
rect -8047 -3789 -7983 -3774
rect -5935 -3676 -5871 -3661
rect -5935 -3774 -5920 -3676
rect -5886 -3774 -5871 -3676
rect -5935 -3789 -5871 -3774
rect -3823 -3676 -3759 -3661
rect -3823 -3774 -3808 -3676
rect -3774 -3774 -3759 -3676
rect -3823 -3789 -3759 -3774
rect -1711 -3676 -1647 -3661
rect -1711 -3774 -1696 -3676
rect -1662 -3774 -1647 -3676
rect -1711 -3789 -1647 -3774
rect 401 -3676 465 -3661
rect 401 -3774 416 -3676
rect 450 -3774 465 -3676
rect 401 -3789 465 -3774
rect 2513 -3676 2577 -3661
rect 2513 -3774 2528 -3676
rect 2562 -3774 2577 -3676
rect 2513 -3789 2577 -3774
rect 4625 -3676 4689 -3661
rect 4625 -3774 4640 -3676
rect 4674 -3774 4689 -3676
rect 4625 -3789 4689 -3774
rect 6737 -3676 6801 -3661
rect 6737 -3774 6752 -3676
rect 6786 -3774 6801 -3676
rect 6737 -3783 6801 -3774
rect 8849 -3676 8913 -3661
rect 8849 -3774 8864 -3676
rect 8898 -3774 8913 -3676
rect 8849 -3789 8913 -3774
<< viali >>
rect -28981 13809 -28921 13843
rect -28921 13809 -6415 13843
rect -6415 13809 -6329 13843
rect -28981 13783 -28947 13809
rect -28981 13370 -28947 13783
rect -29009 -11096 -28981 -10858
rect -28981 -24293 -28947 13164
rect -6363 13757 -6329 13809
rect -11358 11341 -11310 11389
rect -10510 11329 -10396 11370
rect -14938 9923 -7501 9957
rect -15129 1961 -15095 9861
rect -7439 1961 -7405 9861
rect -15033 1865 -7501 1899
rect -6363 536 -6329 13757
rect -4975 13176 -2503 13210
rect -5056 10624 -5022 13150
rect -3945 11686 -3570 11720
rect -3473 11521 -3405 11759
rect -2444 10624 -2410 13150
rect -4983 10564 -2486 10598
rect -2254 7677 -2208 7847
rect -3786 6982 -3738 7030
rect -6363 510 -6329 536
rect -9897 476 -6389 510
rect -6389 476 -6329 510
rect -10352 -5328 -10318 189
rect -5056 -147 -5022 5852
rect -4302 4975 -4254 5023
rect -2582 4863 -2548 5082
rect -4302 4148 -4254 4196
rect -2582 4036 -2548 4255
rect -4309 2003 -4065 2037
rect -2588 1915 -2544 2152
rect -4321 1254 -4188 1288
rect -2122 1149 -2088 1327
rect -961 -147 -927 5852
rect -6500 -1308 -6466 -1210
rect -4388 -1308 -4354 -1210
rect -2276 -1308 -2242 -1210
rect -164 -1308 -130 -1210
rect 1948 -1308 1982 -1210
rect 4060 -1308 4094 -1210
rect 6172 -1308 6206 -1210
rect 8284 -1308 8318 -1210
rect 10396 -1308 10430 -1210
rect 10642 -1378 10690 -1330
rect 11186 -1895 11238 -1843
rect -8032 -2040 -7998 -1942
rect -5920 -2040 -5886 -1942
rect -3808 -2040 -3774 -1942
rect -1696 -2040 -1662 -1942
rect 416 -2040 450 -1942
rect 2528 -2040 2562 -1942
rect 4640 -2040 4674 -1942
rect 6752 -2040 6786 -1942
rect 8864 -2040 8898 -1942
rect -6500 -3042 -6466 -2944
rect -4388 -3042 -4354 -2944
rect -2276 -3042 -2242 -2944
rect -164 -3042 -130 -2944
rect 1948 -3042 1982 -2944
rect 4060 -3042 4094 -2944
rect 6172 -3042 6206 -2944
rect 8284 -3042 8318 -2944
rect 10396 -3042 10430 -2944
rect 10642 -3114 10694 -3062
rect 11203 -3642 11251 -3594
rect -8032 -3774 -7998 -3676
rect -5920 -3774 -5886 -3676
rect -3808 -3774 -3774 -3676
rect -1696 -3774 -1662 -3676
rect 416 -3774 450 -3676
rect 2528 -3774 2562 -3676
rect 4640 -3774 4674 -3676
rect 6752 -3774 6786 -3676
rect 8864 -3774 8898 -3676
rect -10352 -5428 -10318 -5328
rect -10352 -5462 -10214 -5428
rect -10214 -5462 12182 -5428
rect 12182 -5462 12242 -5428
rect 12208 -5488 12242 -5462
rect -28947 -11096 -28771 -10858
rect 12208 -19839 12242 -5488
rect 12208 -19915 12242 -19839
rect -28981 -24319 -28947 -24293
rect -16212 -19949 -16152 -19915
rect -16152 -19949 12182 -19915
rect 12182 -19949 12242 -19915
rect -16212 -19976 -16178 -19949
rect -16212 -24270 -16178 -19976
rect -16212 -24319 -16178 -24270
rect -28981 -24353 -28921 -24319
rect -28921 -24353 -16232 -24319
rect -16232 -24353 -16178 -24319
<< metal1 >>
rect -29001 13843 -6309 13863
rect -29001 13370 -28981 13843
rect -28947 13789 -6363 13809
rect -28947 13370 -28927 13789
rect -29001 13365 -28927 13370
rect -29001 13359 -28751 13365
rect -29001 13211 -28905 13359
rect -28757 13211 -28751 13359
rect -29001 13205 -28751 13211
rect -29001 13164 -28927 13205
rect -29001 -10852 -28981 13164
rect -29021 -10858 -28981 -10852
rect -28947 -10852 -28927 13164
rect -11077 11696 -11071 11844
rect -10923 11696 -10917 11844
rect -8185 11513 -7927 11519
rect -8185 11461 -8179 11513
rect -7933 11461 -7927 11513
rect -8185 11455 -7927 11461
rect -11370 11335 -11364 11395
rect -11304 11335 -11298 11395
rect -10522 11377 -10386 11382
rect -10522 11370 -9993 11377
rect -10522 11329 -10510 11370
rect -10396 11329 -9993 11370
rect -10522 11321 -9993 11329
rect -10522 11317 -10386 11321
rect -15370 10989 -15364 11137
rect -15216 10989 -7665 11137
rect -15135 9957 -7398 9963
rect -15135 9923 -14938 9957
rect -7501 9923 -7398 9957
rect -15135 9917 -7398 9923
rect -15135 9861 -15089 9917
rect -15135 8025 -15129 9861
rect -15155 8016 -15129 8025
rect -15095 8025 -15089 9861
rect -7445 9861 -7398 9917
rect -14727 9400 -14611 9821
rect -13971 9400 -13855 9821
rect -13215 9400 -13099 9821
rect -12459 9400 -12343 9821
rect -11703 9400 -11587 9821
rect -10947 9400 -10831 9821
rect -10191 9400 -10075 9821
rect -9435 9400 -9319 9821
rect -8679 9400 -8563 9821
rect -7923 9400 -7807 9821
rect -15095 8016 -15081 8025
rect -15155 7886 -15146 8016
rect -15090 7886 -15081 8016
rect -15155 7877 -15129 7886
rect -15135 1961 -15129 7877
rect -15095 7877 -15081 7886
rect -15095 1961 -15089 7877
rect -14892 2023 -14886 2087
rect -14822 2023 -14816 2087
rect -14349 2001 -14233 2422
rect -13593 2001 -13477 2422
rect -12837 2001 -12721 2422
rect -12081 2001 -11965 2422
rect -11325 2001 -11209 2422
rect -10569 2001 -10453 2422
rect -9813 2001 -9697 2422
rect -9057 2001 -8941 2422
rect -8301 2001 -8185 2422
rect -7731 2013 -7725 2107
rect -7621 2013 -7615 2107
rect -15135 1905 -15089 1961
rect -7445 1961 -7439 9861
rect -7405 1961 -7398 9861
rect -7445 1905 -7398 1961
rect -15135 1899 -7398 1905
rect -15135 1865 -15033 1899
rect -7501 1865 -7398 1899
rect -15135 1859 -7398 1865
rect -6383 530 -6363 13789
rect -10372 510 -6363 530
rect -10372 476 -9897 510
rect -6329 476 -6309 13843
rect -5076 13210 -2390 13230
rect -5076 13176 -4975 13210
rect -2503 13176 -2390 13210
rect -5076 13156 -2390 13176
rect -5076 13150 -5002 13156
rect -5076 10624 -5056 13150
rect -5022 10624 -5002 13150
rect -2464 13150 -2390 13156
rect -3842 11944 -3676 11959
rect -3842 11808 -3827 11944
rect -3691 11808 -3676 11944
rect -3842 11793 -3676 11808
rect -3488 11898 -3387 11904
rect -3488 11759 -3387 11797
rect -3488 11739 -3473 11759
rect -3968 11720 -3473 11739
rect -3968 11686 -3945 11720
rect -3570 11686 -3473 11720
rect -3968 11667 -3473 11686
rect -3488 11521 -3473 11667
rect -3405 11577 -3387 11759
rect -2464 11577 -2444 13150
rect -3405 11521 -2444 11577
rect -3488 11504 -3387 11521
rect -5076 10618 -5002 10624
rect -2464 10624 -2444 11521
rect -2410 10624 -2390 13150
rect -2464 10618 -2390 10624
rect -5076 10598 -2390 10618
rect -5076 10564 -4983 10598
rect -2486 10564 -2390 10598
rect -5076 10544 -2390 10564
rect -4713 8156 -4707 8284
rect -4579 8156 -2170 8284
rect -2266 7847 -2196 7860
rect -2266 7795 -2254 7847
rect -2208 7795 -2196 7847
rect -2266 7739 -2260 7795
rect -2204 7739 -2196 7795
rect -2266 7677 -2254 7739
rect -2208 7677 -2196 7739
rect -2266 7665 -2196 7677
rect -4282 7529 -2172 7572
rect -5322 7401 -5316 7529
rect -5188 7401 -2172 7529
rect -4282 7327 -2172 7401
rect -4912 7242 -4906 7299
rect -4849 7242 -4174 7299
rect -3798 7036 -3726 7042
rect -3798 6976 -3792 7036
rect -3732 6976 -3726 7036
rect -3798 6970 -3726 6976
rect -4713 6743 -4579 6749
rect -4713 6615 -4707 6743
rect -4579 6615 -2170 6743
rect -4713 6609 -4579 6615
rect -10372 456 -6309 476
rect -5076 5858 -907 5932
rect -5076 5852 -5002 5858
rect -10372 189 -10298 456
rect -10372 -5462 -10352 189
rect -10318 -5408 -10298 189
rect -5076 -147 -5056 5852
rect -5022 2375 -5002 5852
rect -981 5852 -907 5858
rect -4893 5254 -4887 5350
rect -4791 5254 -4350 5350
rect -2598 5082 -2532 5091
rect -4314 5029 -4242 5035
rect -4314 4969 -4308 5029
rect -4248 4969 -4242 5029
rect -4314 4963 -4242 4969
rect -2598 4859 -2590 5082
rect -2538 4859 -2532 5082
rect -2598 4853 -2532 4859
rect -4690 4710 -4684 4806
rect -4588 4710 -4350 4806
rect -4897 4427 -4891 4523
rect -4795 4427 -4350 4523
rect -2598 4255 -2532 4264
rect -4314 4202 -4242 4208
rect -4314 4142 -4308 4202
rect -4248 4142 -4242 4202
rect -4314 4136 -4242 4142
rect -2598 4032 -2590 4255
rect -2538 4032 -2532 4255
rect -2598 4026 -2532 4032
rect -4694 3883 -4688 3979
rect -4592 3883 -4350 3979
rect -4907 3699 -4448 3705
rect -4907 3540 -4899 3699
rect -4785 3540 -4448 3699
rect -4907 3533 -4448 3540
rect -4707 3054 -4420 3059
rect -4707 2897 -4698 3054
rect -4588 2897 -4420 3054
rect -4707 2890 -4420 2897
rect -5022 2374 -4907 2375
rect -5022 2363 -4350 2374
rect -5022 2287 -4898 2363
rect -4791 2287 -4350 2363
rect -5022 2278 -4350 2287
rect -5022 -147 -5002 2278
rect -2594 2153 -2538 2165
rect -4324 2037 -4117 2052
rect -4324 2003 -4309 2037
rect -4324 1992 -4117 2003
rect -4057 1992 -4051 2052
rect -2594 1885 -2538 1898
rect -4707 1824 -4350 1830
rect -4707 1740 -4699 1824
rect -4587 1740 -4350 1824
rect -4707 1734 -4350 1740
rect -4901 1529 -4895 1625
rect -4799 1529 -4350 1625
rect -2138 1334 -2072 1343
rect -4333 1297 -4176 1303
rect -4333 1245 -4327 1297
rect -4184 1245 -4176 1297
rect -4333 1239 -4176 1245
rect -2138 1142 -2130 1334
rect -2078 1142 -2072 1334
rect -2138 1134 -2072 1142
rect -4701 985 -4695 1081
rect -4599 985 -4314 1081
rect -5076 -153 -5002 -147
rect -981 -147 -961 5852
rect -927 -147 -907 5852
rect -981 -153 -907 -147
rect -9058 -350 -9052 -222
rect -8924 -350 -5316 -222
rect -5188 -350 -5182 -222
rect -5076 -227 -907 -153
rect -9258 -593 -9252 -465
rect -9124 -466 -5636 -465
rect -9124 -593 -4907 -466
rect -5762 -594 -4907 -593
rect -4779 -594 -4773 -466
rect -8852 -718 -6055 -712
rect -8852 -854 -8846 -718
rect -8730 -724 -6055 -718
rect -5918 -724 12117 -712
rect -8730 -728 12117 -724
rect -8730 -854 -4707 -728
rect -8852 -856 -4707 -854
rect -4579 -856 12117 -728
rect -8852 -860 12117 -856
rect -6515 -1201 -6451 -1195
rect -6515 -1317 -6509 -1201
rect -6457 -1317 -6451 -1201
rect -6515 -1323 -6451 -1317
rect -4403 -1201 -4339 -1195
rect -4403 -1317 -4397 -1201
rect -4345 -1317 -4339 -1201
rect -4403 -1323 -4339 -1317
rect -2291 -1201 -2227 -1195
rect -2291 -1317 -2285 -1201
rect -2233 -1317 -2227 -1201
rect -2291 -1323 -2227 -1317
rect -179 -1201 -115 -1195
rect -179 -1317 -173 -1201
rect -121 -1317 -115 -1201
rect -179 -1323 -115 -1317
rect 1933 -1201 1997 -1195
rect 1933 -1317 1939 -1201
rect 1991 -1317 1997 -1201
rect 1933 -1323 1997 -1317
rect 4045 -1201 4109 -1195
rect 4045 -1317 4051 -1201
rect 4103 -1317 4109 -1201
rect 4045 -1323 4109 -1317
rect 6157 -1201 6221 -1195
rect 6157 -1317 6163 -1201
rect 6215 -1317 6221 -1201
rect 6157 -1323 6221 -1317
rect 8269 -1201 8333 -1195
rect 8269 -1317 8275 -1201
rect 8327 -1317 8333 -1201
rect 8269 -1323 8333 -1317
rect 10381 -1201 10445 -1195
rect 10381 -1317 10387 -1201
rect 10439 -1317 10445 -1201
rect 10381 -1323 10445 -1317
rect 10630 -1384 10636 -1324
rect 10696 -1384 10702 -1324
rect -9052 -1430 12117 -1424
rect -9052 -1668 -9046 -1430
rect -8930 -1668 12117 -1430
rect -9052 -1674 12117 -1668
rect -9252 -1704 12099 -1702
rect -9252 -1756 -9246 -1704
rect -9130 -1756 12099 -1704
rect -9252 -1759 12099 -1756
rect 11174 -1837 11250 -1831
rect 11174 -1901 11180 -1837
rect 11244 -1901 11250 -1837
rect 11174 -1907 11250 -1901
rect -8047 -1933 -7983 -1927
rect -8047 -2049 -8041 -1933
rect -7989 -2049 -7983 -1933
rect -8047 -2055 -7983 -2049
rect -5935 -1933 -5871 -1927
rect -5935 -2049 -5929 -1933
rect -5877 -2049 -5871 -1933
rect -5935 -2055 -5871 -2049
rect -3823 -1933 -3759 -1927
rect -3823 -2049 -3817 -1933
rect -3765 -2049 -3759 -1933
rect -3823 -2055 -3759 -2049
rect -1711 -1933 -1647 -1927
rect -1711 -2049 -1705 -1933
rect -1653 -2049 -1647 -1933
rect -1711 -2055 -1647 -2049
rect 401 -1933 465 -1927
rect 401 -2049 407 -1933
rect 459 -2049 465 -1933
rect 401 -2055 465 -2049
rect 2513 -1933 2577 -1927
rect 2513 -2049 2519 -1933
rect 2571 -2049 2577 -1933
rect 2513 -2055 2577 -2049
rect 4625 -1933 4689 -1927
rect 4625 -2049 4631 -1933
rect 4683 -2049 4689 -1933
rect 4625 -2055 4689 -2049
rect 6737 -1933 6801 -1927
rect 6737 -2049 6743 -1933
rect 6795 -2049 6801 -1933
rect 6737 -2055 6801 -2049
rect 8849 -1933 8913 -1927
rect 8849 -2049 8855 -1933
rect 8907 -2049 8913 -1933
rect 8849 -2055 8913 -2049
rect -8852 -2242 12117 -2238
rect -8852 -2244 4625 -2242
rect -8852 -2588 -8846 -2244
rect -8730 -2246 4625 -2244
rect -8730 -2310 401 -2246
rect 465 -2248 4625 -2246
rect 465 -2310 2513 -2248
rect -8730 -2312 2513 -2310
rect 2577 -2306 4625 -2248
rect 4689 -2248 12117 -2242
rect 4689 -2306 6737 -2248
rect 2577 -2312 6737 -2306
rect 6801 -2312 12117 -2248
rect -8730 -2588 12117 -2312
rect -8852 -2594 12117 -2588
rect -6515 -2935 -6451 -2929
rect -6515 -3051 -6509 -2935
rect -6457 -3051 -6451 -2935
rect -6515 -3057 -6451 -3051
rect -4403 -2935 -4339 -2929
rect -4403 -3051 -4397 -2935
rect -4345 -3051 -4339 -2935
rect -4403 -3057 -4339 -3051
rect -2291 -2935 -2227 -2929
rect -2291 -3051 -2285 -2935
rect -2233 -3051 -2227 -2935
rect -2291 -3057 -2227 -3051
rect -179 -2935 -115 -2929
rect -179 -3051 -173 -2935
rect -121 -3051 -115 -2935
rect -179 -3057 -115 -3051
rect 1933 -2935 1997 -2929
rect 1933 -3051 1939 -2935
rect 1991 -3051 1997 -2935
rect 1933 -3057 1997 -3051
rect 4045 -2935 4109 -2929
rect 4045 -3051 4051 -2935
rect 4103 -3051 4109 -2935
rect 4045 -3057 4109 -3051
rect 6157 -2935 6221 -2929
rect 6157 -3051 6163 -2935
rect 6215 -3051 6221 -2935
rect 6157 -3057 6221 -3051
rect 8269 -2935 8333 -2929
rect 8269 -3051 8275 -2935
rect 8327 -3051 8333 -2935
rect 8269 -3057 8333 -3051
rect 10381 -2935 10445 -2929
rect 10381 -3051 10387 -2935
rect 10439 -3051 10445 -2935
rect 10381 -3057 10445 -3051
rect 10630 -3120 10636 -3056
rect 10700 -3120 10706 -3056
rect -9052 -3164 12117 -3158
rect -9052 -3402 -9046 -3164
rect -8930 -3402 12117 -3164
rect -9052 -3408 12117 -3402
rect -9252 -3438 12117 -3436
rect -9252 -3490 -9246 -3438
rect -9130 -3490 12117 -3438
rect -9252 -3493 12117 -3490
rect 11191 -3648 11197 -3588
rect 11257 -3648 11263 -3588
rect -8047 -3667 -7983 -3661
rect -8047 -3783 -8041 -3667
rect -7989 -3783 -7983 -3667
rect -8047 -3789 -7983 -3783
rect -5935 -3667 -5871 -3661
rect -5935 -3783 -5929 -3667
rect -5877 -3783 -5871 -3667
rect -5935 -3789 -5871 -3783
rect -3823 -3667 -3759 -3661
rect -3823 -3783 -3817 -3667
rect -3765 -3783 -3759 -3667
rect -3823 -3789 -3759 -3783
rect -1711 -3667 -1647 -3661
rect -1711 -3783 -1705 -3667
rect -1653 -3783 -1647 -3667
rect -1711 -3789 -1647 -3783
rect 401 -3667 465 -3661
rect 401 -3783 407 -3667
rect 459 -3783 465 -3667
rect 401 -3789 465 -3783
rect 2513 -3667 2577 -3661
rect 2513 -3783 2519 -3667
rect 2571 -3783 2577 -3667
rect 2513 -3789 2577 -3783
rect 4625 -3667 4689 -3661
rect 4625 -3783 4631 -3667
rect 4683 -3783 4689 -3667
rect 6737 -3667 6801 -3661
rect 6737 -3783 6743 -3667
rect 6795 -3783 6801 -3667
rect 8849 -3667 8913 -3661
rect 8849 -3783 8855 -3667
rect 8907 -3783 8913 -3667
rect 4625 -3789 4689 -3783
rect 8849 -3789 8913 -3783
rect 395 -3972 401 -3970
rect -8852 -3978 401 -3972
rect -8852 -4082 -8846 -3978
rect -9252 -4114 -8846 -4082
rect -8730 -4034 401 -3978
rect 465 -3972 471 -3970
rect 465 -3980 12117 -3972
rect 465 -3984 6737 -3980
rect 465 -4034 2513 -3984
rect -8730 -4048 2513 -4034
rect 2577 -4048 4625 -3984
rect 4689 -4036 6737 -3984
rect 6793 -4036 12117 -3980
rect 4689 -4048 12117 -4036
rect -8730 -4114 12117 -4048
rect -9252 -4282 12117 -4114
rect -9252 -4344 10468 -4338
rect -9252 -4532 -9246 -4344
rect -9130 -4532 10468 -4344
rect -9252 -4538 10468 -4532
rect -9252 -4600 10468 -4594
rect -9252 -4788 -9046 -4600
rect -8930 -4788 10468 -4600
rect -9252 -4794 10468 -4788
rect -4837 -5408 -4637 -4794
rect -10318 -5428 12262 -5408
rect -10372 -5482 12208 -5462
rect -4837 -6994 -4637 -5482
rect -27806 -10519 -27406 -10513
rect -27806 -10796 -27800 -10519
rect -27412 -10796 -27406 -10519
rect -27806 -10802 -27406 -10796
rect -19274 -10802 -10164 -10552
rect -10355 -10824 -10164 -10802
rect -10355 -10830 -4887 -10824
rect -28947 -10858 -27459 -10852
rect -29021 -11096 -29009 -10858
rect -28771 -11096 -28256 -10858
rect -27868 -11096 -27459 -10858
rect -29021 -11102 -28981 -11096
rect -29001 -24353 -28981 -11102
rect -28947 -11102 -27459 -11096
rect -19020 -11080 -10420 -10854
rect -10355 -11018 -5076 -10830
rect -4893 -11018 -4887 -10830
rect -10355 -11024 -4887 -11018
rect -28947 -24299 -28927 -11102
rect -19020 -11104 -4637 -11080
rect -10614 -11280 -4637 -11104
rect 12188 -19896 12208 -5482
rect -16232 -19915 12208 -19896
rect -16232 -24299 -16212 -19915
rect 12242 -19949 12262 -5428
rect -28947 -24319 -16212 -24299
rect -16178 -19969 12262 -19949
rect -16178 -24353 -16158 -19969
rect 11650 -19970 12262 -19969
rect -10867 -21963 -10766 -21957
rect -10867 -22052 -10861 -21963
rect -10772 -22052 -10766 -21963
rect -10867 -22058 -10766 -22052
rect -10549 -22947 -10409 -22941
rect -10549 -23075 -10543 -22947
rect -10415 -23075 -10409 -22947
rect -10549 -23081 -10409 -23075
rect -29001 -24373 -16158 -24353
<< via1 >>
rect -28905 13211 -28757 13359
rect -11071 11696 -10923 11844
rect -8179 11461 -7933 11513
rect -11364 11389 -11304 11395
rect -11364 11341 -11358 11389
rect -11358 11341 -11310 11389
rect -11310 11341 -11304 11389
rect -11364 11335 -11304 11341
rect -15364 10989 -15216 11137
rect -15146 7886 -15129 8016
rect -15129 7886 -15095 8016
rect -15095 7886 -15090 8016
rect -14886 2023 -14822 2087
rect -7725 2013 -7621 2107
rect -3827 11808 -3691 11944
rect -3488 11797 -3387 11898
rect -4707 8156 -4579 8284
rect -2260 7739 -2254 7795
rect -2254 7739 -2208 7795
rect -2208 7739 -2204 7795
rect -5316 7401 -5188 7529
rect -4906 7242 -4849 7299
rect -3792 7030 -3732 7036
rect -3792 6982 -3786 7030
rect -3786 6982 -3738 7030
rect -3738 6982 -3732 7030
rect -3792 6976 -3732 6982
rect -4707 6615 -4579 6743
rect -4887 5254 -4791 5350
rect -4308 5023 -4248 5029
rect -4308 4975 -4302 5023
rect -4302 4975 -4254 5023
rect -4254 4975 -4248 5023
rect -4308 4969 -4248 4975
rect -2590 4863 -2582 5082
rect -2582 4863 -2548 5082
rect -2548 4863 -2538 5082
rect -2590 4859 -2538 4863
rect -4684 4710 -4588 4806
rect -4891 4427 -4795 4523
rect -4308 4196 -4248 4202
rect -4308 4148 -4302 4196
rect -4302 4148 -4254 4196
rect -4254 4148 -4248 4196
rect -4308 4142 -4248 4148
rect -2590 4036 -2582 4255
rect -2582 4036 -2548 4255
rect -2548 4036 -2538 4255
rect -2590 4032 -2538 4036
rect -4688 3883 -4592 3979
rect -4899 3540 -4785 3699
rect -4698 2897 -4588 3054
rect -4898 2287 -4791 2363
rect -2594 2152 -2538 2153
rect -4117 2037 -4057 2052
rect -4117 2003 -4065 2037
rect -4065 2003 -4057 2037
rect -4117 1992 -4057 2003
rect -2594 1915 -2588 2152
rect -2588 1915 -2544 2152
rect -2544 1915 -2538 2152
rect -2594 1898 -2538 1915
rect -4699 1740 -4587 1824
rect -4895 1529 -4799 1625
rect -4327 1288 -4184 1297
rect -4327 1254 -4321 1288
rect -4321 1254 -4188 1288
rect -4188 1254 -4184 1288
rect -4327 1245 -4184 1254
rect -2130 1327 -2078 1334
rect -2130 1149 -2122 1327
rect -2122 1149 -2088 1327
rect -2088 1149 -2078 1327
rect -2130 1142 -2078 1149
rect -4695 985 -4599 1081
rect -9052 -350 -8924 -222
rect -5316 -350 -5188 -222
rect -9252 -593 -9124 -465
rect -4907 -594 -4779 -466
rect -8846 -854 -8730 -718
rect -4707 -856 -4579 -728
rect -6509 -1210 -6457 -1201
rect -6509 -1308 -6500 -1210
rect -6500 -1308 -6466 -1210
rect -6466 -1308 -6457 -1210
rect -6509 -1317 -6457 -1308
rect -4397 -1210 -4345 -1201
rect -4397 -1308 -4388 -1210
rect -4388 -1308 -4354 -1210
rect -4354 -1308 -4345 -1210
rect -4397 -1317 -4345 -1308
rect -2285 -1210 -2233 -1201
rect -2285 -1308 -2276 -1210
rect -2276 -1308 -2242 -1210
rect -2242 -1308 -2233 -1210
rect -2285 -1317 -2233 -1308
rect -173 -1210 -121 -1201
rect -173 -1308 -164 -1210
rect -164 -1308 -130 -1210
rect -130 -1308 -121 -1210
rect -173 -1317 -121 -1308
rect 1939 -1210 1991 -1201
rect 1939 -1308 1948 -1210
rect 1948 -1308 1982 -1210
rect 1982 -1308 1991 -1210
rect 1939 -1317 1991 -1308
rect 4051 -1210 4103 -1201
rect 4051 -1308 4060 -1210
rect 4060 -1308 4094 -1210
rect 4094 -1308 4103 -1210
rect 4051 -1317 4103 -1308
rect 6163 -1210 6215 -1201
rect 6163 -1308 6172 -1210
rect 6172 -1308 6206 -1210
rect 6206 -1308 6215 -1210
rect 6163 -1317 6215 -1308
rect 8275 -1210 8327 -1201
rect 8275 -1308 8284 -1210
rect 8284 -1308 8318 -1210
rect 8318 -1308 8327 -1210
rect 8275 -1317 8327 -1308
rect 10387 -1210 10439 -1201
rect 10387 -1308 10396 -1210
rect 10396 -1308 10430 -1210
rect 10430 -1308 10439 -1210
rect 10387 -1317 10439 -1308
rect 10636 -1330 10696 -1324
rect 10636 -1378 10642 -1330
rect 10642 -1378 10690 -1330
rect 10690 -1378 10696 -1330
rect 10636 -1384 10696 -1378
rect -9046 -1668 -8930 -1430
rect -9246 -1756 -9130 -1704
rect 11180 -1843 11244 -1837
rect 11180 -1895 11186 -1843
rect 11186 -1895 11238 -1843
rect 11238 -1895 11244 -1843
rect 11180 -1901 11244 -1895
rect -8041 -1942 -7989 -1933
rect -8041 -2040 -8032 -1942
rect -8032 -2040 -7998 -1942
rect -7998 -2040 -7989 -1942
rect -8041 -2049 -7989 -2040
rect -5929 -1942 -5877 -1933
rect -5929 -2040 -5920 -1942
rect -5920 -2040 -5886 -1942
rect -5886 -2040 -5877 -1942
rect -5929 -2049 -5877 -2040
rect -3817 -1942 -3765 -1933
rect -3817 -2040 -3808 -1942
rect -3808 -2040 -3774 -1942
rect -3774 -2040 -3765 -1942
rect -3817 -2049 -3765 -2040
rect -1705 -1942 -1653 -1933
rect -1705 -2040 -1696 -1942
rect -1696 -2040 -1662 -1942
rect -1662 -2040 -1653 -1942
rect -1705 -2049 -1653 -2040
rect 407 -1942 459 -1933
rect 407 -2040 416 -1942
rect 416 -2040 450 -1942
rect 450 -2040 459 -1942
rect 407 -2049 459 -2040
rect 2519 -1942 2571 -1933
rect 2519 -2040 2528 -1942
rect 2528 -2040 2562 -1942
rect 2562 -2040 2571 -1942
rect 2519 -2049 2571 -2040
rect 4631 -1942 4683 -1933
rect 4631 -2040 4640 -1942
rect 4640 -2040 4674 -1942
rect 4674 -2040 4683 -1942
rect 4631 -2049 4683 -2040
rect 6743 -1942 6795 -1933
rect 6743 -2040 6752 -1942
rect 6752 -2040 6786 -1942
rect 6786 -2040 6795 -1942
rect 6743 -2049 6795 -2040
rect 8855 -1942 8907 -1933
rect 8855 -2040 8864 -1942
rect 8864 -2040 8898 -1942
rect 8898 -2040 8907 -1942
rect 8855 -2049 8907 -2040
rect -8846 -2588 -8730 -2244
rect 401 -2310 465 -2246
rect 2513 -2312 2577 -2248
rect 4625 -2306 4689 -2242
rect 6737 -2312 6801 -2248
rect -6509 -2944 -6457 -2935
rect -6509 -3042 -6500 -2944
rect -6500 -3042 -6466 -2944
rect -6466 -3042 -6457 -2944
rect -6509 -3051 -6457 -3042
rect -4397 -2944 -4345 -2935
rect -4397 -3042 -4388 -2944
rect -4388 -3042 -4354 -2944
rect -4354 -3042 -4345 -2944
rect -4397 -3051 -4345 -3042
rect -2285 -2944 -2233 -2935
rect -2285 -3042 -2276 -2944
rect -2276 -3042 -2242 -2944
rect -2242 -3042 -2233 -2944
rect -2285 -3051 -2233 -3042
rect -173 -2944 -121 -2935
rect -173 -3042 -164 -2944
rect -164 -3042 -130 -2944
rect -130 -3042 -121 -2944
rect -173 -3051 -121 -3042
rect 1939 -2944 1991 -2935
rect 1939 -3042 1948 -2944
rect 1948 -3042 1982 -2944
rect 1982 -3042 1991 -2944
rect 1939 -3051 1991 -3042
rect 4051 -2944 4103 -2935
rect 4051 -3042 4060 -2944
rect 4060 -3042 4094 -2944
rect 4094 -3042 4103 -2944
rect 4051 -3051 4103 -3042
rect 6163 -2944 6215 -2935
rect 6163 -3042 6172 -2944
rect 6172 -3042 6206 -2944
rect 6206 -3042 6215 -2944
rect 6163 -3051 6215 -3042
rect 8275 -2944 8327 -2935
rect 8275 -3042 8284 -2944
rect 8284 -3042 8318 -2944
rect 8318 -3042 8327 -2944
rect 8275 -3051 8327 -3042
rect 10387 -2944 10439 -2935
rect 10387 -3042 10396 -2944
rect 10396 -3042 10430 -2944
rect 10430 -3042 10439 -2944
rect 10387 -3051 10439 -3042
rect 10636 -3062 10700 -3056
rect 10636 -3114 10642 -3062
rect 10642 -3114 10694 -3062
rect 10694 -3114 10700 -3062
rect 10636 -3120 10700 -3114
rect -9046 -3402 -8930 -3164
rect -9246 -3490 -9130 -3438
rect 11197 -3594 11257 -3588
rect 11197 -3642 11203 -3594
rect 11203 -3642 11251 -3594
rect 11251 -3642 11257 -3594
rect 11197 -3648 11257 -3642
rect -8041 -3676 -7989 -3667
rect -8041 -3774 -8032 -3676
rect -8032 -3774 -7998 -3676
rect -7998 -3774 -7989 -3676
rect -8041 -3783 -7989 -3774
rect -5929 -3676 -5877 -3667
rect -5929 -3774 -5920 -3676
rect -5920 -3774 -5886 -3676
rect -5886 -3774 -5877 -3676
rect -5929 -3783 -5877 -3774
rect -3817 -3676 -3765 -3667
rect -3817 -3774 -3808 -3676
rect -3808 -3774 -3774 -3676
rect -3774 -3774 -3765 -3676
rect -3817 -3783 -3765 -3774
rect -1705 -3676 -1653 -3667
rect -1705 -3774 -1696 -3676
rect -1696 -3774 -1662 -3676
rect -1662 -3774 -1653 -3676
rect -1705 -3783 -1653 -3774
rect 407 -3676 459 -3667
rect 407 -3774 416 -3676
rect 416 -3774 450 -3676
rect 450 -3774 459 -3676
rect 407 -3783 459 -3774
rect 2519 -3676 2571 -3667
rect 2519 -3774 2528 -3676
rect 2528 -3774 2562 -3676
rect 2562 -3774 2571 -3676
rect 2519 -3783 2571 -3774
rect 4631 -3676 4683 -3667
rect 4631 -3774 4640 -3676
rect 4640 -3774 4674 -3676
rect 4674 -3774 4683 -3676
rect 4631 -3783 4683 -3774
rect 6743 -3676 6795 -3667
rect 6743 -3774 6752 -3676
rect 6752 -3774 6786 -3676
rect 6786 -3774 6795 -3676
rect 6743 -3783 6795 -3774
rect 8855 -3676 8907 -3667
rect 8855 -3774 8864 -3676
rect 8864 -3774 8898 -3676
rect 8898 -3774 8907 -3676
rect 8855 -3783 8907 -3774
rect -8846 -4114 -8730 -3978
rect 401 -4034 465 -3970
rect 2513 -4048 2577 -3984
rect 4625 -4048 4689 -3984
rect 6737 -4036 6793 -3980
rect -9246 -4532 -9130 -4344
rect -9046 -4788 -8930 -4600
rect -27800 -10796 -27412 -10519
rect -28256 -11096 -27868 -10858
rect -5076 -11018 -4893 -10830
rect -4575 -11018 -4387 -10830
rect -10861 -22052 -10772 -21963
rect -10543 -23075 -10415 -22947
<< metal2 >>
rect -27525 13694 -27434 13698
rect -3488 13695 -3387 13701
rect -27529 13689 -27428 13694
rect -27529 13598 -27525 13689
rect -27434 13598 -27428 13689
rect -27529 13433 -27428 13598
rect -3497 13592 -3488 13695
rect -3387 13592 -3378 13695
rect -23906 13490 -23850 13497
rect -3844 13490 -3784 13499
rect -23908 13488 -23848 13490
rect -28911 13359 -28751 13365
rect -28911 13211 -28905 13359
rect -28757 13211 -28751 13359
rect -28911 13205 -28751 13211
rect -28262 13353 -27862 13433
rect -28262 13217 -27929 13353
rect -27868 13217 -27862 13353
rect -28262 -10858 -27862 13217
rect -28262 -10926 -28256 -10858
rect -29373 -11096 -28256 -10926
rect -27868 -11096 -27862 -10858
rect -29373 -11326 -27862 -11096
rect -27806 8019 -27406 13433
rect -23908 13432 -23906 13488
rect -23850 13432 -23848 13488
rect -27042 8356 -26986 8365
rect -27042 8291 -26986 8300
rect -27806 7883 -27478 8019
rect -27412 7883 -27406 8019
rect -27806 1922 -27406 7883
rect -27806 1786 -27478 1922
rect -27412 1786 -27406 1922
rect -27806 -10519 -27406 1786
rect -26907 525 -26851 532
rect -27806 -10796 -27800 -10519
rect -27412 -10796 -27406 -10519
rect -29373 -11876 -28973 -11326
rect -27806 -11400 -27406 -10796
rect -29373 -12014 -29119 -11876
rect -28981 -12014 -28973 -11876
rect -29373 -24340 -28973 -12014
rect -28880 -11800 -27406 -11400
rect -26909 523 -26849 525
rect -26909 467 -26907 523
rect -26851 467 -26849 523
rect -28880 -15261 -28480 -11800
rect -28140 -14554 -28084 -14553
rect -28010 -14562 -27954 -14553
rect -28010 -14627 -27954 -14618
rect -28880 -15317 -28582 -15261
rect -28526 -15317 -28480 -15261
rect -28880 -17210 -28480 -15317
rect -28237 -15321 -28228 -15257
rect -28164 -15321 -28155 -15257
rect -26909 -16276 -26849 467
rect -23908 -1768 -23848 13432
rect -3844 13421 -3784 13430
rect -11066 13359 -10928 13363
rect -11071 13354 -10923 13359
rect -11071 13216 -11066 13354
rect -10928 13216 -10923 13354
rect -11071 11844 -10923 13216
rect -3842 11959 -3786 13421
rect -3842 11944 -3676 11959
rect -3842 11808 -3827 11944
rect -3691 11808 -3676 11944
rect -3488 11898 -3387 13592
rect -3842 11793 -3676 11808
rect -3494 11797 -3488 11898
rect -3387 11797 -3381 11898
rect -11071 11690 -10923 11696
rect -8185 11513 -7927 11519
rect -8185 11461 -8179 11513
rect -7933 11461 -7927 11513
rect -8185 11455 -7927 11461
rect -11364 11395 -11304 11401
rect -15364 11137 -15216 11143
rect -19254 8943 -19180 8952
rect -21437 7290 -21373 7455
rect -19254 607 -19180 8869
rect -17670 8296 -17661 8360
rect -17597 8296 -17588 8360
rect -18588 6727 -18528 6736
rect -23908 -1837 -23848 -1828
rect -26744 -7520 -26688 -7515
rect -26748 -7524 -26684 -7520
rect -26748 -7580 -26744 -7524
rect -26688 -7580 -26684 -7524
rect -26748 -14558 -26684 -7580
rect -18588 -8044 -18528 6667
rect -18293 6529 -18229 6538
rect -18293 2618 -18229 6465
rect -18293 2554 -18177 2618
rect -18241 -2878 -18177 2554
rect -17661 -2678 -17597 8296
rect -17531 605 -17457 753
rect -16331 -763 -16275 8526
rect -15364 8020 -15216 10989
rect -11364 10370 -11304 11335
rect -11364 10314 -11362 10370
rect -11306 10314 -11304 10370
rect -11364 10312 -11304 10314
rect -2262 10372 -2202 10381
rect -11362 10305 -11306 10312
rect -2262 10303 -2202 10312
rect -4707 8284 -4579 8290
rect -15364 7882 -15359 8020
rect -15221 7882 -15216 8020
rect -15364 7877 -15216 7882
rect -15155 8016 -15081 8025
rect -15155 7886 -15146 8016
rect -15090 7886 -15081 8016
rect -15155 7877 -15081 7886
rect -15359 7873 -15221 7877
rect -5316 7529 -5188 7535
rect -5959 4204 -5895 4213
rect -5959 2235 -5895 4140
rect -5568 3253 -5508 3262
rect -7731 2107 -7615 2113
rect -14886 2087 -14822 2093
rect -14886 1002 -14822 2023
rect -7731 2013 -7725 2107
rect -7621 2013 -7615 2107
rect -7725 1595 -7621 2013
rect -7725 1539 -7696 1595
rect -7640 1539 -7621 1595
rect -14886 946 -14882 1002
rect -14826 946 -14822 1002
rect -14886 942 -14822 946
rect -13792 1006 -13728 1015
rect -14882 937 -14826 942
rect -13792 -614 -13728 942
rect -9052 -222 -8924 -216
rect -9252 -465 -9124 -456
rect -13792 -670 -13788 -614
rect -13732 -670 -13728 -614
rect -13792 -674 -13728 -670
rect -11294 -610 -11230 -601
rect -13788 -679 -13732 -674
rect -16333 -772 -16273 -763
rect -11470 -772 -11414 -765
rect -16333 -841 -16273 -832
rect -11472 -774 -11412 -772
rect -11472 -830 -11470 -774
rect -11414 -830 -11412 -774
rect -11648 -900 -11584 -891
rect -11648 -1490 -11584 -964
rect -11653 -1546 -11644 -1490
rect -11588 -1546 -11579 -1490
rect -11648 -1550 -11584 -1546
rect -11472 -1661 -11412 -830
rect -11476 -1670 -11412 -1661
rect -11420 -1726 -11412 -1670
rect -11476 -1735 -11412 -1726
rect -11294 -1841 -11230 -674
rect -11294 -1897 -11292 -1841
rect -11236 -1897 -11230 -1841
rect -11294 -1909 -11230 -1897
rect -9252 -1704 -9124 -593
rect -9252 -1756 -9246 -1704
rect -9130 -1756 -9124 -1704
rect -15351 -2196 -15287 -2068
rect -17666 -2734 -17657 -2678
rect -17601 -2734 -17592 -2678
rect -17661 -2738 -17597 -2734
rect -13162 -2745 -13084 -2709
rect -18588 -8100 -18586 -8044
rect -18530 -8100 -18528 -8044
rect -18588 -8102 -18528 -8100
rect -18586 -8109 -18530 -8102
rect -26748 -14631 -26684 -14622
rect -26909 -16345 -26849 -16336
rect -28880 -17348 -28681 -17210
rect -28543 -17348 -28480 -17210
rect -28880 -23307 -28480 -17348
rect -18235 -18500 -18183 -3862
rect -16891 -4070 -16882 -4006
rect -16818 -4070 -16809 -4006
rect -16882 -11692 -16818 -4070
rect -13162 -7524 -13098 -2745
rect -13162 -7580 -13158 -7524
rect -13102 -7580 -13098 -7524
rect -13162 -7584 -13098 -7580
rect -9252 -3438 -9124 -1756
rect -9252 -3490 -9246 -3438
rect -9130 -3490 -9124 -3438
rect -9252 -4344 -9124 -3490
rect -9252 -4532 -9246 -4344
rect -9130 -4532 -9124 -4344
rect -13158 -7589 -13102 -7584
rect -16924 -11756 -16818 -11692
rect -16924 -14508 -16860 -11756
rect -16485 -11758 -16425 -11756
rect -16492 -11814 -16483 -11758
rect -16427 -11814 -16418 -11758
rect -18239 -18509 -18179 -18500
rect -18239 -18578 -18179 -18569
rect -16485 -18711 -16425 -11814
rect -16485 -18780 -16425 -18771
rect -9252 -21941 -9124 -4532
rect -9052 -1430 -8924 -350
rect -9052 -1668 -9046 -1430
rect -8930 -1668 -8924 -1430
rect -9052 -3164 -8924 -1668
rect -9052 -3402 -9046 -3164
rect -8930 -3402 -8924 -3164
rect -9052 -4600 -8924 -3402
rect -9052 -4788 -9046 -4600
rect -8930 -4788 -8924 -4600
rect -9052 -4794 -8924 -4788
rect -8852 -718 -8724 -712
rect -8852 -854 -8846 -718
rect -8730 -854 -8724 -718
rect -8852 -2244 -8724 -854
rect -8047 -1933 -7983 -1927
rect -8047 -2049 -8041 -1933
rect -7989 -2049 -7983 -1933
rect -8047 -2119 -7983 -2049
rect -8852 -2588 -8846 -2244
rect -8730 -2588 -8724 -2244
rect -8852 -3978 -8724 -2588
rect -8047 -3667 -7983 -3661
rect -8047 -3783 -8041 -3667
rect -7989 -3783 -7983 -3667
rect -8047 -3853 -7983 -3783
rect -8852 -4114 -8846 -3978
rect -8730 -4114 -8724 -3978
rect -8852 -8902 -8724 -4114
rect -7725 -6600 -7621 1539
rect -6515 -1201 -6451 -1195
rect -6515 -1317 -6509 -1201
rect -6457 -1317 -6451 -1201
rect -6515 -2796 -6451 -1317
rect -5957 -1592 -5897 2235
rect -5568 1595 -5508 3193
rect -5568 1539 -5566 1595
rect -5510 1539 -5508 1595
rect -5568 1537 -5508 1539
rect -5566 1530 -5510 1537
rect -5316 -222 -5188 7401
rect -4906 7299 -4849 7305
rect -5316 -356 -5188 -350
rect -4907 7242 -4906 7294
rect -4849 7242 -4779 7294
rect -4907 5350 -4779 7242
rect -4907 5254 -4887 5350
rect -4791 5254 -4779 5350
rect -4907 4523 -4779 5254
rect -4907 4427 -4891 4523
rect -4795 4427 -4779 4523
rect -4907 3699 -4779 4427
rect -4907 3540 -4899 3699
rect -4785 3540 -4779 3699
rect -4907 2363 -4779 3540
rect -4907 2287 -4898 2363
rect -4791 2287 -4779 2363
rect -4907 1625 -4779 2287
rect -4907 1529 -4895 1625
rect -4799 1529 -4779 1625
rect -4907 -466 -4779 1529
rect -4907 -600 -4779 -594
rect -4707 6743 -4579 8156
rect -2260 7795 -2204 10303
rect -2266 7739 -2260 7795
rect -2204 7739 -2198 7795
rect -4707 4806 -4579 6615
rect -4707 4710 -4684 4806
rect -4588 4710 -4579 4806
rect -4707 3979 -4579 4710
rect -4707 3883 -4688 3979
rect -4592 3883 -4579 3979
rect -4707 3054 -4579 3883
rect -4707 2897 -4698 3054
rect -4588 2897 -4579 3054
rect -4707 1824 -4579 2897
rect -4707 1740 -4699 1824
rect -4587 1740 -4579 1824
rect -4707 1081 -4579 1740
rect -4480 7036 -4420 7045
rect -3790 7042 -3734 7043
rect -4480 5027 -4420 6976
rect -3798 7036 -3726 7042
rect -3798 6976 -3792 7036
rect -3732 6976 -3726 7036
rect -3798 6970 -3726 6976
rect -3790 6969 -3734 6970
rect -2598 5082 -2532 5091
rect -4306 5035 -4250 5036
rect -4480 4971 -4478 5027
rect -4422 4971 -4420 5027
rect -4480 1300 -4420 4971
rect -4314 5029 -4242 5035
rect -4314 4969 -4308 5029
rect -4248 4969 -4242 5029
rect -4314 4963 -4242 4969
rect -4306 4962 -4250 4963
rect -2598 4859 -2590 5082
rect -2538 5002 -2532 5082
rect -2538 4950 -2438 5002
rect -2538 4859 -2532 4950
rect -2598 4853 -2532 4859
rect -2598 4255 -2532 4264
rect -4306 4208 -4250 4209
rect -4314 4202 -4242 4208
rect -4314 4142 -4308 4202
rect -4248 4142 -4242 4202
rect -4314 4136 -4242 4142
rect -4306 4135 -4250 4136
rect -2598 4032 -2590 4255
rect -2538 4175 -2532 4255
rect -2538 4123 -2438 4175
rect -2538 4032 -2532 4123
rect -2598 4026 -2532 4032
rect -4060 3261 -4004 3360
rect -4062 3252 -4004 3261
rect -4006 3196 -4004 3252
rect -4062 3187 -4004 3196
rect -4060 3129 -4004 3187
rect -3651 2836 -3595 2843
rect -3653 2834 -3593 2836
rect -3653 2778 -3651 2834
rect -3595 2778 -3593 2834
rect -3653 2553 -3593 2778
rect -4117 2551 -4057 2553
rect -4124 2495 -4115 2551
rect -4059 2495 -4050 2551
rect -4117 2052 -4057 2495
rect -3653 2484 -3593 2493
rect -2599 2153 -2532 2165
rect -2599 2044 -2594 2153
rect -4117 1986 -4057 1992
rect -2600 1988 -2594 2044
rect -2599 1898 -2594 1988
rect -2538 2044 -2532 2153
rect -2538 1988 -2411 2044
rect -2538 1898 -2532 1988
rect -2599 1886 -2532 1898
rect -2138 1334 -2072 1343
rect -4300 1303 -4244 1307
rect -4480 1231 -4420 1240
rect -4333 1298 -4176 1303
rect -4333 1297 -4300 1298
rect -4244 1297 -4176 1298
rect -4333 1245 -4327 1297
rect -4184 1245 -4176 1297
rect -4333 1242 -4300 1245
rect -4244 1242 -4176 1245
rect -4333 1239 -4176 1242
rect -4300 1233 -4223 1239
rect -4279 1160 -4223 1233
rect -2138 1142 -2130 1334
rect -2078 1269 -2072 1334
rect -2078 1213 -1997 1269
rect -2078 1142 -2072 1213
rect -2138 1134 -2072 1142
rect -4707 985 -4695 1081
rect -4599 985 -4579 1081
rect -4707 -728 -4579 985
rect -4707 -862 -4579 -856
rect -6101 -1652 -5897 -1592
rect -4403 -1201 -4339 -1195
rect -4403 -1317 -4397 -1201
rect -4345 -1317 -4339 -1201
rect -6101 -1845 -6041 -1652
rect -6101 -1914 -6041 -1905
rect -5935 -1933 -5871 -1927
rect -5935 -2049 -5929 -1933
rect -5877 -2049 -5871 -1933
rect -5935 -2119 -5871 -2049
rect -4403 -2767 -4339 -1317
rect -4279 -2589 -4223 954
rect -2291 -1201 -2227 -1195
rect -2291 -1317 -2285 -1201
rect -2233 -1317 -2227 -1201
rect -3823 -1933 -3759 -1927
rect -3823 -2049 -3817 -1933
rect -3765 -2049 -3759 -1933
rect -3823 -2119 -3759 -2049
rect -4279 -2645 -4061 -2589
rect -6515 -2860 -6341 -2796
rect -4403 -2831 -4223 -2767
rect -7725 -6713 -7621 -6704
rect -6515 -2935 -6451 -2929
rect -6515 -3051 -6509 -2935
rect -6457 -3051 -6451 -2935
rect -6515 -7297 -6451 -3051
rect -6405 -7158 -6341 -2860
rect -4403 -2935 -4339 -2929
rect -4403 -3051 -4397 -2935
rect -4345 -3051 -4339 -2935
rect -4403 -3489 -4339 -3051
rect -4287 -3470 -4223 -2831
rect -4117 -3345 -4061 -2645
rect -2291 -2745 -2227 -1317
rect -179 -1201 -115 -1195
rect -179 -1317 -173 -1201
rect -121 -1317 -115 -1201
rect -1711 -1933 -1647 -1927
rect -1711 -2049 -1705 -1933
rect -1653 -2049 -1647 -1933
rect -1711 -2119 -1647 -2049
rect -179 -2724 -115 -1317
rect 1933 -1201 1997 -1195
rect 1933 -1317 1939 -1201
rect 1991 -1317 1997 -1201
rect 401 -1933 465 -1927
rect 401 -2049 407 -1933
rect 459 -2049 465 -1933
rect 401 -2246 465 -2049
rect 401 -2316 465 -2310
rect -2291 -2809 -2111 -2745
rect -179 -2788 44 -2724
rect -2291 -2935 -2227 -2929
rect -2291 -3051 -2285 -2935
rect -2233 -3051 -2227 -2935
rect -4119 -3354 -4059 -3345
rect -4119 -3423 -4059 -3414
rect -4403 -3529 -4338 -3489
rect -4287 -3519 -4222 -3470
rect -5935 -3667 -5871 -3661
rect -5935 -3783 -5929 -3667
rect -5877 -3783 -5871 -3667
rect -4402 -3702 -4338 -3529
rect -4286 -3569 -4222 -3519
rect -4286 -3625 -4282 -3569
rect -4226 -3625 -4222 -3569
rect -4286 -3629 -4222 -3625
rect -2618 -3565 -2554 -3556
rect -4282 -3634 -4226 -3629
rect -4402 -3758 -4398 -3702
rect -4342 -3758 -4338 -3702
rect -4402 -3762 -4338 -3758
rect -3823 -3667 -3759 -3661
rect -4398 -3767 -4342 -3762
rect -5935 -3853 -5871 -3783
rect -3823 -3783 -3817 -3667
rect -3765 -3783 -3759 -3667
rect -3823 -3853 -3759 -3783
rect -3146 -3698 -3082 -3689
rect -3666 -7152 -3610 -7147
rect -6405 -7231 -6341 -7222
rect -3670 -7156 -3606 -7152
rect -3670 -7212 -3666 -7156
rect -3610 -7212 -3606 -7156
rect -6515 -7370 -6451 -7361
rect -4212 -7302 -4156 -7293
rect -4212 -7367 -4156 -7358
rect -3670 -7371 -3606 -7212
rect -3146 -7382 -3082 -3762
rect -2618 -7374 -2554 -3629
rect -2291 -4510 -2227 -3051
rect -2175 -4344 -2111 -2809
rect -179 -2935 -115 -2929
rect -179 -3051 -173 -2935
rect -121 -3051 -115 -2935
rect -1711 -3667 -1647 -3661
rect -1711 -3783 -1705 -3667
rect -1653 -3783 -1647 -3667
rect -1711 -3853 -1647 -3783
rect -2175 -4417 -2111 -4408
rect -1533 -4344 -1469 -4335
rect -2291 -4583 -2227 -4574
rect -2083 -4511 -2019 -4502
rect -2083 -7374 -2019 -4575
rect -1533 -7374 -1469 -4408
rect -1003 -4826 -934 -4817
rect -1003 -7367 -934 -4895
rect -179 -4830 -115 -3051
rect -179 -4889 -173 -4830
rect -117 -4889 -115 -4830
rect -179 -4899 -115 -4889
rect -20 -4872 44 -2788
rect 1933 -2782 1997 -1317
rect 4045 -1201 4109 -1195
rect 4045 -1317 4051 -1201
rect 4103 -1317 4109 -1201
rect 2513 -1933 2577 -1927
rect 2513 -2049 2519 -1933
rect 2571 -2049 2577 -1933
rect 2513 -2248 2577 -2049
rect 2513 -2318 2577 -2312
rect 4045 -2778 4109 -1317
rect 6157 -1201 6221 -1195
rect 6157 -1317 6163 -1201
rect 6215 -1317 6221 -1201
rect 4625 -1933 4689 -1927
rect 4625 -2049 4631 -1933
rect 4683 -2049 4689 -1933
rect 4625 -2242 4689 -2049
rect 4625 -2312 4689 -2306
rect 6157 -2771 6221 -1317
rect 8269 -1201 8333 -1195
rect 8269 -1317 8275 -1201
rect 8327 -1317 8333 -1201
rect 6737 -1933 6801 -1927
rect 6737 -2049 6743 -1933
rect 6795 -2049 6801 -1933
rect 6737 -2248 6801 -2049
rect 6737 -2318 6801 -2312
rect 8269 -2742 8333 -1317
rect 10381 -1201 10445 -1195
rect 10381 -1317 10387 -1201
rect 10439 -1317 10445 -1201
rect 10381 -1486 10445 -1317
rect 10381 -1559 10445 -1550
rect 10636 -1324 10696 -1318
rect 10636 -1670 10696 -1384
rect 10629 -1726 10638 -1670
rect 10694 -1726 10703 -1670
rect 10636 -1728 10696 -1726
rect 11174 -1837 11250 -1831
rect 11174 -1901 11180 -1837
rect 11244 -1901 11250 -1837
rect 11174 -1907 11250 -1901
rect 8849 -1933 8913 -1927
rect 8849 -2049 8855 -1933
rect 8907 -2049 8913 -1933
rect 8849 -2119 8913 -2049
rect 1933 -2846 2149 -2782
rect 4045 -2842 4247 -2778
rect 6157 -2835 6367 -2771
rect 8269 -2806 8480 -2742
rect 1933 -2935 1997 -2929
rect 1933 -3051 1939 -2935
rect 1991 -3051 1997 -2935
rect 401 -3667 465 -3661
rect 401 -3783 407 -3667
rect 459 -3783 465 -3667
rect 401 -3970 465 -3783
rect 1076 -3859 1132 -3854
rect 1933 -3859 1997 -3051
rect 401 -4040 465 -4034
rect 1072 -3863 1136 -3859
rect 1072 -3919 1076 -3863
rect 1132 -3919 1136 -3863
rect -20 -4899 47 -4872
rect -479 -5097 -470 -5033
rect -406 -5097 -397 -5033
rect -17 -5037 47 -4899
rect -17 -5093 -13 -5037
rect 43 -5093 47 -5037
rect -17 -5097 47 -5093
rect -470 -7382 -406 -5097
rect -13 -5102 43 -5097
rect 72 -5202 136 -5193
rect 1072 -5206 1136 -3919
rect 1933 -3932 1997 -3923
rect 1597 -3997 1653 -3992
rect 2085 -3997 2149 -2846
rect 4045 -2935 4109 -2929
rect 4045 -3051 4051 -2935
rect 4103 -3051 4109 -2935
rect 1593 -4001 1657 -3997
rect 1593 -4057 1597 -4001
rect 1653 -4057 1657 -4001
rect 1593 -4872 1657 -4057
rect 2513 -3667 2577 -3661
rect 2513 -3783 2519 -3667
rect 2571 -3783 2577 -3667
rect 2513 -3984 2577 -3783
rect 2513 -4054 2577 -4048
rect 2085 -4070 2149 -4061
rect 2140 -4157 2196 -4152
rect 4045 -4157 4109 -3051
rect 2136 -4161 2200 -4157
rect 2136 -4217 2140 -4161
rect 2196 -4217 2200 -4161
rect 2136 -4830 2200 -4217
rect 4045 -4230 4109 -4221
rect 2669 -4311 2725 -4306
rect 4183 -4311 4247 -2842
rect 6157 -2935 6221 -2929
rect 6157 -3051 6163 -2935
rect 6215 -3051 6221 -2935
rect 4625 -3667 4689 -3661
rect 4625 -3783 4631 -3667
rect 4683 -3783 4689 -3667
rect 4625 -3984 4689 -3783
rect 4625 -4054 4689 -4048
rect 2665 -4315 2729 -4311
rect 2665 -4371 2669 -4315
rect 2725 -4371 2729 -4315
rect 1593 -4899 1658 -4872
rect 2136 -4899 2201 -4830
rect 1072 -5262 1076 -5206
rect 1132 -5262 1136 -5206
rect 1072 -5266 1136 -5262
rect 72 -7374 136 -5266
rect 1076 -5271 1132 -5266
rect 593 -5367 657 -5358
rect 1594 -5371 1658 -4899
rect 1594 -5427 1598 -5371
rect 1654 -5427 1658 -5371
rect 1594 -5431 1658 -5427
rect 593 -7367 657 -5431
rect 1598 -5436 1654 -5431
rect 1136 -5543 1200 -5534
rect 2137 -5547 2201 -4899
rect 2137 -5603 2141 -5547
rect 2197 -5603 2201 -5547
rect 2137 -5607 2201 -5603
rect 1136 -7332 1200 -5607
rect 2141 -5612 2197 -5607
rect 1665 -5732 1729 -5723
rect 2665 -5736 2729 -4371
rect 4183 -4384 4247 -4375
rect 3205 -4458 3261 -4453
rect 6157 -4458 6221 -3051
rect 3201 -4462 3265 -4458
rect 3201 -4518 3205 -4462
rect 3261 -4518 3265 -4462
rect 3201 -4802 3265 -4518
rect 6157 -4531 6221 -4522
rect 3747 -4612 3803 -4607
rect 6303 -4612 6367 -2835
rect 8269 -2935 8333 -2929
rect 8269 -3051 8275 -2935
rect 8327 -3051 8333 -2935
rect 6737 -3667 6801 -3661
rect 6737 -3783 6743 -3667
rect 6795 -3783 6801 -3667
rect 6737 -3980 6793 -3783
rect 6737 -4042 6793 -4036
rect 3743 -4616 3807 -4612
rect 3743 -4672 3747 -4616
rect 3803 -4672 3807 -4616
rect 3743 -4791 3807 -4672
rect 6303 -4685 6367 -4676
rect 3201 -4899 3267 -4802
rect 3743 -4899 3810 -4791
rect 4275 -4796 4331 -4791
rect 8269 -4796 8333 -3051
rect 4271 -4800 4335 -4796
rect 4271 -4856 4275 -4800
rect 4331 -4856 4335 -4800
rect 4271 -4861 4335 -4856
rect 4271 -4899 4336 -4861
rect 8269 -4869 8333 -4860
rect 8416 -4850 8480 -2806
rect 10381 -2935 10445 -2929
rect 10381 -3051 10387 -2935
rect 10439 -3051 10445 -2935
rect 8849 -3667 8913 -3661
rect 8849 -3783 8855 -3667
rect 8907 -3783 8913 -3667
rect 8849 -3853 8913 -3783
rect 10381 -4841 10445 -3051
rect 10636 -3056 10700 -3050
rect 10636 -3688 10700 -3120
rect 11199 -3354 11255 -3347
rect 11197 -3356 11257 -3354
rect 11197 -3412 11199 -3356
rect 11255 -3412 11257 -3356
rect 11197 -3588 11257 -3412
rect 11197 -3654 11257 -3648
rect 10636 -3744 10640 -3688
rect 10696 -3744 10700 -3688
rect 10636 -3748 10700 -3744
rect 10640 -3753 10696 -3748
rect 8416 -4899 8481 -4850
rect 2665 -5792 2669 -5736
rect 2725 -5792 2729 -5736
rect 2665 -5796 2729 -5792
rect 1665 -7375 1729 -5796
rect 2669 -5801 2725 -5796
rect 2201 -5925 2265 -5916
rect 3203 -5929 3267 -4899
rect 3203 -5985 3207 -5929
rect 3263 -5985 3267 -5929
rect 3203 -5989 3267 -5985
rect 2201 -7382 2265 -5989
rect 3207 -5994 3263 -5989
rect 2743 -6094 2807 -6085
rect 3746 -6098 3810 -4899
rect 3746 -6154 3750 -6098
rect 3806 -6154 3810 -6098
rect 3746 -6158 3810 -6154
rect 2743 -7390 2807 -6158
rect 3750 -6163 3806 -6158
rect 3271 -6270 3335 -6261
rect 4272 -6274 4336 -4899
rect 4272 -6330 4276 -6274
rect 4332 -6330 4336 -6274
rect 4272 -6334 4336 -6330
rect 4424 -4984 4488 -4975
rect 8417 -4988 8481 -4899
rect 8417 -5044 8421 -4988
rect 8477 -5044 8481 -4988
rect 8417 -5048 8481 -5044
rect 10380 -4899 10445 -4841
rect 3271 -7368 3335 -6334
rect 4276 -6339 4332 -6334
rect 3801 -6421 3865 -6412
rect 4424 -6425 4488 -5048
rect 8421 -5053 8477 -5048
rect 4424 -6481 4428 -6425
rect 4484 -6481 4488 -6425
rect 4424 -6485 4488 -6481
rect 4571 -5188 4635 -5179
rect 10380 -5192 10444 -4899
rect 10380 -5248 10384 -5192
rect 10440 -5248 10444 -5192
rect 10380 -5252 10444 -5248
rect 3801 -7368 3865 -6485
rect 4428 -6490 4484 -6485
rect -5084 -7520 -5028 -7515
rect -5088 -7524 -5024 -7520
rect -5088 -7580 -5084 -7524
rect -5028 -7580 -5024 -7524
rect -5088 -8780 -5024 -7580
rect 4571 -7524 4635 -5252
rect 10384 -5257 10440 -5252
rect 4571 -7580 4575 -7524
rect 4631 -7580 4635 -7524
rect 4571 -7584 4635 -7580
rect 4575 -7589 4631 -7584
rect -4390 -8042 -4330 -8033
rect -4390 -8904 -4330 -8102
rect -4390 -8960 -4388 -8904
rect -4332 -8960 -4330 -8904
rect -4390 -8962 -4330 -8960
rect -4388 -8969 -4332 -8962
rect -10867 -21963 -10766 -21957
rect -10867 -22052 -10861 -21963
rect -10772 -22052 -10766 -21963
rect -10867 -22058 -10766 -22052
rect -9261 -22069 -9252 -21941
rect -9124 -22069 -9115 -21941
rect -10877 -22354 -10817 -22202
rect -14211 -22492 -14151 -22364
rect -10549 -22947 -10409 -22941
rect -8852 -22947 -8724 -9030
rect -7484 -9963 -7380 -9815
rect -5082 -10830 -4381 -10824
rect -5082 -11018 -5076 -10830
rect -4893 -11018 -4575 -10830
rect -4387 -11018 -4381 -10830
rect -5082 -11024 -4381 -11018
rect 427 -11747 483 -9708
rect 425 -11756 485 -11747
rect 425 -11825 485 -11816
rect -10549 -23075 -10543 -22947
rect -10415 -23075 -10409 -22947
rect -8861 -23075 -8852 -22947
rect -8724 -23075 -8715 -22947
rect -10549 -23081 -10409 -23075
rect -28880 -23445 -28677 -23307
rect -28539 -23445 -28480 -23307
rect -28880 -24350 -28480 -23445
<< via2 >>
rect -27525 13598 -27434 13689
rect -3488 13592 -3387 13695
rect -28900 13216 -28762 13354
rect -27929 13217 -27868 13353
rect -23906 13432 -23850 13488
rect -27042 8300 -26986 8356
rect -27478 7883 -27412 8019
rect -27478 1786 -27412 1922
rect -29119 -12014 -28981 -11876
rect -26907 467 -26851 523
rect -28010 -14618 -27954 -14562
rect -28582 -15317 -28526 -15261
rect -28228 -15321 -28164 -15257
rect -3844 13430 -3784 13490
rect -11066 13216 -10928 13354
rect -19254 8869 -19180 8943
rect -17661 8296 -17597 8360
rect -18588 6667 -18528 6727
rect -23908 -1828 -23848 -1768
rect -26744 -7580 -26688 -7524
rect -18293 6465 -18229 6529
rect -11362 10314 -11306 10370
rect -2262 10312 -2202 10372
rect -15359 7882 -15221 8020
rect -15146 7886 -15090 8016
rect -5959 4140 -5895 4204
rect -5568 3193 -5508 3253
rect -7696 1539 -7640 1595
rect -14882 946 -14826 1002
rect -13792 942 -13728 1006
rect -13788 -670 -13732 -614
rect -11294 -674 -11230 -610
rect -16333 -832 -16273 -772
rect -11470 -830 -11414 -774
rect -11648 -964 -11584 -900
rect -11644 -1546 -11588 -1490
rect -11476 -1726 -11420 -1670
rect -11292 -1897 -11236 -1841
rect -17657 -2734 -17601 -2678
rect -18586 -8100 -18530 -8044
rect -26748 -14622 -26684 -14558
rect -26909 -16336 -26849 -16276
rect -28681 -17348 -28543 -17210
rect -16882 -4070 -16818 -4006
rect -13158 -7580 -13102 -7524
rect -16483 -11814 -16427 -11758
rect -18239 -18569 -18179 -18509
rect -16485 -18771 -16425 -18711
rect -5566 1539 -5510 1595
rect -4480 6976 -4420 7036
rect -3790 6978 -3734 7034
rect -4478 4971 -4422 5027
rect -4306 4971 -4250 5027
rect -4306 4144 -4250 4200
rect -4062 3196 -4006 3252
rect -3651 2778 -3595 2834
rect -4115 2495 -4059 2551
rect -3653 2493 -3593 2553
rect -4480 1240 -4420 1300
rect -4300 1297 -4244 1298
rect -4300 1245 -4244 1297
rect -4300 1242 -4244 1245
rect -6101 -1905 -6041 -1845
rect -7725 -6704 -7621 -6600
rect -4119 -3414 -4059 -3354
rect -4282 -3625 -4226 -3569
rect -2618 -3629 -2554 -3565
rect -4398 -3758 -4342 -3702
rect -3146 -3762 -3082 -3698
rect -6405 -7222 -6341 -7158
rect -3666 -7212 -3610 -7156
rect -6515 -7361 -6451 -7297
rect -4212 -7358 -4156 -7302
rect -2175 -4408 -2111 -4344
rect -1533 -4408 -1469 -4344
rect -2291 -4574 -2227 -4510
rect -2083 -4575 -2019 -4511
rect -1003 -4895 -934 -4826
rect -173 -4889 -117 -4830
rect 10381 -1550 10445 -1486
rect 10638 -1726 10694 -1670
rect 11184 -1897 11240 -1841
rect 1076 -3919 1132 -3863
rect -470 -5097 -406 -5033
rect -13 -5093 43 -5037
rect 72 -5266 136 -5202
rect 1933 -3923 1997 -3859
rect 1597 -4057 1653 -4001
rect 2085 -4061 2149 -3997
rect 2140 -4217 2196 -4161
rect 4045 -4221 4109 -4157
rect 2669 -4371 2725 -4315
rect 1076 -5262 1132 -5206
rect 593 -5431 657 -5367
rect 1598 -5427 1654 -5371
rect 1136 -5607 1200 -5543
rect 2141 -5603 2197 -5547
rect 1665 -5796 1729 -5732
rect 4183 -4375 4247 -4311
rect 3205 -4518 3261 -4462
rect 6157 -4522 6221 -4458
rect 3747 -4672 3803 -4616
rect 6303 -4676 6367 -4612
rect 4275 -4856 4331 -4800
rect 8269 -4860 8333 -4796
rect 11199 -3412 11255 -3356
rect 10640 -3744 10696 -3688
rect 2669 -5792 2725 -5736
rect 2201 -5989 2265 -5925
rect 3207 -5985 3263 -5929
rect 2743 -6158 2807 -6094
rect 3750 -6154 3806 -6098
rect 3271 -6334 3335 -6270
rect 4276 -6330 4332 -6274
rect 4424 -5048 4488 -4984
rect 8421 -5044 8477 -4988
rect 3801 -6485 3865 -6421
rect 4428 -6481 4484 -6425
rect 4571 -5252 4635 -5188
rect 10384 -5248 10440 -5192
rect -5084 -7580 -5028 -7524
rect 4575 -7580 4631 -7524
rect -4390 -8102 -4330 -8042
rect -8852 -9030 -8724 -8902
rect -4388 -8960 -4332 -8904
rect -10856 -22047 -10777 -21968
rect -9252 -22069 -9124 -21941
rect 425 -11816 485 -11756
rect -10538 -23070 -10420 -22952
rect -8852 -23075 -8724 -22947
rect -28677 -23445 -28539 -23307
<< metal3 >>
rect -3493 13695 -3382 13700
rect -3493 13694 -3488 13695
rect -27530 13689 -3488 13694
rect -27530 13598 -27525 13689
rect -27434 13598 -3488 13689
rect -27530 13593 -3488 13598
rect -3493 13592 -3488 13593
rect -3387 13592 -3382 13695
rect -3493 13587 -3382 13592
rect -23911 13490 -23845 13493
rect -3849 13490 -3779 13495
rect -23911 13488 -3844 13490
rect -23911 13432 -23906 13488
rect -23850 13432 -3844 13488
rect -23911 13430 -3844 13432
rect -3784 13430 -3779 13490
rect -23911 13427 -23845 13430
rect -3849 13425 -3779 13430
rect -28905 13354 -27136 13359
rect -28905 13216 -28900 13354
rect -28762 13353 -27136 13354
rect -28762 13217 -27929 13353
rect -27868 13217 -27136 13353
rect -28762 13216 -27136 13217
rect -28905 13211 -27136 13216
rect -16022 13354 -10923 13359
rect -16022 13216 -11066 13354
rect -10928 13216 -10923 13354
rect -16022 13211 -10923 13216
rect -11367 10372 -11301 10375
rect -2267 10372 -2197 10377
rect -11367 10370 -2262 10372
rect -11367 10314 -11362 10370
rect -11306 10314 -2262 10370
rect -11367 10312 -2262 10314
rect -2202 10312 -2197 10372
rect -11367 10309 -11301 10312
rect -2267 10307 -2197 10312
rect -19259 8943 -19175 8948
rect -27181 8869 -19254 8943
rect -19180 8869 -19175 8943
rect -19259 8864 -19175 8869
rect -27047 8360 -26981 8361
rect -17666 8360 -17592 8365
rect -27047 8356 -17661 8360
rect -27047 8300 -27042 8356
rect -26986 8300 -17661 8356
rect -27047 8296 -17661 8300
rect -17597 8296 -17592 8360
rect -27047 8295 -26981 8296
rect -17666 8291 -17592 8296
rect -27484 8019 -27166 8025
rect -27484 7883 -27478 8019
rect -27412 7883 -27166 8019
rect -27484 7877 -27166 7883
rect -15503 8020 -15081 8025
rect -15503 7882 -15359 8020
rect -15221 8016 -15081 8020
rect -15221 7886 -15146 8016
rect -15090 7886 -15081 8016
rect -15221 7882 -15081 7886
rect -15503 7877 -15081 7882
rect -4485 7036 -4415 7041
rect -3795 7036 -3729 7039
rect -4485 6976 -4480 7036
rect -4420 7034 -3729 7036
rect -4420 6978 -3790 7034
rect -3734 6978 -3729 7034
rect -4420 6976 -3729 6978
rect -4485 6971 -4415 6976
rect -3795 6973 -3729 6976
rect -18593 6727 -18523 6732
rect -18593 6667 -18588 6727
rect -18528 6667 -18523 6727
rect -18593 6662 -18523 6667
rect -18298 6529 -18224 6534
rect -18298 6465 -18293 6529
rect -18229 6465 -18224 6529
rect -18298 6460 -18224 6465
rect -4483 5029 -4417 5032
rect -4311 5029 -4245 5032
rect -4483 5027 -4245 5029
rect -4483 4971 -4478 5027
rect -4422 4971 -4306 5027
rect -4250 4971 -4245 5027
rect -4483 4969 -4245 4971
rect -4483 4966 -4417 4969
rect -4311 4966 -4245 4969
rect -5964 4204 -5890 4209
rect -5964 4140 -5959 4204
rect -5895 4202 -4919 4204
rect -4311 4202 -4245 4205
rect -5895 4200 -4245 4202
rect -5895 4144 -4306 4200
rect -4250 4144 -4245 4200
rect -5895 4142 -4245 4144
rect -5895 4140 -4919 4142
rect -5964 4135 -5890 4140
rect -4311 4139 -4245 4142
rect -5573 3253 -5503 3258
rect -4067 3254 -4001 3257
rect -5057 3253 -4001 3254
rect -5573 3193 -5568 3253
rect -5508 3252 -4001 3253
rect -5508 3196 -4062 3252
rect -4006 3196 -4001 3252
rect -5508 3194 -4001 3196
rect -5508 3193 -4947 3194
rect -5573 3188 -5503 3193
rect -4067 3191 -4001 3194
rect -3656 2836 -3590 2839
rect -3656 2834 -3395 2836
rect -3656 2778 -3651 2834
rect -3595 2778 -3395 2834
rect -3656 2776 -3395 2778
rect -3656 2773 -3590 2776
rect -4120 2553 -4054 2556
rect -3658 2553 -3588 2558
rect -4120 2551 -3653 2553
rect -4120 2495 -4115 2551
rect -4059 2495 -3653 2551
rect -4120 2493 -3653 2495
rect -3593 2493 -3588 2553
rect -4120 2490 -4054 2493
rect -3658 2488 -3588 2493
rect -27484 1922 -26420 1928
rect -27484 1786 -27478 1922
rect -27412 1786 -26420 1922
rect -27484 1780 -26420 1786
rect -7701 1597 -7635 1600
rect -5571 1597 -5505 1600
rect -7701 1595 -5505 1597
rect -7701 1539 -7696 1595
rect -7640 1539 -5566 1595
rect -5510 1539 -5505 1595
rect -7701 1537 -5505 1539
rect -7701 1534 -7635 1537
rect -5571 1534 -5505 1537
rect -4485 1300 -4415 1305
rect -4305 1300 -4239 1303
rect -4485 1240 -4480 1300
rect -4420 1298 -4239 1300
rect -4420 1242 -4300 1298
rect -4244 1242 -4239 1298
rect -4420 1240 -4239 1242
rect -4485 1235 -4415 1240
rect -4305 1237 -4239 1240
rect -14887 1006 -14821 1007
rect -13797 1006 -13723 1011
rect -14887 1002 -13792 1006
rect -14887 946 -14882 1002
rect -14826 946 -13792 1002
rect -14887 942 -13792 946
rect -13728 942 -13723 1006
rect -14887 941 -14821 942
rect -13797 937 -13723 942
rect -17297 655 -14099 715
rect -26912 525 -26846 528
rect -17297 525 -17237 655
rect -26912 523 -17237 525
rect -26912 467 -26907 523
rect -26851 467 -17237 523
rect -26912 465 -17237 467
rect -26912 462 -26846 465
rect -13793 -610 -13727 -609
rect -11299 -610 -11225 -605
rect -13793 -614 -11294 -610
rect -13793 -670 -13788 -614
rect -13732 -670 -11294 -614
rect -13793 -674 -11294 -670
rect -11230 -674 -11225 -610
rect -13793 -675 -13727 -674
rect -11299 -679 -11225 -674
rect -16338 -772 -16268 -767
rect -11475 -772 -11409 -769
rect -16338 -832 -16333 -772
rect -16273 -774 -11409 -772
rect -16273 -830 -11470 -774
rect -11414 -830 -11409 -774
rect -16273 -832 -11409 -830
rect -16338 -837 -16268 -832
rect -11475 -835 -11409 -832
rect -11653 -900 -11579 -895
rect -11771 -964 -11648 -900
rect -11584 -964 -11579 -900
rect -11653 -969 -11579 -964
rect -11649 -1486 -11583 -1485
rect 10376 -1486 10450 -1481
rect -11649 -1490 10381 -1486
rect -11649 -1546 -11644 -1490
rect -11588 -1546 10381 -1490
rect -11649 -1550 10381 -1546
rect 10445 -1550 10450 -1486
rect -11649 -1551 -11583 -1550
rect 10376 -1555 10450 -1550
rect -11481 -1668 -11415 -1665
rect 10633 -1668 10699 -1665
rect -11481 -1670 10699 -1668
rect -11481 -1726 -11476 -1670
rect -11420 -1726 10638 -1670
rect 10694 -1726 10699 -1670
rect -11481 -1728 10699 -1726
rect -11481 -1731 -11415 -1728
rect 10633 -1731 10699 -1728
rect -23913 -1768 -23843 -1763
rect -23913 -1828 -23908 -1768
rect -23848 -1828 -23843 -1768
rect -23913 -1833 -23843 -1828
rect -11297 -1837 -11231 -1836
rect 11174 -1837 11250 -1831
rect -11297 -1841 11250 -1837
rect -11297 -1897 -11292 -1841
rect -11236 -1845 11184 -1841
rect -11236 -1897 -6101 -1845
rect -11297 -1901 -6101 -1897
rect -11297 -1902 -11231 -1901
rect -6106 -1905 -6101 -1901
rect -6041 -1897 11184 -1845
rect 11240 -1897 11250 -1841
rect -6041 -1901 11250 -1897
rect -6041 -1905 -6036 -1901
rect -6106 -1910 -6036 -1905
rect 11174 -1907 11250 -1901
rect -17662 -2674 -17596 -2673
rect -17662 -2678 -15348 -2674
rect -17662 -2734 -17657 -2678
rect -17601 -2734 -15348 -2678
rect -17662 -2738 -15348 -2734
rect -17662 -2739 -17596 -2738
rect -15414 -2793 -15348 -2738
rect -15414 -2858 -15412 -2793
rect -4124 -3354 -4054 -3349
rect 11194 -3354 11260 -3351
rect -4124 -3414 -4119 -3354
rect -4059 -3356 11260 -3354
rect -4059 -3412 11199 -3356
rect 11255 -3412 11260 -3356
rect -4059 -3414 11260 -3412
rect -4124 -3419 -4054 -3414
rect 11194 -3417 11260 -3414
rect -4287 -3565 -4221 -3564
rect -2623 -3565 -2549 -3560
rect -4287 -3569 -2618 -3565
rect -4287 -3625 -4282 -3569
rect -4226 -3625 -2618 -3569
rect -4287 -3629 -2618 -3625
rect -2554 -3629 -2549 -3565
rect -4287 -3630 -4221 -3629
rect -2623 -3634 -2549 -3629
rect 10635 -3684 10701 -3683
rect 732 -3688 10701 -3684
rect -4403 -3698 -4337 -3697
rect -3151 -3698 -3077 -3693
rect -4403 -3702 -3146 -3698
rect -4403 -3758 -4398 -3702
rect -4342 -3758 -3146 -3702
rect -4403 -3762 -3146 -3758
rect -3082 -3762 -3077 -3698
rect -4403 -3763 -4337 -3762
rect -3151 -3767 -3077 -3762
rect 732 -3744 10640 -3688
rect 10696 -3744 10701 -3688
rect 732 -3748 10701 -3744
rect -16887 -4006 -16813 -4001
rect 732 -4006 796 -3748
rect 10635 -3749 10701 -3748
rect 1071 -3859 1137 -3858
rect 1928 -3859 2002 -3854
rect 1071 -3863 1933 -3859
rect 1071 -3919 1076 -3863
rect 1132 -3919 1933 -3863
rect 1071 -3923 1933 -3919
rect 1997 -3923 2002 -3859
rect 1071 -3924 1137 -3923
rect 1928 -3928 2002 -3923
rect -16887 -4070 -16882 -4006
rect -16818 -4070 796 -4006
rect 1592 -3997 1658 -3996
rect 2080 -3997 2154 -3992
rect 1592 -4001 2085 -3997
rect 1592 -4057 1597 -4001
rect 1653 -4057 2085 -4001
rect 1592 -4061 2085 -4057
rect 2149 -4061 2154 -3997
rect 1592 -4062 1658 -4061
rect 2080 -4066 2154 -4061
rect -16887 -4075 -16813 -4070
rect 2135 -4157 2201 -4156
rect 4040 -4157 4114 -4152
rect 2135 -4161 4045 -4157
rect 2135 -4217 2140 -4161
rect 2196 -4217 4045 -4161
rect 2135 -4221 4045 -4217
rect 4109 -4221 4114 -4157
rect 2135 -4222 2201 -4221
rect 4040 -4226 4114 -4221
rect 2664 -4311 2730 -4310
rect 4178 -4311 4252 -4306
rect 2664 -4315 4183 -4311
rect -2180 -4344 -2106 -4339
rect -1538 -4344 -1464 -4339
rect -2180 -4408 -2175 -4344
rect -2111 -4408 -1533 -4344
rect -1469 -4408 -1464 -4344
rect 2664 -4371 2669 -4315
rect 2725 -4371 4183 -4315
rect 2664 -4375 4183 -4371
rect 4247 -4375 4252 -4311
rect 2664 -4376 2730 -4375
rect 4178 -4380 4252 -4375
rect -2180 -4413 -2106 -4408
rect -1538 -4413 -1464 -4408
rect 3200 -4458 3266 -4457
rect 6152 -4458 6226 -4453
rect 3200 -4462 6157 -4458
rect -2296 -4510 -2222 -4505
rect -2088 -4510 -2014 -4506
rect -2296 -4574 -2291 -4510
rect -2227 -4511 -2014 -4510
rect -2227 -4574 -2083 -4511
rect -2296 -4579 -2222 -4574
rect -2088 -4575 -2083 -4574
rect -2019 -4575 -2014 -4511
rect 3200 -4518 3205 -4462
rect 3261 -4518 6157 -4462
rect 3200 -4522 6157 -4518
rect 6221 -4522 6226 -4458
rect 3200 -4523 3266 -4522
rect 6152 -4527 6226 -4522
rect -2088 -4580 -2014 -4575
rect 3742 -4612 3808 -4611
rect 6298 -4612 6372 -4607
rect 3742 -4616 6303 -4612
rect 3742 -4672 3747 -4616
rect 3803 -4672 6303 -4616
rect 3742 -4676 6303 -4672
rect 6367 -4676 6372 -4612
rect 3742 -4677 3808 -4676
rect 6298 -4681 6372 -4676
rect 4270 -4796 4336 -4795
rect 8264 -4796 8338 -4791
rect 4270 -4800 8269 -4796
rect -1008 -4825 -929 -4821
rect -1008 -4826 -112 -4825
rect -1008 -4895 -1003 -4826
rect -934 -4830 -112 -4826
rect -934 -4889 -173 -4830
rect -117 -4889 -112 -4830
rect 4270 -4856 4275 -4800
rect 4331 -4856 8269 -4800
rect 4270 -4860 8269 -4856
rect 8333 -4860 8338 -4796
rect 4270 -4861 4336 -4860
rect 8264 -4865 8338 -4860
rect -934 -4894 -112 -4889
rect -934 -4895 -929 -4894
rect -1008 -4900 -929 -4895
rect 4419 -4984 4493 -4979
rect 8416 -4984 8482 -4983
rect -475 -5033 -401 -5028
rect -18 -5033 48 -5032
rect -475 -5097 -470 -5033
rect -406 -5037 48 -5033
rect -406 -5093 -13 -5037
rect 43 -5093 48 -5037
rect 4419 -5048 4424 -4984
rect 4488 -4988 8482 -4984
rect 4488 -5044 8421 -4988
rect 8477 -5044 8482 -4988
rect 4488 -5048 8482 -5044
rect 4419 -5053 4493 -5048
rect 8416 -5049 8482 -5048
rect -406 -5097 48 -5093
rect -475 -5102 -401 -5097
rect -18 -5098 48 -5097
rect 4566 -5188 4640 -5183
rect 10379 -5188 10445 -5187
rect 67 -5202 141 -5197
rect 1071 -5202 1137 -5201
rect 67 -5266 72 -5202
rect 136 -5206 1137 -5202
rect 136 -5262 1076 -5206
rect 1132 -5262 1137 -5206
rect 4566 -5252 4571 -5188
rect 4635 -5192 10445 -5188
rect 4635 -5248 10384 -5192
rect 10440 -5248 10445 -5192
rect 4635 -5252 10445 -5248
rect 4566 -5257 4640 -5252
rect 10379 -5253 10445 -5252
rect 136 -5266 1137 -5262
rect 67 -5271 141 -5266
rect 1071 -5267 1137 -5266
rect 588 -5367 662 -5362
rect 1593 -5367 1659 -5366
rect 588 -5431 593 -5367
rect 657 -5371 1659 -5367
rect 657 -5427 1598 -5371
rect 1654 -5427 1659 -5371
rect 657 -5431 1659 -5427
rect 588 -5436 662 -5431
rect 1593 -5432 1659 -5431
rect 1131 -5543 1205 -5538
rect 2136 -5543 2202 -5542
rect 1131 -5607 1136 -5543
rect 1200 -5547 2202 -5543
rect 1200 -5603 2141 -5547
rect 2197 -5603 2202 -5547
rect 1200 -5607 2202 -5603
rect 1131 -5612 1205 -5607
rect 2136 -5608 2202 -5607
rect 1660 -5732 1734 -5727
rect 2664 -5732 2730 -5731
rect 1660 -5796 1665 -5732
rect 1729 -5736 2730 -5732
rect 1729 -5792 2669 -5736
rect 2725 -5792 2730 -5736
rect 1729 -5796 2730 -5792
rect 1660 -5801 1734 -5796
rect 2664 -5797 2730 -5796
rect 2196 -5925 2270 -5920
rect 3202 -5925 3268 -5924
rect 2196 -5989 2201 -5925
rect 2265 -5929 3268 -5925
rect 2265 -5985 3207 -5929
rect 3263 -5985 3268 -5929
rect 2265 -5989 3268 -5985
rect 2196 -5994 2270 -5989
rect 3202 -5990 3268 -5989
rect 2738 -6094 2812 -6089
rect 3745 -6094 3811 -6093
rect 2738 -6158 2743 -6094
rect 2807 -6098 3811 -6094
rect 2807 -6154 3750 -6098
rect 3806 -6154 3811 -6098
rect 2807 -6158 3811 -6154
rect 2738 -6163 2812 -6158
rect 3745 -6159 3811 -6158
rect 3266 -6270 3340 -6265
rect 4271 -6270 4337 -6269
rect 3266 -6334 3271 -6270
rect 3335 -6274 4337 -6270
rect 3335 -6330 4276 -6274
rect 4332 -6330 4337 -6274
rect 3335 -6334 4337 -6330
rect 3266 -6339 3340 -6334
rect 4271 -6335 4337 -6334
rect 3796 -6421 3870 -6416
rect 4423 -6421 4489 -6420
rect 3796 -6485 3801 -6421
rect 3865 -6425 4489 -6421
rect 3865 -6481 4428 -6425
rect 4484 -6481 4489 -6425
rect 3865 -6485 4489 -6481
rect 3796 -6490 3870 -6485
rect 4423 -6486 4489 -6485
rect -7730 -6600 -7616 -6595
rect -7730 -6704 -7725 -6600
rect -7621 -6704 11086 -6600
rect 11190 -6704 11196 -6600
rect -7730 -6709 -7616 -6704
rect -3671 -7152 -3605 -7151
rect -6410 -7156 -3605 -7152
rect -6410 -7158 -3666 -7156
rect -6410 -7222 -6405 -7158
rect -6341 -7212 -3666 -7158
rect -3610 -7212 -3605 -7156
rect -6341 -7216 -3605 -7212
rect -6341 -7222 -6336 -7216
rect -3671 -7217 -3605 -7216
rect -6410 -7227 -6336 -7222
rect -6520 -7297 -6446 -7292
rect -6520 -7361 -6515 -7297
rect -6451 -7298 -6446 -7297
rect -4217 -7298 -4151 -7297
rect -6451 -7302 -4151 -7298
rect -6451 -7358 -4212 -7302
rect -4156 -7358 -4151 -7302
rect -6451 -7361 -4151 -7358
rect -6520 -7362 -4151 -7361
rect -6520 -7366 -6446 -7362
rect -4217 -7363 -4151 -7362
rect -26749 -7520 -26683 -7519
rect -13163 -7520 -13097 -7519
rect -5089 -7520 -5023 -7519
rect 4570 -7520 4636 -7519
rect -26749 -7524 4636 -7520
rect -26749 -7580 -26744 -7524
rect -26688 -7580 -13158 -7524
rect -13102 -7580 -5084 -7524
rect -5028 -7580 4575 -7524
rect 4631 -7580 4636 -7524
rect -26749 -7584 4636 -7580
rect -26749 -7585 -26683 -7584
rect -13163 -7585 -13097 -7584
rect -5089 -7585 -5023 -7584
rect 4570 -7585 4636 -7584
rect -18591 -8042 -18525 -8039
rect -4395 -8042 -4325 -8037
rect -18591 -8044 -4390 -8042
rect -18591 -8100 -18586 -8044
rect -18530 -8100 -4390 -8044
rect -18591 -8102 -4390 -8100
rect -4330 -8102 -4325 -8042
rect -18591 -8105 -18525 -8102
rect -4395 -8107 -4325 -8102
rect -8863 -9035 -8857 -8897
rect -8729 -8902 -8719 -8897
rect -8724 -9030 -8719 -8902
rect -4393 -8902 -4327 -8899
rect -4393 -8904 -3729 -8902
rect -4393 -8960 -4388 -8904
rect -4332 -8960 -3729 -8904
rect -4393 -8962 -3729 -8960
rect 3724 -8962 3784 -8902
rect -4393 -8965 -4327 -8962
rect -8729 -9035 -8719 -9030
rect -16488 -11756 -16422 -11753
rect 420 -11756 490 -11751
rect -16488 -11758 425 -11756
rect -16488 -11814 -16483 -11758
rect -16427 -11814 425 -11758
rect -16488 -11816 425 -11814
rect 485 -11816 490 -11756
rect -16488 -11819 -16422 -11816
rect 420 -11821 490 -11816
rect -29124 -11876 -27982 -11871
rect -29124 -12014 -29119 -11876
rect -28981 -12014 -27982 -11876
rect -29124 -12019 -27982 -12014
rect -28015 -14558 -27949 -14557
rect -26753 -14558 -26679 -14553
rect -28015 -14562 -27674 -14558
rect -28015 -14618 -28010 -14562
rect -27954 -14618 -27674 -14562
rect -28015 -14622 -27674 -14618
rect -27566 -14622 -26748 -14558
rect -26684 -14622 -26679 -14558
rect -28015 -14623 -27949 -14622
rect -26753 -14627 -26679 -14622
rect -28587 -15257 -28521 -15256
rect -28233 -15257 -28159 -15252
rect -28587 -15261 -28228 -15257
rect -28587 -15317 -28582 -15261
rect -28526 -15317 -28228 -15261
rect -28587 -15321 -28228 -15317
rect -28164 -15321 -28159 -15257
rect -28587 -15322 -28521 -15321
rect -28233 -15326 -28159 -15321
rect -26914 -16276 -26844 -16271
rect -28135 -16336 -26909 -16276
rect -26849 -16336 -26844 -16276
rect -26914 -16341 -26844 -16336
rect -28686 -17210 -27544 -17205
rect -28686 -17348 -28681 -17210
rect -28543 -17348 -27544 -17210
rect -28686 -17353 -27544 -17348
rect -18244 -18509 -18174 -18504
rect -19239 -18569 -18239 -18509
rect -18179 -18569 -18174 -18509
rect -18244 -18574 -18174 -18569
rect -16490 -18711 -16420 -18706
rect -19239 -18771 -16485 -18711
rect -16425 -18771 -16420 -18711
rect -16490 -18776 -16420 -18771
rect -9257 -21941 -9119 -21936
rect -9257 -21963 -9252 -21941
rect -10861 -21968 -9252 -21963
rect -10861 -22047 -10856 -21968
rect -10777 -22047 -9252 -21968
rect -10861 -22052 -9252 -22047
rect -9257 -22069 -9252 -22052
rect -9124 -22069 -9119 -21941
rect -9257 -22074 -9119 -22069
rect -8857 -22947 -8719 -22942
rect -10543 -22952 -8852 -22947
rect -10543 -23070 -10538 -22952
rect -10420 -23070 -8852 -22952
rect -10543 -23075 -8852 -23070
rect -8724 -23075 -8719 -22947
rect -8857 -23080 -8719 -23075
rect -28682 -23307 -27348 -23302
rect -28682 -23445 -28677 -23307
rect -28539 -23445 -27348 -23307
rect -28682 -23450 -27348 -23445
<< via3 >>
rect 11086 -6704 11190 -6600
rect -8857 -8902 -8729 -8897
rect -8857 -9030 -8852 -8902
rect -8852 -9030 -8729 -8902
rect -8857 -9035 -8729 -9030
<< metal4 >>
rect 11085 -6600 11191 -6599
rect 11085 -6704 11086 -6600
rect 11190 -6704 11191 -6600
rect 11085 -6705 11191 -6704
rect 11086 -12043 11190 -6705
rect 11081 -12112 11190 -12043
rect 11081 -12941 11185 -12112
<< via4 >>
rect -8953 -8897 -8633 -8806
rect -8953 -9035 -8857 -8897
rect -8857 -9035 -8729 -8897
rect -8729 -9035 -8633 -8897
rect -8953 -9126 -8633 -9035
rect 10973 -13261 11293 -12941
<< metal5 >>
rect -8977 -8806 -8609 -8782
rect -8977 -9126 -8953 -8806
rect -8633 -9126 -8609 -8806
rect -8977 -9458 -8609 -9126
rect 10949 -12938 11317 -12917
rect 10345 -12941 11317 -12938
rect 10345 -13258 10973 -12941
rect 10949 -13261 10973 -13258
rect 11293 -13261 11317 -12941
rect 10949 -13285 11317 -13261
use comparator  comparator_0
timestamp 1713454396
transform 1 0 -27530 0 1 -21626
box -811 -2117 11035 9755
use comparator  comparator_1
timestamp 1713454396
transform 1 0 -26517 0 1 3604
box -811 -2117 11035 9755
use ibias_gen  ibias_gen_0
timestamp 1713454396
transform 1 0 -27321 0 1 -10450
box -138 -652 15828 11500
use rc_osc_por  rc_osc_por_0
timestamp 1713454396
transform 1 0 -12543 0 1 -23191
box -14232 -2658 25847 4148
use rstring_mux  rstring_mux_0
timestamp 1713454396
transform 1 0 -16753 0 1 -15968
box 464 -3512 27160 9182
use schmitt_trigger  schmitt_trigger_0
timestamp 1713454396
transform 1 0 -4393 0 1 2578
box -91 -52 2297 1163
use sky130_fd_pr__cap_mim_m3_2_LUWKLG  sky130_fd_pr__cap_mim_m3_2_LUWKLG_0
timestamp 1712463840
transform 0 -1 -8855 1 0 -12829
box -3349 -19200 3371 19200
use sky130_fd_pr__res_xhigh_po_1p41_DVQADA  sky130_fd_pr__res_xhigh_po_1p41_DVQADA_0
timestamp 1712352531
transform 1 0 -11267 0 1 5911
box -3898 -4082 3898 4082
use sky130_fd_pr__rf_pnp_05v5_W0p68L0p68  sky130_fd_pr__rf_pnp_05v5_W0p68L0p68_0 $PDKPATH/libs.ref/sky130_fd_pr/mag
timestamp 1712845802
transform 1 0 -4157 0 1 11478
box 0 0 796 796
use sky130_fd_sc_hd__inv_4  sky130_fd_sc_hd__inv_4_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712845802
transform 1 0 -4350 0 1 1782
box -38 -48 498 592
use sky130_fd_sc_hd__inv_4  sky130_fd_sc_hd__inv_4_1
timestamp 1712845802
transform 1 0 -3890 0 1 1033
box -38 -48 498 592
use sky130_fd_sc_hd__inv_4  sky130_fd_sc_hd__inv_4_2
timestamp 1712845802
transform 1 0 -4350 0 1 1033
box -38 -48 498 592
use sky130_fd_sc_hd__inv_4  sky130_fd_sc_hd__inv_4_3
timestamp 1712845802
transform 1 0 -4350 0 1 3931
box -38 -48 498 592
use sky130_fd_sc_hd__inv_4  sky130_fd_sc_hd__inv_4_4
timestamp 1712845802
transform 1 0 -4350 0 1 4758
box -38 -48 498 592
use sky130_fd_sc_hd__inv_16  sky130_fd_sc_hd__inv_16_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712845802
transform 1 0 -3890 0 1 1782
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_16  sky130_fd_sc_hd__inv_16_1
timestamp 1712845802
transform 1 0 -3430 0 1 1033
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_16  sky130_fd_sc_hd__inv_16_2
timestamp 1712845802
transform 1 0 -3890 0 1 3931
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_16  sky130_fd_sc_hd__inv_16_3
timestamp 1712845802
transform 1 0 -3890 0 1 4758
box -38 -48 1510 592
use sky130_fd_sc_hvl__inv_1  sky130_fd_sc_hvl__inv_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1712845802
transform 1 0 -11417 0 1 11008
box -66 -43 354 897
use sky130_fd_sc_hvl__inv_4  sky130_fd_sc_hvl__inv_4_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1712845802
transform 1 0 -11129 0 1 11008
box -66 -43 834 897
use sky130_fd_sc_hvl__inv_16  sky130_fd_sc_hvl__inv_16_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1712845802
transform 1 0 -10361 0 1 11008
box -66 -43 2754 897
use sky130_fd_sc_hvl__lsbufhv2lv_1  sky130_fd_sc_hvl__lsbufhv2lv_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1712845802
transform 1 0 10485 0 1 -2363
box -66 -43 1698 1671
use sky130_fd_sc_hvl__lsbufhv2lv_1  sky130_fd_sc_hvl__lsbufhv2lv_1_1
timestamp 1712845802
transform 1 0 10484 0 1 -4097
box -66 -43 1698 1671
use sky130_fd_sc_hvl__lsbuflv2hv_1  sky130_fd_sc_hvl__lsbuflv2hv_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
array 0 8 2112 0 1 1734
timestamp 1712845802
transform 1 0 -8523 0 1 -4097
box -66 -43 2178 1671
use sky130_fd_sc_hvl__lsbuflv2hv_1  sky130_fd_sc_hvl__lsbuflv2hv_1_1
timestamp 1712845802
transform 1 0 -4282 0 1 6638
box -66 -43 2178 1671
<< labels >>
flabel metal1 s -4580 -7558 -4580 -7558 0 FreeSans 1200 0 0 0 avss
port 13 nsew
flabel metal2 -17531 753 -17531 753 0 FreeSans 1200 0 0 0 itest
port 12 nsew
flabel metal2 s -18241 -2814 -18241 -2814 0 FreeSans 1200 0 0 0 vbg_1v2
port 10 nsew
flabel metal2 -15287 -2068 -15287 -2068 0 FreeSans 1200 0 0 0 ibg_200n
port 14 nsew
flabel metal3 10912 -1837 10912 -1837 0 FreeSans 800 0 0 0 vl
flabel metal2 s 8849 -2119 8909 -2059 0 FreeSans 1200 0 0 0 isrc_sel
port 19 nsew
flabel metal1 s -3836 -4436 -3836 -4436 0 FreeSans 1200 0 0 0 dvdd
port 16 nsew
flabel metal1 s -3836 -4646 -3836 -4646 0 FreeSans 1200 0 0 0 avdd
port 11 nsew
flabel metal2 s -8047 -2119 -8047 -2119 0 FreeSans 1200 0 0 0 otrip_decoded[1]
port 8 nsew
flabel metal2 s -5935 -2119 -5935 -2119 0 FreeSans 1200 0 0 0 otrip_decoded[3]
port 6 nsew
flabel metal2 s -3823 -2119 -3823 -2119 0 FreeSans 1200 0 0 0 otrip_decoded[5]
port 4 nsew
flabel metal2 s -1711 -2119 -1711 -2119 0 FreeSans 1200 0 0 0 otrip_decoded[7]
port 2 nsew
flabel metal2 s -1711 -3853 -1711 -3853 0 FreeSans 1200 0 0 0 otrip_decoded[6]
port 3 nsew
flabel metal2 s -3823 -3853 -3823 -3853 0 FreeSans 1200 0 0 0 otrip_decoded[4]
port 5 nsew
flabel metal2 s -5935 -3853 -5935 -3853 0 FreeSans 1200 0 0 0 otrip_decoded[2]
port 7 nsew
flabel metal2 s -8047 -3853 -8047 -3853 0 FreeSans 1200 0 0 0 otrip_decoded[0]
port 9 nsew
flabel metal3 s 10400 -1728 10400 -1728 0 FreeSans 800 0 0 0 dcomp3v3
flabel metal3 s 10506 -3684 10506 -3684 0 FreeSans 800 0 0 0 dcomp3v3uv
flabel metal2 s -2438 4175 -2438 4175 0 FreeSans 1200 0 0 0 dcomp
port 18 nsew
flabel metal2 s -10817 -22202 -10817 -22202 0 FreeSans 1200 0 0 0 osc_ck
port 21 nsew
flabel metal2 -14211 -22364 -14211 -22364 0 FreeSans 1200 0 0 0 osc_ena
port 22 nsew
flabel metal2 s 8849 -3853 8909 -3793 0 FreeSans 1200 0 0 0 force_pdnb
port 15 nsew
flabel metal2 -2411 1988 -2411 1988 0 FreeSans 1200 0 0 0 pwup_filt
port 20 nsew
flabel metal2 s -2438 5002 -2438 5002 0 FreeSans 1200 0 0 0 por
port 25 nsew
flabel metal2 s -7927 11519 -7927 11519 0 FreeSans 1200 0 0 0 porb_h
port 23 nsew
flabel metal3 s -2178 -8855 -2178 -8855 0 FreeSans 1200 0 0 0 vin
port 1 nsew
flabel metal2 -4579 1551 -4579 1551 0 FreeSans 1200 0 0 0 dvss
port 17 nsew
flabel metal2 s -1997 1269 -1997 1269 0 FreeSans 1200 0 0 0 porb
port 26 nsew
flabel metal2 s -4279 1160 -4279 1160 0 FreeSans 1200 0 0 0 por_unbuf
port 24 nsew
<< properties >>
string MASKHINTS_PSDM -8549 -2512 12143 -2320
<< end >>
