* XSpice netlist created from SPICE and liberty sources by spi2xspice.py
* NGSPICE file created from por_dig.ext - technology: sky130A
* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt por_dig a_VGND a_VPWR a_force_pdn a_force_pdnb a_force_rc_osc a_force_short_oneshot a_osc_ck a_osc_ena a_otrip_0_ a_otrip_1_ a_otrip_2_ a_otrip_decoded_0_ a_otrip_decoded_1_ a_otrip_decoded_2_ a_otrip_decoded_3_ a_otrip_decoded_4_ a_otrip_decoded_5_ a_otrip_decoded_6_ a_otrip_decoded_7_ a_por_timed_out a_por_unbuf a_pwup_filt a_startup_timed_out
A_062_ [net6 net4 net5] net12 d_lut_sky130_fd_sc_hd__nor3b_1
A_114_ _005_ clknet_1_1__leaf_osc_ck NULL ~net23 cnt_por\_0\_ NULL ddflop
Aoutput20 [net20] startup_timed_out d_lut_sky130_fd_sc_hd__buf_2
A_113_ _004_ clknet_1_1__leaf_osc_ck NULL ~net23 cnt_st\_4\_ NULL ddflop
A_061_ [net6 net5 net4] net11 d_lut_sky130_fd_sc_hd__nor3b_1
Aoutput8 [net8] force_pdnb d_lut_sky130_fd_sc_hd__buf_2
Aoutput10 [net10] otrip_decoded_0_ d_lut_sky130_fd_sc_hd__buf_2
A_060_ [net6 net5 net4] net10 d_lut_sky130_fd_sc_hd__nor3_1
A_112_ _003_ clknet_1_1__leaf_osc_ck NULL ~net23 cnt_st\_3\_ NULL ddflop
Ahold10 [cnt_por\_8\_] net34 d_lut_sky130_fd_sc_hd__dlygate4sd3_1
Aoutput9 [net9] osc_ena d_lut_sky130_fd_sc_hd__buf_2
Aoutput11 [net11] otrip_decoded_1_ d_lut_sky130_fd_sc_hd__buf_2
A_111_ _002_ clknet_1_1__leaf_osc_ck NULL ~net23 cnt_st\_2\_ NULL ddflop
Ahold11 [cnt_por\_1\_] net35 d_lut_sky130_fd_sc_hd__dlygate4sd3_1
Aoutput12 [net12] otrip_decoded_2_ d_lut_sky130_fd_sc_hd__buf_2
A_125__240 net24 done
A_125__241 _125__24/LO dzero
Ahold12 [cnt_st\_4\_] net36 d_lut_sky130_fd_sc_hd__dlygate4sd3_1
A_110_ _001_ clknet_1_1__leaf_osc_ck NULL ~net22 cnt_st\_1\_ NULL ddflop
Aoutput13 [net13] otrip_decoded_3_ d_lut_sky130_fd_sc_hd__buf_2
Ahold13 [cnt_por\_0\_] net37 d_lut_sky130_fd_sc_hd__dlygate4sd3_1
Aoutput14 [net14] otrip_decoded_4_ d_lut_sky130_fd_sc_hd__buf_2
A_099_ [_017_ _018_] _010_ d_lut_sky130_fd_sc_hd__nor2_1
Aoutput15 [net15] otrip_decoded_5_ d_lut_sky130_fd_sc_hd__buf_2
A_098_ [net21 _016_ net32] _018_ d_lut_sky130_fd_sc_hd__a21oi_1
Aoutput16 [net16] otrip_decoded_6_ d_lut_sky130_fd_sc_hd__buf_2
A_097_ [cnt_por\_5\_ net21 _016_] _017_ d_lut_sky130_fd_sc_hd__and3_1
Aoutput17 [net17] otrip_decoded_7_ d_lut_sky130_fd_sc_hd__buf_2
A_096_ [cnt_por\_4\_ _026_ _027_ net3] _016_ d_lut_sky130_fd_sc_hd__a31o_1
Aoutput18 [net18] por_timed_out d_lut_sky130_fd_sc_hd__buf_2
A_079_ [net31 _035_ _037_] _003_ d_lut_sky130_fd_sc_hd__o21ai_1
A_095_ [net3 net21 _047_] _009_ d_lut_sky130_fd_sc_hd__a21o_1
Aoutput19 [net19] por_unbuf d_lut_sky130_fd_sc_hd__clkbuf_4
A_078_ [net31 _035_ net20] _037_ d_lut_sky130_fd_sc_hd__a21oi_1
Afanout21 [net19] net21 d_lut_sky130_fd_sc_hd__clkbuf_2
A_094_ [cnt_por\_4\_ _046_] _047_ d_lut_sky130_fd_sc_hd__xor2_1
A_077_ [_035_ _036_ net20] _002_ d_lut_sky130_fd_sc_hd__a21o_1
A_093_ [_045_ _046_ net3 net21] _008_ d_lut_sky130_fd_sc_hd__a2bb2o_1
Afanout22 [net25] net22 d_lut_sky130_fd_sc_hd__clkbuf_4
Ainput1 [force_pdn] net1 d_lut_sky130_fd_sc_hd__clkbuf_1
A_076_ [cnt_st\_2\_ _032_] _036_ d_lut_sky130_fd_sc_hd__or2_1
A_059_ [_028_ _031_] net18 d_lut_sky130_fd_sc_hd__nor2_1
Afanout23 [net25] net23 d_lut_sky130_fd_sc_hd__clkbuf_2
A_092_ [_028_ _031_ net20 _026_ _027_] _046_ d_lut_sky130_fd_sc_hd__o2111a_1
Ainput2 [force_rc_osc] net2 d_lut_sky130_fd_sc_hd__clkbuf_1
A_058_ [_029_ _030_] _031_ d_lut_sky130_fd_sc_hd__nand2_1
A_127_ net27 clknet_1_0__leaf_osc_ck NULL ~net7 cnt_rsb NULL ddflop
A_075_ [cnt_st\_2\_ _032_] _035_ d_lut_sky130_fd_sc_hd__nand2_1
A_091_ [cnt_por\_2\_ _026_ net21 cnt_por\_3\_] _045_ d_lut_sky130_fd_sc_hd__a31oi_1
Ainput3 [force_short_oneshot] net3 d_lut_sky130_fd_sc_hd__clkbuf_2
A_074_ [_033_ _034_ net20] _001_ d_lut_sky130_fd_sc_hd__a21o_1
A_126_ net26 clknet_1_0__leaf_osc_ck NULL ~net7 cnt_rsb_stg2 NULL ddflop
A_057_ [cnt_por\_7\_ cnt_por\_9\_ cnt_por\_8\_ cnt_por\_10\_] _030_ d_lut_sky130_fd_sc_hd__and4_1
A_109_ _000_ clknet_1_1__leaf_osc_ck NULL ~net22 cnt_st\_0\_ NULL ddflop
A_090_ [net3 net19 _043_ _044_] _007_ d_lut_sky130_fd_sc_hd__a22o_1
Ainput4 [otrip_0_] net4 d_lut_sky130_fd_sc_hd__dlymetal6s2s_1
A_056_ [cnt_por\_5\_ cnt_por\_6\_] _029_ d_lut_sky130_fd_sc_hd__and2_1
A_125_ net24 clknet_1_0__leaf_osc_ck NULL ~net7 cnt_rsb_stg1 NULL ddflop
A_073_ [cnt_st\_1\_ cnt_st\_0\_ net3] _034_ d_lut_sky130_fd_sc_hd__or3_1
A_108_ [net29 _022_] _015_ d_lut_sky130_fd_sc_hd__xor2_1
Ainput5 [otrip_1_] net5 d_lut_sky130_fd_sc_hd__dlymetal6s2s_1
A_072_ [_032_] _033_ d_lut_sky130_fd_sc_hd__inv_2
A_055_ [cnt_por\_4\_ _026_ _027_] _028_ d_lut_sky130_fd_sc_hd__nand3_1
A_124_ _015_ clknet_1_1__leaf_osc_ck NULL ~net22 cnt_por\_10\_ NULL ddflop
A_107_ [net30 _020_] _014_ d_lut_sky130_fd_sc_hd__xor2_1
Ainput6 [otrip_2_] net6 d_lut_sky130_fd_sc_hd__dlymetal6s2s_1
A_071_ [cnt_st\_0\_ net3 cnt_st\_1\_] _032_ d_lut_sky130_fd_sc_hd__o21a_1
A_054_ [cnt_por\_3\_ cnt_por\_2\_] _027_ d_lut_sky130_fd_sc_hd__and2_1
A_123_ _014_ clknet_1_0__leaf_osc_ck NULL ~net22 cnt_por\_9\_ NULL ddflop
A_106_ [cnt_por\_7\_ cnt_por\_9\_ cnt_por\_8\_ _019_] _022_ d_lut_sky130_fd_sc_hd__and4_1
Ainput7 [pwup_filt] net7 d_lut_sky130_fd_sc_hd__dlymetal6s2s_1
A_070_ [net3 net20 cnt_st\_0\_] _000_ d_lut_sky130_fd_sc_hd__or3b_1
A_053_ [cnt_por\_1\_ cnt_por\_0\_] _026_ d_lut_sky130_fd_sc_hd__and2_2
A_122_ _013_ clknet_1_0__leaf_osc_ck NULL ~net22 cnt_por\_8\_ NULL ddflop
A_105_ [_020_ _021_] _013_ d_lut_sky130_fd_sc_hd__nor2_1
Aclkbuf_1_1__f_osc_ck [clknet_0_osc_ck] clknet_1_1__leaf_osc_ck d_lut_sky130_fd_sc_hd__clkbuf_16
A_052_ [cnt_st\_4\_ _025_] net20 d_lut_sky130_fd_sc_hd__and2_2
A_121_ _012_ clknet_1_0__leaf_osc_ck NULL ~net22 cnt_por\_7\_ NULL ddflop
A_104_ [cnt_por\_7\_ _019_ net34] _021_ d_lut_sky130_fd_sc_hd__a21oi_1
A_120_ _011_ clknet_1_0__leaf_osc_ck NULL ~net22 cnt_por\_6\_ NULL ddflop
A_051_ [cnt_st\_1\_ cnt_st\_0\_ cnt_st\_2\_ cnt_st\_3\_] _025_ d_lut_sky130_fd_sc_hd__and4_1
A_103_ [cnt_por\_7\_ cnt_por\_8\_ _019_] _020_ d_lut_sky130_fd_sc_hd__and3_1
Ahold1 [cnt_rsb] net25 d_lut_sky130_fd_sc_hd__dlygate4sd3_1
Aclkbuf_0_osc_ck [osc_ck] clknet_0_osc_ck d_lut_sky130_fd_sc_hd__clkbuf_16
A_050_ [net7] _024_ d_lut_sky130_fd_sc_hd__inv_2
A_102_ [net33 _019_] _012_ d_lut_sky130_fd_sc_hd__xor2_1
Ahold2 [cnt_rsb_stg1] net26 d_lut_sky130_fd_sc_hd__dlygate4sd3_1
A_101_ [net28 _017_] _011_ d_lut_sky130_fd_sc_hd__xor2_1
Ahold3 [cnt_rsb_stg2] net27 d_lut_sky130_fd_sc_hd__dlygate4sd3_1
A_100_ [_028_ _031_ _016_ _029_ net20] _019_ d_lut_sky130_fd_sc_hd__o2111a_1
Ahold4 [cnt_por\_6\_] net28 d_lut_sky130_fd_sc_hd__dlygate4sd3_1
Ahold5 [cnt_por\_10\_] net29 d_lut_sky130_fd_sc_hd__dlygate4sd3_1
A_089_ [_026_ net19 cnt_por\_2\_] _044_ d_lut_sky130_fd_sc_hd__a21o_1
Ahold6 [cnt_por\_9\_] net30 d_lut_sky130_fd_sc_hd__dlygate4sd3_1
A_088_ [cnt_por\_2\_ _026_ net19] _043_ d_lut_sky130_fd_sc_hd__nand3_1
Ahold7 [cnt_st\_3\_] net31 d_lut_sky130_fd_sc_hd__dlygate4sd3_1
Ahold8 [cnt_por\_5\_] net32 d_lut_sky130_fd_sc_hd__dlygate4sd3_1
A_087_ [net3 net21 _041_ _042_] _006_ d_lut_sky130_fd_sc_hd__a22o_1
Aclkbuf_1_0__f_osc_ck [clknet_0_osc_ck] clknet_1_0__leaf_osc_ck d_lut_sky130_fd_sc_hd__clkbuf_16
A_086_ [cnt_por\_0\_ net21 net35] _042_ d_lut_sky130_fd_sc_hd__a21o_1
A_069_ [_028_ _031_ net20] net19 d_lut_sky130_fd_sc_hd__o21a_1
Ahold9 [cnt_por\_7\_] net33 d_lut_sky130_fd_sc_hd__dlygate4sd3_1
A_085_ [_026_ net21] _041_ d_lut_sky130_fd_sc_hd__nand2_1
A_068_ [_024_ net18 net2] net9 d_lut_sky130_fd_sc_hd__o21bai_1
A_084_ [net21 _040_ net37] _005_ d_lut_sky130_fd_sc_hd__mux2_1
A_067_ [net6 net5 net4] net17 d_lut_sky130_fd_sc_hd__and3_1
A_119_ _010_ clknet_1_0__leaf_osc_ck NULL ~net22 cnt_por\_5\_ NULL ddflop
A_083_ [net3 net21] _040_ d_lut_sky130_fd_sc_hd__nand2b_1
A_049_ [net1] net8 d_lut_sky130_fd_sc_hd__inv_2
A_118_ _009_ clknet_1_1__leaf_osc_ck NULL ~net22 cnt_por\_4\_ NULL ddflop
A_066_ [net4 net5 net6] net16 d_lut_sky130_fd_sc_hd__and3b_1
A_082_ [_023_ _038_ _039_] _004_ d_lut_sky130_fd_sc_hd__o21ai_1
A_065_ [net5 net4 net6] net15 d_lut_sky130_fd_sc_hd__and3b_1
A_117_ _008_ clknet_1_1__leaf_osc_ck NULL ~net22 cnt_por\_3\_ NULL ddflop
A_048_ [net36] _023_ d_lut_sky130_fd_sc_hd__inv_2
A_081_ [_023_ _038_ _025_] _039_ d_lut_sky130_fd_sc_hd__a21oi_1
A_064_ [net5 net4 net6] net14 d_lut_sky130_fd_sc_hd__nor3b_1
A_116_ _007_ clknet_1_1__leaf_osc_ck NULL ~net23 cnt_por\_2\_ NULL ddflop
A_080_ [cnt_st\_1\_ cnt_st\_2\_ cnt_st\_3\_ net3] _038_ d_lut_sky130_fd_sc_hd__and4_1
A_063_ [net6 net5 net4] net13 d_lut_sky130_fd_sc_hd__and3b_1
A_115_ _006_ clknet_1_1__leaf_osc_ck NULL ~net23 cnt_por\_1\_ NULL ddflop

.model todig_1v8 adc_bridge(in_high=1.2 in_low=0.6 rise_delay=10n fall_delay=10n)
.model toana_1v8 dac_bridge(out_high=1.8 out_low=0)

.model ddflop d_dff(ic=0 rise_delay=1n fall_delay=1n)
.model dlatch d_dlatch(ic=0 rise_delay=1n fall_delay=1n)
.model dzero d_pulldown(load=1p)
.model done d_pullup(load=1p)

AA2D1 [a_VGND] [VGND] todig_1v8
AA2D2 [a_VPWR] [VPWR] todig_1v8
AA2D3 [a_force_pdn] [force_pdn] todig_1v8
AD2A1 [force_pdnb] [a_force_pdnb] toana_1v8
AA2D4 [a_force_rc_osc] [force_rc_osc] todig_1v8
AA2D5 [a_force_short_oneshot] [force_short_oneshot] todig_1v8
AA2D6 [a_osc_ck] [osc_ck] todig_1v8
AD2A2 [osc_ena] [a_osc_ena] toana_1v8
AA2D7 [a_otrip_0_] [otrip_0_] todig_1v8
AA2D8 [a_otrip_1_] [otrip_1_] todig_1v8
AA2D9 [a_otrip_2_] [otrip_2_] todig_1v8
AD2A3 [otrip_decoded_0_] [a_otrip_decoded_0_] toana_1v8
AD2A4 [otrip_decoded_1_] [a_otrip_decoded_1_] toana_1v8
AD2A5 [otrip_decoded_2_] [a_otrip_decoded_2_] toana_1v8
AD2A6 [otrip_decoded_3_] [a_otrip_decoded_3_] toana_1v8
AD2A7 [otrip_decoded_4_] [a_otrip_decoded_4_] toana_1v8
AD2A8 [otrip_decoded_5_] [a_otrip_decoded_5_] toana_1v8
AD2A9 [otrip_decoded_6_] [a_otrip_decoded_6_] toana_1v8
AD2A10 [otrip_decoded_7_] [a_otrip_decoded_7_] toana_1v8
AD2A11 [por_timed_out] [a_por_timed_out] toana_1v8
AD2A12 [por_unbuf] [a_por_unbuf] toana_1v8
AA2D10 [a_pwup_filt] [pwup_filt] todig_1v8
AD2A13 [startup_timed_out] [a_startup_timed_out] toana_1v8

.ends


* sky130_fd_sc_hd__nor3b_1 (!A&!B&C_N)
.model d_lut_sky130_fd_sc_hd__nor3b_1 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "00001000")
* sky130_fd_sc_hd__fill_2 (no function)
* sky130_fd_sc_hd__decap_8 (no function)
* sky130_fd_sc_hd__dfrtp_1 IQ
* sky130_fd_sc_hd__fill_1 (no function)
* sky130_fd_sc_hd__buf_2 (A)
.model d_lut_sky130_fd_sc_hd__buf_2 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "01")
* sky130_fd_sc_hd__decap_4 (no function)
* sky130_fd_sc_hd__decap_3 (no function)
* sky130_fd_sc_hd__tapvpwrvgnd_1 (no function)
* sky130_fd_sc_hd__nor3_1 (!A&!B&!C)
.model d_lut_sky130_fd_sc_hd__nor3_1 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "10000000")
* sky130_fd_sc_hd__dlygate4sd3_1 (A)
.model d_lut_sky130_fd_sc_hd__dlygate4sd3_1 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "01")
* sky130_ef_sc_hd__decap_12 (no function)
* sky130_fd_sc_hd__conb_1 1
* sky130_fd_sc_hd__nor2_1 (!A&!B)
.model d_lut_sky130_fd_sc_hd__nor2_1 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "1000")
* sky130_fd_sc_hd__a21oi_1 (!A1&!B1) | (!A2&!B1)
.model d_lut_sky130_fd_sc_hd__a21oi_1 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "11100000")
* sky130_fd_sc_hd__and3_1 (A&B&C)
.model d_lut_sky130_fd_sc_hd__and3_1 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "00000001")
* sky130_fd_sc_hd__a31o_1 (A1&A2&A3) | (B1)
.model d_lut_sky130_fd_sc_hd__a31o_1 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "0000000111111111")
* sky130_fd_sc_hd__o21ai_1 (!A1&!A2) | (!B1)
.model d_lut_sky130_fd_sc_hd__o21ai_1 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "11111000")
* sky130_fd_sc_hd__a21o_1 (A1&A2) | (B1)
.model d_lut_sky130_fd_sc_hd__a21o_1 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "00011111")
* sky130_fd_sc_hd__clkbuf_4 (A)
.model d_lut_sky130_fd_sc_hd__clkbuf_4 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "01")
* sky130_fd_sc_hd__clkbuf_2 (A)
.model d_lut_sky130_fd_sc_hd__clkbuf_2 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "01")
* sky130_fd_sc_hd__xor2_1 (A&!B) | (!A&B)
.model d_lut_sky130_fd_sc_hd__xor2_1 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "0110")
* sky130_fd_sc_hd__a2bb2o_1 (B1&B2) | (!A1_N&!A2_N)
.model d_lut_sky130_fd_sc_hd__a2bb2o_1 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "1000100010001111")
* sky130_fd_sc_hd__clkbuf_1 (A)
.model d_lut_sky130_fd_sc_hd__clkbuf_1 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "01")
* sky130_fd_sc_hd__or2_1 (A) | (B)
.model d_lut_sky130_fd_sc_hd__or2_1 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "0111")
* sky130_fd_sc_hd__o2111a_1 (A1&B1&C1&D1) | (A2&B1&C1&D1)
.model d_lut_sky130_fd_sc_hd__o2111a_1 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "00000000000000000000000000000111")
* sky130_fd_sc_hd__nand2_1 (!A) | (!B)
.model d_lut_sky130_fd_sc_hd__nand2_1 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "1110")
* sky130_fd_sc_hd__a31oi_1 (!A1&!B1) | (!A2&!B1) | (!A3&!B1)
.model d_lut_sky130_fd_sc_hd__a31oi_1 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "1111111000000000")
* sky130_fd_sc_hd__and4_1 (A&B&C&D)
.model d_lut_sky130_fd_sc_hd__and4_1 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "0000000000000001")
* sky130_fd_sc_hd__a22o_1 (B1&B2) | (A1&A2)
.model d_lut_sky130_fd_sc_hd__a22o_1 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "0001000100011111")
* sky130_fd_sc_hd__dlymetal6s2s_1 (A)
.model d_lut_sky130_fd_sc_hd__dlymetal6s2s_1 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "01")
* sky130_fd_sc_hd__and2_1 (A&B)
.model d_lut_sky130_fd_sc_hd__and2_1 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "0001")
* sky130_fd_sc_hd__or3_1 (A) | (B) | (C)
.model d_lut_sky130_fd_sc_hd__or3_1 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "01111111")
* sky130_fd_sc_hd__decap_6 (no function)
* sky130_fd_sc_hd__inv_2 (!A)
.model d_lut_sky130_fd_sc_hd__inv_2 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "10")
* sky130_fd_sc_hd__nand3_1 (!A) | (!B) | (!C)
.model d_lut_sky130_fd_sc_hd__nand3_1 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "11111110")
* sky130_fd_sc_hd__o21a_1 (A1&B1) | (A2&B1)
.model d_lut_sky130_fd_sc_hd__o21a_1 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "00000111")
* sky130_fd_sc_hd__or3b_1 (A) | (B) | (!C_N)
.model d_lut_sky130_fd_sc_hd__or3b_1 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "11110111")
* sky130_fd_sc_hd__and2_2 (A&B)
.model d_lut_sky130_fd_sc_hd__and2_2 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "0001")
* sky130_fd_sc_hd__clkbuf_16 (A)
.model d_lut_sky130_fd_sc_hd__clkbuf_16 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "01")
* sky130_fd_sc_hd__o21bai_1 (!A1&!A2) | (B1_N)
.model d_lut_sky130_fd_sc_hd__o21bai_1 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "10001111")
* sky130_fd_sc_hd__mux2_1 (A0&!S) | (A1&S)
.model d_lut_sky130_fd_sc_hd__mux2_1 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "01010011")
* sky130_fd_sc_hd__nand2b_1 (A_N) | (!B)
.model d_lut_sky130_fd_sc_hd__nand2b_1 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "1101")
* sky130_fd_sc_hd__and3b_1 (!A_N&B&C)
.model d_lut_sky130_fd_sc_hd__and3b_1 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "00000010")
.end
