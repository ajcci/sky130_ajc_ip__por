xspice/por_dig.out.spice