* NGSPICE file created from por_dig.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

.subckt por_dig VGND VPWR force_pdn force_pdnb force_rc_osc force_short_oneshot osc_ck
+ osc_ck_256 osc_ena otrip[0] otrip[1] otrip[2] otrip_decoded[0] otrip_decoded[1]
+ otrip_decoded[2] otrip_decoded[3] otrip_decoded[4] otrip_decoded[5] otrip_decoded[6]
+ otrip_decoded[7] por_timed_out por_unbuf pwup_filt startup_timed_out
XFILLER_0_2_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_229__29 VGND VGND VPWR VPWR net29 _229__29/LO sky130_fd_sc_hd__conb_1
XFILLER_0_18_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_131_ cnt_ck_256\[6\] _045_ VGND VGND VPWR VPWR _047_ sky130_fd_sc_hd__nand2_1
X_200_ clknet_2_2__leaf_osc_ck _010_ net25 VGND VGND VPWR VPWR cnt_st\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_5_56 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_114_ cnt_st\[1\] cnt_st\[0\] cnt_st\[3\] cnt_st\[2\] VGND VGND VPWR VPWR _037_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_20_87 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_76 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput20 net24 VGND VGND VPWR VPWR por_unbuf sky130_fd_sc_hd__buf_2
XFILLER_0_13_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_21_Right_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_130_ _045_ _046_ VGND VGND VPWR VPWR _005_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_12_Right_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_5_57 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_113_ cnt_st\[1\] cnt_st\[0\] cnt_st\[2\] VGND VGND VPWR VPWR _036_ sky130_fd_sc_hd__and3_1
Xclkbuf_2_3__f_osc_ck clknet_0_osc_ck VGND VGND VPWR VPWR clknet_2_3__leaf_osc_ck
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_21_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_107 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold20 cnt_st\[2\] VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_16_Left_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_15_77 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput10 net10 VGND VGND VPWR VPWR osc_ena sky130_fd_sc_hd__buf_2
Xoutput8 net8 VGND VGND VPWR VPWR force_pdnb sky130_fd_sc_hd__buf_2
Xoutput21 net21 VGND VGND VPWR VPWR startup_timed_out sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_19_Left_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_4_Left_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_189_ net47 _082_ _083_ VGND VGND VPWR VPWR _027_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_10_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_112_ cnt_st\[1\] cnt_st\[0\] VGND VGND VPWR VPWR _035_ sky130_fd_sc_hd__nand2_1
XFILLER_0_21_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold10 cnt_ck_256\[5\] VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__dlygate4sd3_1
Xhold21 cnt_st\[4\] VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput11 net11 VGND VGND VPWR VPWR otrip_decoded[0] sky130_fd_sc_hd__clkbuf_4
Xoutput9 net9 VGND VGND VPWR VPWR osc_ck_256 sky130_fd_sc_hd__buf_2
XFILLER_0_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_20_Left_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_188_ cnt_por\[9\] cnt_por\[10\] net23 _080_ VGND VGND VPWR VPWR _083_ sky130_fd_sc_hd__and4_1
XFILLER_0_10_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_111_ _087_ net19 net2 VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__o21bai_1
Xhold11 cnt_ck_256\[1\] VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__dlygate4sd3_1
Xhold22 cnt_por\[9\] VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__dlygate4sd3_1
Xoutput12 net12 VGND VGND VPWR VPWR otrip_decoded[1] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_5_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_187_ _081_ _082_ VGND VGND VPWR VPWR _026_ sky130_fd_sc_hd__nor2_1
XFILLER_0_10_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_110_ cnt_por\[12\] cnt_por\[13\] _032_ VGND VGND VPWR VPWR _034_ sky130_fd_sc_hd__and3_1
Xhold12 cnt_por\[11\] VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__dlygate4sd3_1
Xhold23 cnt_por\[3\] VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__dlygate4sd3_1
Xoutput13 net13 VGND VGND VPWR VPWR otrip_decoded[2] sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_21_90 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_19_Right_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_186_ cnt_por\[9\] net23 _080_ VGND VGND VPWR VPWR _082_ sky130_fd_sc_hd__and3_1
XFILLER_0_19_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_169_ _069_ _070_ _063_ VGND VGND VPWR VPWR _020_ sky130_fd_sc_hd__a21o_1
Xhold13 cnt_ck_256\[3\] VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__dlygate4sd3_1
Xhold24 cnt_por\[7\] VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_18_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_91 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput14 net14 VGND VGND VPWR VPWR otrip_decoded[3] sky130_fd_sc_hd__buf_2
XFILLER_0_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_185_ net23 _080_ net51 VGND VGND VPWR VPWR _081_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_10_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_099_ net5 net4 net6 VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__nor3b_1
X_168_ _088_ net22 VGND VGND VPWR VPWR _070_ sky130_fd_sc_hd__nand2_1
Xhold14 cnt_por\[8\] VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__dlygate4sd3_1
Xhold25 cnt_por\[4\] VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_11_Left_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_115 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput15 net15 VGND VGND VPWR VPWR otrip_decoded[4] sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_184_ net3 _091_ VGND VGND VPWR VPWR _080_ sky130_fd_sc_hd__or2_1
XFILLER_0_21_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_098_ net6 net5 net4 VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__and3b_1
X_167_ cnt_por\[0\] cnt_por\[1\] cnt_por\[2\] net22 net52 VGND VGND VPWR VPWR _069_
+ sky130_fd_sc_hd__a41o_1
XFILLER_0_1_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold15 cnt_por\[12\] VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_219_ clknet_2_3__leaf_osc_ck _022_ net28 VGND VGND VPWR VPWR cnt_por\[5\] sky130_fd_sc_hd__dfrtp_1
Xoutput16 net16 VGND VGND VPWR VPWR otrip_decoded[5] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_7_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_15_Right_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_3_52 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_116 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_72 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_183_ net43 _078_ _079_ _063_ VGND VGND VPWR VPWR _025_ sky130_fd_sc_hd__a211o_1
XFILLER_0_21_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_097_ net6 net4 net5 VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__nor3b_1
XFILLER_0_11_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_166_ _067_ _068_ _063_ VGND VGND VPWR VPWR _019_ sky130_fd_sc_hd__a21o_1
XFILLER_0_15_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold16 cnt_st\[0\] VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__dlygate4sd3_1
X_218_ clknet_2_3__leaf_osc_ck _021_ net28 VGND VGND VPWR VPWR cnt_por\[4\] sky130_fd_sc_hd__dfrtp_1
X_149_ cnt_st\[6\] _054_ VGND VGND VPWR VPWR _058_ sky130_fd_sc_hd__or2_1
Xoutput17 net17 VGND VGND VPWR VPWR otrip_decoded[6] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_7_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_53 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_13_73 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_182_ cnt_por\[8\] _089_ _090_ net24 VGND VGND VPWR VPWR _079_ sky130_fd_sc_hd__and4b_1
XFILLER_0_21_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_096_ net6 net5 net4 VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__nor3b_1
XFILLER_0_1_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_165_ cnt_por\[0\] cnt_por\[1\] net22 cnt_por\[2\] VGND VGND VPWR VPWR _068_ sky130_fd_sc_hd__a31o_1
Xhold17 cnt_st\[8\] VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_217_ clknet_2_2__leaf_osc_ck _020_ net27 VGND VGND VPWR VPWR cnt_por\[3\] sky130_fd_sc_hd__dfrtp_1
X_148_ cnt_st\[6\] _054_ VGND VGND VPWR VPWR _057_ sky130_fd_sc_hd__nand2_1
XFILLER_0_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput18 net18 VGND VGND VPWR VPWR otrip_decoded[7] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_4_104 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_15_Left_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_2_2__f_osc_ck clknet_0_osc_ck VGND VGND VPWR VPWR clknet_2_2__leaf_osc_ck
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_19_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_18_Left_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_44 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_181_ _077_ _078_ _063_ VGND VGND VPWR VPWR _024_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_9_64 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_3_Left_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_095_ net6 net5 net4 VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__nor3_1
X_164_ cnt_por\[0\] cnt_por\[1\] cnt_por\[2\] net22 VGND VGND VPWR VPWR _067_ sky130_fd_sc_hd__nand4_1
Xhold18 cnt_por\[10\] VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_19_84 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_216_ clknet_2_3__leaf_osc_ck _019_ net27 VGND VGND VPWR VPWR cnt_por\[2\] sky130_fd_sc_hd__dfrtp_1
X_147_ _055_ _056_ net21 VGND VGND VPWR VPWR _012_ sky130_fd_sc_hd__a21o_1
Xoutput19 net19 VGND VGND VPWR VPWR por_timed_out sky130_fd_sc_hd__buf_2
XFILLER_0_4_116 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_20_Right_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_180_ _089_ _090_ net24 VGND VGND VPWR VPWR _078_ sky130_fd_sc_hd__nand3_1
XFILLER_0_19_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_45 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_65 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_094_ net35 VGND VGND VPWR VPWR _000_ sky130_fd_sc_hd__inv_2
X_163_ _065_ _066_ _064_ VGND VGND VPWR VPWR _018_ sky130_fd_sc_hd__o21ai_1
Xhold19 cnt_st\[3\] VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_19_85 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_146_ net3 cnt_st\[5\] _038_ VGND VGND VPWR VPWR _056_ sky130_fd_sc_hd__or3_1
X_215_ clknet_2_3__leaf_osc_ck _018_ net28 VGND VGND VPWR VPWR cnt_por\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_7_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_129_ net38 _043_ net39 VGND VGND VPWR VPWR _046_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_17_94 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout22 net23 VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_0_46 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_231_ clknet_2_1__leaf_osc_ck net31 net7 VGND VGND VPWR VPWR cnt_rsb sky130_fd_sc_hd__dfrtp_1
X_093_ net7 VGND VGND VPWR VPWR _087_ sky130_fd_sc_hd__inv_2
X_162_ cnt_por\[0\] cnt_por\[1\] net22 VGND VGND VPWR VPWR _066_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_10_66 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput1 force_pdn VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__clkbuf_1
X_214_ clknet_2_2__leaf_osc_ck _017_ net27 VGND VGND VPWR VPWR cnt_por\[0\] sky130_fd_sc_hd__dfrtp_2
X_145_ _054_ VGND VGND VPWR VPWR _055_ sky130_fd_sc_hd__inv_2
X_128_ cnt_ck_256\[4\] cnt_ck_256\[5\] _043_ VGND VGND VPWR VPWR _045_ sky130_fd_sc_hd__and3_1
XFILLER_0_17_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_47 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout23 net24 VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__clkbuf_2
X_230_ clknet_2_1__leaf_osc_ck net32 net7 VGND VGND VPWR VPWR cnt_rsb_stg2 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_161_ cnt_por\[0\] net22 cnt_por\[1\] VGND VGND VPWR VPWR _065_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_1_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_092_ net1 VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__inv_2
Xinput2 force_rc_osc VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_7_Left_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_67 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_213_ clknet_2_1__leaf_osc_ck _016_ net27 VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__dfrtp_1
X_144_ net3 _038_ cnt_st\[5\] VGND VGND VPWR VPWR _054_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_21_88 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_127_ net38 _043_ VGND VGND VPWR VPWR _004_ sky130_fd_sc_hd__xor2_1
XFILLER_0_0_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout24 net20 VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__clkbuf_2
X_160_ net3 net22 VGND VGND VPWR VPWR _064_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_18_Right_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput3 force_short_oneshot VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__clkbuf_2
X_212_ clknet_2_1__leaf_osc_ck _006_ net27 VGND VGND VPWR VPWR cnt_ck_256\[6\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_6_58 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_143_ _038_ _053_ _049_ VGND VGND VPWR VPWR _011_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_21_89 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_126_ _043_ _044_ VGND VGND VPWR VPWR _003_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_10_Left_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_16_78 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_109_ _091_ _033_ VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__and2_1
Xfanout25 net26 VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_1_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput4 otrip[0] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__dlymetal6s2s_1
X_211_ clknet_2_1__leaf_osc_ck _005_ net27 VGND VGND VPWR VPWR cnt_ck_256\[5\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_6_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_142_ net50 _037_ VGND VGND VPWR VPWR _053_ sky130_fd_sc_hd__nor2_1
X_125_ net42 _041_ VGND VGND VPWR VPWR _044_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_16_79 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_108_ cnt_por\[12\] cnt_por\[13\] cnt_por\[14\] _032_ VGND VGND VPWR VPWR _033_ sky130_fd_sc_hd__and4_1
XFILLER_0_14_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout26 net30 VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__buf_2
XFILLER_0_5_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput5 otrip[1] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__dlymetal6s2s_1
X_210_ clknet_2_0__leaf_osc_ck _004_ net25 VGND VGND VPWR VPWR cnt_ck_256\[4\] sky130_fd_sc_hd__dfrtp_1
X_141_ _037_ _052_ _049_ VGND VGND VPWR VPWR _010_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_11_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_124_ cnt_ck_256\[3\] _041_ VGND VGND VPWR VPWR _043_ sky130_fd_sc_hd__and2_1
XFILLER_0_17_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_107_ cnt_por\[9\] cnt_por\[10\] cnt_por\[11\] VGND VGND VPWR VPWR _032_ sky130_fd_sc_hd__and3_1
Xfanout27 net30 VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_18_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput6 otrip[2] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__dlymetal6s2s_1
X_140_ net48 _036_ VGND VGND VPWR VPWR _052_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_14_Right_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_123_ _041_ net37 VGND VGND VPWR VPWR _002_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_7_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_106_ cnt_por\[4\] cnt_por\[8\] _088_ _090_ VGND VGND VPWR VPWR _091_ sky130_fd_sc_hd__and4_1
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_14_Left_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_17_80 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout28 net30 VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput7 pwup_filt VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__dlymetal6s2s_1
XPHY_EDGE_ROW_2_Left_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_199_ clknet_2_0__leaf_osc_ck _009_ net25 VGND VGND VPWR VPWR cnt_st\[2\] sky130_fd_sc_hd__dfrtp_1
X_122_ cnt_ck_256\[1\] cnt_ck_256\[0\] net36 VGND VGND VPWR VPWR _042_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_7_61 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_2_1__f_osc_ck clknet_0_osc_ck VGND VGND VPWR VPWR clknet_2_1__leaf_osc_ck
+ sky130_fd_sc_hd__clkbuf_16
X_105_ cnt_por\[5\] cnt_por\[6\] cnt_por\[7\] VGND VGND VPWR VPWR _090_ sky130_fd_sc_hd__and3_1
XFILLER_0_8_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_17_81 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_198_ clknet_2_0__leaf_osc_ck _008_ net25 VGND VGND VPWR VPWR cnt_st\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_121_ cnt_ck_256\[1\] cnt_ck_256\[0\] cnt_ck_256\[2\] VGND VGND VPWR VPWR _041_ sky130_fd_sc_hd__and3_1
XFILLER_0_17_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_104_ cnt_por\[4\] _088_ VGND VGND VPWR VPWR _089_ sky130_fd_sc_hd__and2_2
XFILLER_0_5_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_197_ clknet_2_0__leaf_osc_ck _007_ net25 VGND VGND VPWR VPWR cnt_st\[0\] sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_120_ net40 net35 VGND VGND VPWR VPWR _001_ sky130_fd_sc_hd__xor2_1
XFILLER_0_17_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_103_ cnt_por\[0\] cnt_por\[1\] cnt_por\[2\] cnt_por\[3\] VGND VGND VPWR VPWR _088_
+ sky130_fd_sc_hd__and4_1
Xhold1 cnt_rsb VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_196_ net34 _085_ VGND VGND VPWR VPWR _031_ sky130_fd_sc_hd__xor2_1
XPHY_EDGE_ROW_6_Left_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_179_ cnt_por\[5\] cnt_por\[6\] _089_ net24 net53 VGND VGND VPWR VPWR _077_ sky130_fd_sc_hd__a41o_1
XFILLER_0_17_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_102_ net6 net5 net4 VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__and3_1
Xclkbuf_0_osc_ck osc_ck VGND VGND VPWR VPWR clknet_0_osc_ck sky130_fd_sc_hd__clkbuf_16
XFILLER_0_19_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_9_Left_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_4_54 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2 cnt_rsb_stg2 VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_17_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_74 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_195_ _085_ _086_ VGND VGND VPWR VPWR _030_ sky130_fd_sc_hd__and2b_1
XFILLER_0_11_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_178_ _075_ _076_ _063_ VGND VGND VPWR VPWR _023_ sky130_fd_sc_hd__a21o_1
X_101_ net4 net5 net6 VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_4_55 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3 cnt_rsb_stg1 VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_75 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_194_ cnt_por\[12\] _032_ net23 _080_ cnt_por\[13\] VGND VGND VPWR VPWR _086_ sky130_fd_sc_hd__a41o_1
X_177_ cnt_por\[5\] cnt_por\[6\] _089_ net24 VGND VGND VPWR VPWR _076_ sky130_fd_sc_hd__nand4_1
X_100_ net5 net4 net6 VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__and3b_1
X_229_ clknet_2_1__leaf_osc_ck net29 net7 VGND VGND VPWR VPWR cnt_rsb_stg1 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold4 net9 VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_17_Right_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_193_ _034_ net23 _080_ VGND VGND VPWR VPWR _085_ sky130_fd_sc_hd__and3_1
XFILLER_0_6_105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_176_ cnt_por\[5\] _089_ net24 cnt_por\[6\] VGND VGND VPWR VPWR _075_ sky130_fd_sc_hd__a31o_1
X_228_ clknet_2_0__leaf_osc_ck _031_ net26 VGND VGND VPWR VPWR cnt_por\[14\] sky130_fd_sc_hd__dfrtp_1
X_159_ net3 net22 VGND VGND VPWR VPWR _063_ sky130_fd_sc_hd__and2_1
XFILLER_0_20_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold5 cnt_por\[14\] VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_17_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_192_ net44 _084_ VGND VGND VPWR VPWR _029_ sky130_fd_sc_hd__xor2_1
XFILLER_0_6_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_175_ _073_ _074_ _064_ VGND VGND VPWR VPWR _022_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_18_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_227_ clknet_2_0__leaf_osc_ck _030_ net25 VGND VGND VPWR VPWR cnt_por\[13\] sky130_fd_sc_hd__dfrtp_1
X_158_ cnt_por\[0\] net22 _062_ VGND VGND VPWR VPWR _017_ sky130_fd_sc_hd__o21a_1
XFILLER_0_20_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold6 cnt_ck_256\[0\] VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_13_Left_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_1_48 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_191_ net41 _083_ _084_ VGND VGND VPWR VPWR _028_ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_11_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_1_Left_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_174_ cnt_por\[5\] _089_ net24 VGND VGND VPWR VPWR _074_ sky130_fd_sc_hd__and3_1
XFILLER_0_3_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_226_ clknet_2_0__leaf_osc_ck _029_ net27 VGND VGND VPWR VPWR cnt_por\[12\] sky130_fd_sc_hd__dfrtp_1
X_157_ net3 cnt_por\[0\] net22 VGND VGND VPWR VPWR _062_ sky130_fd_sc_hd__nand3b_1
Xhold7 cnt_ck_256\[2\] VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_209_ clknet_2_1__leaf_osc_ck _003_ net25 VGND VGND VPWR VPWR cnt_ck_256\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_13_Right_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_1_49 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_2_0__f_osc_ck clknet_0_osc_ck VGND VGND VPWR VPWR clknet_2_0__leaf_osc_ck
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_6_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_190_ _032_ net23 _080_ VGND VGND VPWR VPWR _084_ sky130_fd_sc_hd__and3_1
XFILLER_0_10_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_11_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_173_ _089_ net24 cnt_por\[5\] VGND VGND VPWR VPWR _073_ sky130_fd_sc_hd__a21oi_1
X_156_ net33 _047_ VGND VGND VPWR VPWR _016_ sky130_fd_sc_hd__xnor2_1
X_225_ clknet_2_1__leaf_osc_ck _028_ net27 VGND VGND VPWR VPWR cnt_por\[11\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold8 _042_ VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_208_ clknet_2_0__leaf_osc_ck _002_ net25 VGND VGND VPWR VPWR cnt_ck_256\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_139_ _036_ _051_ _049_ VGND VGND VPWR VPWR _009_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_172_ _071_ _072_ _063_ VGND VGND VPWR VPWR _021_ sky130_fd_sc_hd__a21o_1
X_224_ clknet_2_1__leaf_osc_ck _027_ net27 VGND VGND VPWR VPWR cnt_por\[10\] sky130_fd_sc_hd__dfrtp_1
X_155_ _040_ _061_ VGND VGND VPWR VPWR _015_ sky130_fd_sc_hd__nand2_1
XFILLER_0_18_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold9 cnt_ck_256\[4\] VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__dlygate4sd3_1
X_207_ clknet_2_0__leaf_osc_ck _001_ net25 VGND VGND VPWR VPWR cnt_ck_256\[1\] sky130_fd_sc_hd__dfrtp_1
X_138_ cnt_st\[1\] cnt_st\[0\] net49 VGND VGND VPWR VPWR _051_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_0_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_17_Left_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_2_50 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_171_ _088_ net23 net54 VGND VGND VPWR VPWR _072_ sky130_fd_sc_hd__a21o_1
XFILLER_0_3_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_5_Left_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_223_ clknet_2_1__leaf_osc_ck _026_ net27 VGND VGND VPWR VPWR cnt_por\[9\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_12_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_154_ net46 _060_ VGND VGND VPWR VPWR _061_ sky130_fd_sc_hd__xor2_1
X_206_ clknet_2_0__leaf_osc_ck _000_ net25 VGND VGND VPWR VPWR cnt_ck_256\[0\] sky130_fd_sc_hd__dfrtp_1
X_137_ _035_ _050_ net21 net3 VGND VGND VPWR VPWR _008_ sky130_fd_sc_hd__a211o_1
XFILLER_0_9_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_8_Left_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_51 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_170_ _089_ net23 VGND VGND VPWR VPWR _071_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_21_Left_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_12_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_222_ clknet_2_3__leaf_osc_ck _025_ net28 VGND VGND VPWR VPWR cnt_por\[8\] sky130_fd_sc_hd__dfrtp_1
X_153_ _040_ _059_ _060_ net21 VGND VGND VPWR VPWR _014_ sky130_fd_sc_hd__a31o_1
X_136_ cnt_st\[1\] cnt_st\[0\] VGND VGND VPWR VPWR _050_ sky130_fd_sc_hd__or2_1
X_205_ clknet_2_2__leaf_osc_ck _015_ net26 VGND VGND VPWR VPWR cnt_st\[8\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_119_ _091_ _033_ net21 VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__a21boi_1
XFILLER_0_6_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_8_62 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_152_ net3 _039_ VGND VGND VPWR VPWR _060_ sky130_fd_sc_hd__nand2_1
X_221_ clknet_2_3__leaf_osc_ck _024_ net28 VGND VGND VPWR VPWR cnt_por\[7\] sky130_fd_sc_hd__dfrtp_1
X_204_ clknet_2_2__leaf_osc_ck _014_ net26 VGND VGND VPWR VPWR cnt_st\[7\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_135_ net45 _049_ VGND VGND VPWR VPWR _007_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_18_82 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_118_ cnt_st\[8\] cnt_st\[4\] _037_ _039_ VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__and4_2
XFILLER_0_8_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_151_ cnt_st\[6\] _054_ cnt_st\[7\] VGND VGND VPWR VPWR _059_ sky130_fd_sc_hd__a21o_1
X_220_ clknet_2_3__leaf_osc_ck _023_ net28 VGND VGND VPWR VPWR cnt_por\[6\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_8_63 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_134_ net3 net21 VGND VGND VPWR VPWR _049_ sky130_fd_sc_hd__nor2_1
X_203_ clknet_2_2__leaf_osc_ck _013_ net26 VGND VGND VPWR VPWR cnt_st\[6\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_83 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_117_ _038_ _039_ VGND VGND VPWR VPWR _040_ sky130_fd_sc_hd__nand2_1
XFILLER_0_15_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_150_ _057_ _058_ net21 VGND VGND VPWR VPWR _013_ sky130_fd_sc_hd__a21o_1
XFILLER_0_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_16_Right_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_133_ _047_ _048_ VGND VGND VPWR VPWR _006_ sky130_fd_sc_hd__and2_1
X_202_ clknet_2_2__leaf_osc_ck _012_ net26 VGND VGND VPWR VPWR cnt_st\[5\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_12_Left_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_116_ cnt_st\[6\] cnt_st\[7\] cnt_st\[5\] VGND VGND VPWR VPWR _039_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_0_Left_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_132_ cnt_ck_256\[6\] _045_ VGND VGND VPWR VPWR _048_ sky130_fd_sc_hd__or2_1
X_201_ clknet_2_2__leaf_osc_ck _011_ net26 VGND VGND VPWR VPWR cnt_st\[4\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_115_ cnt_st\[4\] _037_ VGND VGND VPWR VPWR _038_ sky130_fd_sc_hd__and2_1
XFILLER_0_21_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_86 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
.ends

