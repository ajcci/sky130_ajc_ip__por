magic
tech sky130A
magscale 1 2
timestamp 1712975145
<< pwell >>
rect -2008 -11682 2008 11682
<< psubdiff >>
rect -1972 11612 -1876 11646
rect 1876 11612 1972 11646
rect -1972 11550 -1938 11612
rect 1938 11550 1972 11612
rect -1972 -11612 -1938 -11550
rect 1938 -11612 1972 -11550
rect -1972 -11646 -1876 -11612
rect 1876 -11646 1972 -11612
<< psubdiffcont >>
rect -1876 11612 1876 11646
rect -1972 -11550 -1938 11550
rect 1938 -11550 1972 11550
rect -1876 -11646 1876 -11612
<< xpolycontact >>
rect -1842 11084 -1560 11516
rect -1842 -11516 -1560 -11084
rect -1464 11084 -1182 11516
rect -1464 -11516 -1182 -11084
rect -1086 11084 -804 11516
rect -1086 -11516 -804 -11084
rect -708 11084 -426 11516
rect -708 -11516 -426 -11084
rect -330 11084 -48 11516
rect -330 -11516 -48 -11084
rect 48 11084 330 11516
rect 48 -11516 330 -11084
rect 426 11084 708 11516
rect 426 -11516 708 -11084
rect 804 11084 1086 11516
rect 804 -11516 1086 -11084
rect 1182 11084 1464 11516
rect 1182 -11516 1464 -11084
rect 1560 11084 1842 11516
rect 1560 -11516 1842 -11084
<< xpolyres >>
rect -1842 -11084 -1560 11084
rect -1464 -11084 -1182 11084
rect -1086 -11084 -804 11084
rect -708 -11084 -426 11084
rect -330 -11084 -48 11084
rect 48 -11084 330 11084
rect 426 -11084 708 11084
rect 804 -11084 1086 11084
rect 1182 -11084 1464 11084
rect 1560 -11084 1842 11084
<< locali >>
rect -1972 11612 -1876 11646
rect 1876 11612 1972 11646
rect -1972 11550 -1938 11612
rect 1938 11550 1972 11612
rect -1972 -11612 -1938 -11550
rect 1938 -11612 1972 -11550
rect -1972 -11646 -1876 -11612
rect 1876 -11646 1972 -11612
<< viali >>
rect -1826 11101 -1576 11498
rect -1448 11101 -1198 11498
rect -1070 11101 -820 11498
rect -692 11101 -442 11498
rect -314 11101 -64 11498
rect 64 11101 314 11498
rect 442 11101 692 11498
rect 820 11101 1070 11498
rect 1198 11101 1448 11498
rect 1576 11101 1826 11498
rect -1826 -11498 -1576 -11101
rect -1448 -11498 -1198 -11101
rect -1070 -11498 -820 -11101
rect -692 -11498 -442 -11101
rect -314 -11498 -64 -11101
rect 64 -11498 314 -11101
rect 442 -11498 692 -11101
rect 820 -11498 1070 -11101
rect 1198 -11498 1448 -11101
rect 1576 -11498 1826 -11101
<< metal1 >>
rect -1832 11498 -1570 11510
rect -1832 11101 -1826 11498
rect -1576 11101 -1570 11498
rect -1832 11089 -1570 11101
rect -1454 11498 -1192 11510
rect -1454 11101 -1448 11498
rect -1198 11101 -1192 11498
rect -1454 11089 -1192 11101
rect -1076 11498 -814 11510
rect -1076 11101 -1070 11498
rect -820 11101 -814 11498
rect -1076 11089 -814 11101
rect -698 11498 -436 11510
rect -698 11101 -692 11498
rect -442 11101 -436 11498
rect -698 11089 -436 11101
rect -320 11498 -58 11510
rect -320 11101 -314 11498
rect -64 11101 -58 11498
rect -320 11089 -58 11101
rect 58 11498 320 11510
rect 58 11101 64 11498
rect 314 11101 320 11498
rect 58 11089 320 11101
rect 436 11498 698 11510
rect 436 11101 442 11498
rect 692 11101 698 11498
rect 436 11089 698 11101
rect 814 11498 1076 11510
rect 814 11101 820 11498
rect 1070 11101 1076 11498
rect 814 11089 1076 11101
rect 1192 11498 1454 11510
rect 1192 11101 1198 11498
rect 1448 11101 1454 11498
rect 1192 11089 1454 11101
rect 1570 11498 1832 11510
rect 1570 11101 1576 11498
rect 1826 11101 1832 11498
rect 1570 11089 1832 11101
rect -1832 -11101 -1570 -11089
rect -1832 -11498 -1826 -11101
rect -1576 -11498 -1570 -11101
rect -1832 -11510 -1570 -11498
rect -1454 -11101 -1192 -11089
rect -1454 -11498 -1448 -11101
rect -1198 -11498 -1192 -11101
rect -1454 -11510 -1192 -11498
rect -1076 -11101 -814 -11089
rect -1076 -11498 -1070 -11101
rect -820 -11498 -814 -11101
rect -1076 -11510 -814 -11498
rect -698 -11101 -436 -11089
rect -698 -11498 -692 -11101
rect -442 -11498 -436 -11101
rect -698 -11510 -436 -11498
rect -320 -11101 -58 -11089
rect -320 -11498 -314 -11101
rect -64 -11498 -58 -11101
rect -320 -11510 -58 -11498
rect 58 -11101 320 -11089
rect 58 -11498 64 -11101
rect 314 -11498 320 -11101
rect 58 -11510 320 -11498
rect 436 -11101 698 -11089
rect 436 -11498 442 -11101
rect 692 -11498 698 -11101
rect 436 -11510 698 -11498
rect 814 -11101 1076 -11089
rect 814 -11498 820 -11101
rect 1070 -11498 1076 -11101
rect 814 -11510 1076 -11498
rect 1192 -11101 1454 -11089
rect 1192 -11498 1198 -11101
rect 1448 -11498 1454 -11101
rect 1192 -11510 1454 -11498
rect 1570 -11101 1832 -11089
rect 1570 -11498 1576 -11101
rect 1826 -11498 1832 -11101
rect 1570 -11510 1832 -11498
<< properties >>
string FIXED_BBOX -1955 -11629 1955 11629
string gencell sky130_fd_pr__res_xhigh_po_1p41
string library sky130
string parameters w 1.410 l 111 m 1 nx 10 wmin 1.410 lmin 0.50 rho 2000 val 157.713k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 1.410 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
