magic
tech sky130A
magscale 1 2
timestamp 1713190415
<< viali >>
rect 6009 11305 6043 11339
rect 5641 11237 5675 11271
rect 4721 11101 4755 11135
rect 4997 11101 5031 11135
rect 5089 11101 5123 11135
rect 5365 11101 5399 11135
rect 6193 11101 6227 11135
rect 6929 11101 6963 11135
rect 4905 11033 4939 11067
rect 5457 11033 5491 11067
rect 5641 11033 5675 11067
rect 5273 10965 5307 10999
rect 6377 10965 6411 10999
rect 5917 10761 5951 10795
rect 2329 10625 2363 10659
rect 4169 10625 4203 10659
rect 6193 10625 6227 10659
rect 2605 10557 2639 10591
rect 4445 10557 4479 10591
rect 6377 10557 6411 10591
rect 6653 10557 6687 10591
rect 8769 10557 8803 10591
rect 4077 10421 4111 10455
rect 6101 10421 6135 10455
rect 8125 10421 8159 10455
rect 8217 10421 8251 10455
rect 4813 10217 4847 10251
rect 5365 10217 5399 10251
rect 1869 10081 1903 10115
rect 3617 10081 3651 10115
rect 5457 10081 5491 10115
rect 6193 10081 6227 10115
rect 8033 10081 8067 10115
rect 4445 10013 4479 10047
rect 4938 10013 4972 10047
rect 5733 10013 5767 10047
rect 8493 10013 8527 10047
rect 8677 10013 8711 10047
rect 2145 9945 2179 9979
rect 5917 9945 5951 9979
rect 6469 9945 6503 9979
rect 8217 9945 8251 9979
rect 8401 9945 8435 9979
rect 3801 9877 3835 9911
rect 4997 9877 5031 9911
rect 5549 9877 5583 9911
rect 7941 9877 7975 9911
rect 8493 9877 8527 9911
rect 6561 9673 6595 9707
rect 6929 9673 6963 9707
rect 7389 9673 7423 9707
rect 3249 9605 3283 9639
rect 7021 9605 7055 9639
rect 7665 9605 7699 9639
rect 7875 9605 7909 9639
rect 8309 9605 8343 9639
rect 2145 9537 2179 9571
rect 3341 9537 3375 9571
rect 3433 9537 3467 9571
rect 4077 9537 4111 9571
rect 4813 9537 4847 9571
rect 4997 9537 5031 9571
rect 5181 9537 5215 9571
rect 5365 9535 5399 9569
rect 5641 9537 5675 9571
rect 5825 9537 5859 9571
rect 7573 9537 7607 9571
rect 7758 9537 7792 9571
rect 8401 9537 8435 9571
rect 8493 9537 8527 9571
rect 1777 9469 1811 9503
rect 2237 9469 2271 9503
rect 2421 9469 2455 9503
rect 3985 9469 4019 9503
rect 4445 9469 4479 9503
rect 5549 9469 5583 9503
rect 7205 9469 7239 9503
rect 8033 9469 8067 9503
rect 2697 9401 2731 9435
rect 3617 9401 3651 9435
rect 6009 9401 6043 9435
rect 8677 9401 8711 9435
rect 2881 9333 2915 9367
rect 3065 9333 3099 9367
rect 4537 9333 4571 9367
rect 4813 9333 4847 9367
rect 8125 9333 8159 9367
rect 2893 9129 2927 9163
rect 4721 9129 4755 9163
rect 5549 9129 5583 9163
rect 7665 9129 7699 9163
rect 5733 9061 5767 9095
rect 5917 9061 5951 9095
rect 3157 8993 3191 9027
rect 3985 8993 4019 9027
rect 5181 8993 5215 9027
rect 7021 8993 7055 9027
rect 3617 8925 3651 8959
rect 4077 8925 4111 8959
rect 4445 8925 4479 8959
rect 4721 8925 4755 8959
rect 5089 8925 5123 8959
rect 5825 8925 5859 8959
rect 6101 8925 6135 8959
rect 6377 8925 6411 8959
rect 6561 8925 6595 8959
rect 6653 8925 6687 8959
rect 6745 8925 6779 8959
rect 7297 8925 7331 8959
rect 7481 8925 7515 8959
rect 7757 8925 7791 8959
rect 8033 8925 8067 8959
rect 1409 8789 1443 8823
rect 3433 8789 3467 8823
rect 3801 8789 3835 8823
rect 4261 8789 4295 8823
rect 4353 8789 4387 8823
rect 4537 8789 4571 8823
rect 5549 8789 5583 8823
rect 7113 8789 7147 8823
rect 8585 8789 8619 8823
rect 2697 8585 2731 8619
rect 3065 8585 3099 8619
rect 3249 8585 3283 8619
rect 4445 8585 4479 8619
rect 6745 8585 6779 8619
rect 9045 8585 9079 8619
rect 1501 8449 1535 8483
rect 1685 8449 1719 8483
rect 2973 8449 3007 8483
rect 3341 8449 3375 8483
rect 3893 8449 3927 8483
rect 4261 8449 4295 8483
rect 4997 8449 5031 8483
rect 5089 8449 5123 8483
rect 5457 8449 5491 8483
rect 6101 8449 6135 8483
rect 6377 8449 6411 8483
rect 6561 8449 6595 8483
rect 8493 8449 8527 8483
rect 8677 8449 8711 8483
rect 9048 8449 9082 8483
rect 1961 8381 1995 8415
rect 2605 8381 2639 8415
rect 2881 8381 2915 8415
rect 3801 8381 3835 8415
rect 5181 8381 5215 8415
rect 5273 8381 5307 8415
rect 5549 8381 5583 8415
rect 8217 8381 8251 8415
rect 8585 8381 8619 8415
rect 1869 8313 1903 8347
rect 6469 8313 6503 8347
rect 9229 8313 9263 8347
rect 4261 8245 4295 8279
rect 4813 8245 4847 8279
rect 2329 8041 2363 8075
rect 2973 7973 3007 8007
rect 8401 7973 8435 8007
rect 1685 7905 1719 7939
rect 2145 7905 2179 7939
rect 6653 7905 6687 7939
rect 9505 7905 9539 7939
rect 1409 7837 1443 7871
rect 2053 7837 2087 7871
rect 2697 7837 2731 7871
rect 3157 7837 3191 7871
rect 3433 7837 3467 7871
rect 3617 7837 3651 7871
rect 3985 7837 4019 7871
rect 4629 7837 4663 7871
rect 4813 7837 4847 7871
rect 2513 7769 2547 7803
rect 2881 7769 2915 7803
rect 4077 7769 4111 7803
rect 6929 7769 6963 7803
rect 1593 7701 1627 7735
rect 2605 7701 2639 7735
rect 3893 7701 3927 7735
rect 6101 7701 6135 7735
rect 8953 7701 8987 7735
rect 1501 7497 1535 7531
rect 1869 7497 1903 7531
rect 2881 7497 2915 7531
rect 6193 7497 6227 7531
rect 6745 7497 6779 7531
rect 9045 7497 9079 7531
rect 4353 7429 4387 7463
rect 4721 7429 4755 7463
rect 7757 7429 7791 7463
rect 1685 7361 1719 7395
rect 4445 7361 4479 7395
rect 6561 7361 6595 7395
rect 6929 7361 6963 7395
rect 7205 7361 7239 7395
rect 7389 7361 7423 7395
rect 7665 7361 7699 7395
rect 2421 7293 2455 7327
rect 6469 7157 6503 7191
rect 7573 7157 7607 7191
rect 1672 6953 1706 6987
rect 5549 6953 5583 6987
rect 5641 6953 5675 6987
rect 6561 6953 6595 6987
rect 7205 6953 7239 6987
rect 7481 6953 7515 6987
rect 6377 6885 6411 6919
rect 8033 6885 8067 6919
rect 8309 6885 8343 6919
rect 1409 6817 1443 6851
rect 3801 6817 3835 6851
rect 4077 6817 4111 6851
rect 8953 6817 8987 6851
rect 3525 6749 3559 6783
rect 5917 6749 5951 6783
rect 6009 6749 6043 6783
rect 6101 6749 6135 6783
rect 6285 6749 6319 6783
rect 6929 6749 6963 6783
rect 8585 6749 8619 6783
rect 9137 6749 9171 6783
rect 7021 6681 7055 6715
rect 7665 6681 7699 6715
rect 9321 6681 9355 6715
rect 3157 6613 3191 6647
rect 3341 6613 3375 6647
rect 6561 6613 6595 6647
rect 7221 6613 7255 6647
rect 7389 6613 7423 6647
rect 7757 6613 7791 6647
rect 7849 6613 7883 6647
rect 8125 6613 8159 6647
rect 4629 6409 4663 6443
rect 6377 6409 6411 6443
rect 3157 6341 3191 6375
rect 4873 6341 4907 6375
rect 5089 6341 5123 6375
rect 7113 6341 7147 6375
rect 1593 6273 1627 6307
rect 1685 6273 1719 6307
rect 1869 6273 1903 6307
rect 2881 6273 2915 6307
rect 5825 6273 5859 6307
rect 6561 6273 6595 6307
rect 7297 6273 7331 6307
rect 7481 6273 7515 6307
rect 7573 6273 7607 6307
rect 7665 6273 7699 6307
rect 8033 6273 8067 6307
rect 8217 6273 8251 6307
rect 1777 6205 1811 6239
rect 2789 6205 2823 6239
rect 6653 6205 6687 6239
rect 2145 6137 2179 6171
rect 4721 6137 4755 6171
rect 7113 6137 7147 6171
rect 2053 6069 2087 6103
rect 4905 6069 4939 6103
rect 5273 6069 5307 6103
rect 7941 6069 7975 6103
rect 8217 6069 8251 6103
rect 1672 5865 1706 5899
rect 3433 5865 3467 5899
rect 3985 5865 4019 5899
rect 4353 5865 4387 5899
rect 7021 5865 7055 5899
rect 8505 5865 8539 5899
rect 1409 5729 1443 5763
rect 3801 5729 3835 5763
rect 4905 5729 4939 5763
rect 6940 5729 6974 5763
rect 8769 5729 8803 5763
rect 3249 5661 3283 5695
rect 3893 5661 3927 5695
rect 4261 5661 4295 5695
rect 10149 5661 10183 5695
rect 6653 5593 6687 5627
rect 3157 5525 3191 5559
rect 4169 5525 4203 5559
rect 5181 5525 5215 5559
rect 9965 5525 9999 5559
rect 1961 5321 1995 5355
rect 6193 5321 6227 5355
rect 6377 5321 6411 5355
rect 1409 5185 1443 5219
rect 1869 5185 1903 5219
rect 2145 5185 2179 5219
rect 2605 5185 2639 5219
rect 4445 5185 4479 5219
rect 6561 5185 6595 5219
rect 6837 5185 6871 5219
rect 7021 5185 7055 5219
rect 8861 5185 8895 5219
rect 2881 5117 2915 5151
rect 4721 5117 4755 5151
rect 7113 5117 7147 5151
rect 8585 5117 8619 5151
rect 1593 5049 1627 5083
rect 4353 5049 4387 5083
rect 6653 5049 6687 5083
rect 6745 5049 6779 5083
rect 2329 4981 2363 5015
rect 3157 4777 3191 4811
rect 3801 4777 3835 4811
rect 3985 4777 4019 4811
rect 5457 4777 5491 4811
rect 6837 4777 6871 4811
rect 8033 4777 8067 4811
rect 6745 4709 6779 4743
rect 1409 4641 1443 4675
rect 4537 4641 4571 4675
rect 6469 4641 6503 4675
rect 6929 4641 6963 4675
rect 7665 4641 7699 4675
rect 4077 4573 4111 4607
rect 4353 4573 4387 4607
rect 5181 4573 5215 4607
rect 5457 4573 5491 4607
rect 5641 4573 5675 4607
rect 6653 4573 6687 4607
rect 7849 4573 7883 4607
rect 1685 4505 1719 4539
rect 5089 4437 5123 4471
rect 5917 4437 5951 4471
rect 7113 4437 7147 4471
rect 1777 4233 1811 4267
rect 4169 4233 4203 4267
rect 5273 4233 5307 4267
rect 4445 4165 4479 4199
rect 5457 4165 5491 4199
rect 1685 4097 1719 4131
rect 2053 4097 2087 4131
rect 5181 4097 5215 4131
rect 5641 4097 5675 4131
rect 7021 4097 7055 4131
rect 2145 4029 2179 4063
rect 7113 4029 7147 4063
rect 7389 4029 7423 4063
rect 1501 3961 1535 3995
rect 5457 3961 5491 3995
rect 5825 3961 5859 3995
rect 1593 3689 1627 3723
rect 5549 3689 5583 3723
rect 6009 3553 6043 3587
rect 1409 3485 1443 3519
rect 3985 3485 4019 3519
rect 4629 3485 4663 3519
rect 6101 3485 6135 3519
rect 5503 3451 5537 3485
rect 5733 3417 5767 3451
rect 5825 3417 5859 3451
rect 4169 3349 4203 3383
rect 4813 3349 4847 3383
rect 5365 3349 5399 3383
rect 6101 3349 6135 3383
rect 3709 3145 3743 3179
rect 4721 3145 4755 3179
rect 6193 3145 6227 3179
rect 6009 3077 6043 3111
rect 6745 3077 6779 3111
rect 4077 3009 4111 3043
rect 4445 3009 4479 3043
rect 4537 3009 4571 3043
rect 4997 3009 5031 3043
rect 6377 3009 6411 3043
rect 3893 2941 3927 2975
rect 3985 2941 4019 2975
rect 4353 2941 4387 2975
rect 5089 2941 5123 2975
rect 5181 2941 5215 2975
rect 5641 2941 5675 2975
rect 4813 2805 4847 2839
rect 6009 2805 6043 2839
rect 6745 2805 6779 2839
rect 6929 2805 6963 2839
rect 6009 2601 6043 2635
rect 5641 2533 5675 2567
rect 2973 2465 3007 2499
rect 4077 2465 4111 2499
rect 9413 2465 9447 2499
rect 2697 2397 2731 2431
rect 3801 2397 3835 2431
rect 4905 2397 4939 2431
rect 5273 2397 5307 2431
rect 6561 2397 6595 2431
rect 7205 2397 7239 2431
rect 7849 2397 7883 2431
rect 8493 2397 8527 2431
rect 9137 2397 9171 2431
rect 6009 2329 6043 2363
rect 5089 2261 5123 2295
rect 5457 2261 5491 2295
rect 6193 2261 6227 2295
rect 6745 2261 6779 2295
rect 7389 2261 7423 2295
rect 8033 2261 8067 2295
rect 8677 2261 8711 2295
<< metal1 >>
rect 1104 11450 10488 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 10488 11450
rect 1104 11376 10488 11398
rect 5810 11296 5816 11348
rect 5868 11336 5874 11348
rect 5997 11339 6055 11345
rect 5997 11336 6009 11339
rect 5868 11308 6009 11336
rect 5868 11296 5874 11308
rect 5997 11305 6009 11308
rect 6043 11305 6055 11339
rect 5997 11299 6055 11305
rect 5626 11228 5632 11280
rect 5684 11228 5690 11280
rect 5810 11200 5816 11212
rect 5092 11172 5816 11200
rect 4706 11092 4712 11144
rect 4764 11092 4770 11144
rect 5092 11141 5120 11172
rect 5810 11160 5816 11172
rect 5868 11160 5874 11212
rect 4985 11135 5043 11141
rect 4985 11132 4997 11135
rect 4816 11104 4997 11132
rect 4246 11024 4252 11076
rect 4304 11064 4310 11076
rect 4816 11064 4844 11104
rect 4985 11101 4997 11104
rect 5031 11101 5043 11135
rect 4985 11095 5043 11101
rect 5077 11135 5135 11141
rect 5077 11101 5089 11135
rect 5123 11101 5135 11135
rect 5077 11095 5135 11101
rect 5353 11135 5411 11141
rect 5353 11101 5365 11135
rect 5399 11132 5411 11135
rect 5534 11132 5540 11144
rect 5399 11104 5540 11132
rect 5399 11101 5411 11104
rect 5353 11095 5411 11101
rect 5534 11092 5540 11104
rect 5592 11092 5598 11144
rect 6086 11092 6092 11144
rect 6144 11132 6150 11144
rect 6181 11135 6239 11141
rect 6181 11132 6193 11135
rect 6144 11104 6193 11132
rect 6144 11092 6150 11104
rect 6181 11101 6193 11104
rect 6227 11101 6239 11135
rect 6181 11095 6239 11101
rect 6917 11135 6975 11141
rect 6917 11101 6929 11135
rect 6963 11101 6975 11135
rect 6917 11095 6975 11101
rect 4304 11036 4844 11064
rect 4304 11024 4310 11036
rect 4890 11024 4896 11076
rect 4948 11024 4954 11076
rect 5442 11024 5448 11076
rect 5500 11024 5506 11076
rect 5629 11067 5687 11073
rect 5629 11033 5641 11067
rect 5675 11064 5687 11067
rect 5994 11064 6000 11076
rect 5675 11036 6000 11064
rect 5675 11033 5687 11036
rect 5629 11027 5687 11033
rect 5994 11024 6000 11036
rect 6052 11064 6058 11076
rect 6932 11064 6960 11095
rect 6052 11036 6960 11064
rect 6052 11024 6058 11036
rect 4154 10956 4160 11008
rect 4212 10996 4218 11008
rect 5261 10999 5319 11005
rect 5261 10996 5273 10999
rect 4212 10968 5273 10996
rect 4212 10956 4218 10968
rect 5261 10965 5273 10968
rect 5307 10965 5319 10999
rect 5261 10959 5319 10965
rect 5902 10956 5908 11008
rect 5960 10996 5966 11008
rect 6365 10999 6423 11005
rect 6365 10996 6377 10999
rect 5960 10968 6377 10996
rect 5960 10956 5966 10968
rect 6365 10965 6377 10968
rect 6411 10965 6423 10999
rect 6365 10959 6423 10965
rect 1104 10906 10488 10928
rect 1104 10854 4874 10906
rect 4926 10854 4938 10906
rect 4990 10854 5002 10906
rect 5054 10854 5066 10906
rect 5118 10854 5130 10906
rect 5182 10854 10488 10906
rect 1104 10832 10488 10854
rect 2774 10792 2780 10804
rect 2332 10764 2780 10792
rect 2332 10665 2360 10764
rect 2774 10752 2780 10764
rect 2832 10792 2838 10804
rect 2832 10764 3924 10792
rect 2832 10752 2838 10764
rect 2317 10659 2375 10665
rect 2317 10625 2329 10659
rect 2363 10625 2375 10659
rect 2317 10619 2375 10625
rect 3694 10616 3700 10668
rect 3752 10616 3758 10668
rect 3896 10656 3924 10764
rect 3970 10752 3976 10804
rect 4028 10792 4034 10804
rect 5905 10795 5963 10801
rect 4028 10764 5580 10792
rect 4028 10752 4034 10764
rect 4157 10659 4215 10665
rect 4157 10656 4169 10659
rect 3896 10628 4169 10656
rect 4157 10625 4169 10628
rect 4203 10625 4215 10659
rect 4157 10619 4215 10625
rect 2593 10591 2651 10597
rect 2593 10557 2605 10591
rect 2639 10588 2651 10591
rect 4433 10591 4491 10597
rect 2639 10560 4200 10588
rect 2639 10557 2651 10560
rect 2593 10551 2651 10557
rect 4172 10532 4200 10560
rect 4433 10557 4445 10591
rect 4479 10588 4491 10591
rect 4798 10588 4804 10600
rect 4479 10560 4804 10588
rect 4479 10557 4491 10560
rect 4433 10551 4491 10557
rect 4798 10548 4804 10560
rect 4856 10548 4862 10600
rect 5552 10588 5580 10764
rect 5905 10761 5917 10795
rect 5951 10792 5963 10795
rect 5994 10792 6000 10804
rect 5951 10764 6000 10792
rect 5951 10761 5963 10764
rect 5905 10755 5963 10761
rect 5994 10752 6000 10764
rect 6052 10752 6058 10804
rect 5810 10684 5816 10736
rect 5868 10684 5874 10736
rect 7190 10684 7196 10736
rect 7248 10684 7254 10736
rect 5828 10656 5856 10684
rect 6181 10659 6239 10665
rect 6181 10656 6193 10659
rect 5828 10628 6193 10656
rect 6181 10625 6193 10628
rect 6227 10625 6239 10659
rect 6181 10619 6239 10625
rect 5552 10560 6224 10588
rect 4154 10480 4160 10532
rect 4212 10480 4218 10532
rect 4062 10412 4068 10464
rect 4120 10452 4126 10464
rect 4246 10452 4252 10464
rect 4120 10424 4252 10452
rect 4120 10412 4126 10424
rect 4246 10412 4252 10424
rect 4304 10412 4310 10464
rect 6086 10412 6092 10464
rect 6144 10412 6150 10464
rect 6196 10452 6224 10560
rect 6270 10548 6276 10600
rect 6328 10588 6334 10600
rect 6365 10591 6423 10597
rect 6365 10588 6377 10591
rect 6328 10560 6377 10588
rect 6328 10548 6334 10560
rect 6365 10557 6377 10560
rect 6411 10557 6423 10591
rect 6365 10551 6423 10557
rect 6641 10591 6699 10597
rect 6641 10557 6653 10591
rect 6687 10588 6699 10591
rect 7374 10588 7380 10600
rect 6687 10560 7380 10588
rect 6687 10557 6699 10560
rect 6641 10551 6699 10557
rect 7374 10548 7380 10560
rect 7432 10548 7438 10600
rect 8757 10591 8815 10597
rect 8757 10588 8769 10591
rect 8128 10560 8769 10588
rect 8128 10464 8156 10560
rect 8757 10557 8769 10560
rect 8803 10557 8815 10591
rect 8757 10551 8815 10557
rect 6730 10452 6736 10464
rect 6196 10424 6736 10452
rect 6730 10412 6736 10424
rect 6788 10412 6794 10464
rect 8110 10412 8116 10464
rect 8168 10412 8174 10464
rect 8202 10412 8208 10464
rect 8260 10412 8266 10464
rect 1104 10362 10488 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 10488 10362
rect 1104 10288 10488 10310
rect 4798 10208 4804 10260
rect 4856 10208 4862 10260
rect 5353 10251 5411 10257
rect 5353 10217 5365 10251
rect 5399 10248 5411 10251
rect 6086 10248 6092 10260
rect 5399 10220 6092 10248
rect 5399 10217 5411 10220
rect 5353 10211 5411 10217
rect 6086 10208 6092 10220
rect 6144 10208 6150 10260
rect 6270 10208 6276 10260
rect 6328 10208 6334 10260
rect 1857 10115 1915 10121
rect 1857 10081 1869 10115
rect 1903 10112 1915 10115
rect 2774 10112 2780 10124
rect 1903 10084 2780 10112
rect 1903 10081 1915 10084
rect 1857 10075 1915 10081
rect 2774 10072 2780 10084
rect 2832 10072 2838 10124
rect 3605 10115 3663 10121
rect 3605 10081 3617 10115
rect 3651 10112 3663 10115
rect 5445 10115 5503 10121
rect 3651 10084 4476 10112
rect 3651 10081 3663 10084
rect 3605 10075 3663 10081
rect 4448 10056 4476 10084
rect 5445 10081 5457 10115
rect 5491 10112 5503 10115
rect 5902 10112 5908 10124
rect 5491 10084 5908 10112
rect 5491 10081 5503 10084
rect 5445 10075 5503 10081
rect 5902 10072 5908 10084
rect 5960 10072 5966 10124
rect 6181 10115 6239 10121
rect 6181 10081 6193 10115
rect 6227 10112 6239 10115
rect 6288 10112 6316 10208
rect 6227 10084 6316 10112
rect 6227 10081 6239 10084
rect 6181 10075 6239 10081
rect 7650 10072 7656 10124
rect 7708 10112 7714 10124
rect 8021 10115 8079 10121
rect 8021 10112 8033 10115
rect 7708 10084 8033 10112
rect 7708 10072 7714 10084
rect 8021 10081 8033 10084
rect 8067 10081 8079 10115
rect 8021 10075 8079 10081
rect 3234 10004 3240 10056
rect 3292 10044 3298 10056
rect 3694 10044 3700 10056
rect 3292 10016 3700 10044
rect 3292 10004 3298 10016
rect 3694 10004 3700 10016
rect 3752 10004 3758 10056
rect 4430 10004 4436 10056
rect 4488 10004 4494 10056
rect 4890 10004 4896 10056
rect 4948 10053 4954 10056
rect 4948 10047 4984 10053
rect 4972 10044 4984 10047
rect 4972 10016 5580 10044
rect 4972 10013 4984 10016
rect 4948 10007 4984 10013
rect 4948 10004 4954 10007
rect 1762 9936 1768 9988
rect 1820 9976 1826 9988
rect 2133 9979 2191 9985
rect 2133 9976 2145 9979
rect 1820 9948 2145 9976
rect 1820 9936 1826 9948
rect 2133 9945 2145 9948
rect 2179 9945 2191 9979
rect 5552 9976 5580 10016
rect 5626 10004 5632 10056
rect 5684 10044 5690 10056
rect 5721 10047 5779 10053
rect 5721 10044 5733 10047
rect 5684 10016 5733 10044
rect 5684 10004 5690 10016
rect 5721 10013 5733 10016
rect 5767 10013 5779 10047
rect 8481 10047 8539 10053
rect 8481 10044 8493 10047
rect 5721 10007 5779 10013
rect 8220 10016 8493 10044
rect 5552 9948 5764 9976
rect 2133 9939 2191 9945
rect 5736 9920 5764 9948
rect 5902 9936 5908 9988
rect 5960 9936 5966 9988
rect 6454 9936 6460 9988
rect 6512 9936 6518 9988
rect 6730 9936 6736 9988
rect 6788 9976 6794 9988
rect 6788 9948 6946 9976
rect 6788 9936 6794 9948
rect 8110 9936 8116 9988
rect 8168 9976 8174 9988
rect 8220 9985 8248 10016
rect 8481 10013 8493 10016
rect 8527 10013 8539 10047
rect 8481 10007 8539 10013
rect 8665 10047 8723 10053
rect 8665 10013 8677 10047
rect 8711 10044 8723 10047
rect 8711 10016 8745 10044
rect 8711 10013 8723 10016
rect 8665 10007 8723 10013
rect 8205 9979 8263 9985
rect 8205 9976 8217 9979
rect 8168 9948 8217 9976
rect 8168 9936 8174 9948
rect 8205 9945 8217 9948
rect 8251 9945 8263 9979
rect 8205 9939 8263 9945
rect 8389 9979 8447 9985
rect 8389 9945 8401 9979
rect 8435 9976 8447 9979
rect 8680 9976 8708 10007
rect 9030 9976 9036 9988
rect 8435 9948 9036 9976
rect 8435 9945 8447 9948
rect 8389 9939 8447 9945
rect 9030 9936 9036 9948
rect 9088 9936 9094 9988
rect 3786 9868 3792 9920
rect 3844 9868 3850 9920
rect 4985 9911 5043 9917
rect 4985 9877 4997 9911
rect 5031 9908 5043 9911
rect 5537 9911 5595 9917
rect 5537 9908 5549 9911
rect 5031 9880 5549 9908
rect 5031 9877 5043 9880
rect 4985 9871 5043 9877
rect 5537 9877 5549 9880
rect 5583 9877 5595 9911
rect 5537 9871 5595 9877
rect 5718 9868 5724 9920
rect 5776 9908 5782 9920
rect 6638 9908 6644 9920
rect 5776 9880 6644 9908
rect 5776 9868 5782 9880
rect 6638 9868 6644 9880
rect 6696 9868 6702 9920
rect 7466 9868 7472 9920
rect 7524 9908 7530 9920
rect 7929 9911 7987 9917
rect 7929 9908 7941 9911
rect 7524 9880 7941 9908
rect 7524 9868 7530 9880
rect 7929 9877 7941 9880
rect 7975 9908 7987 9911
rect 8018 9908 8024 9920
rect 7975 9880 8024 9908
rect 7975 9877 7987 9880
rect 7929 9871 7987 9877
rect 8018 9868 8024 9880
rect 8076 9868 8082 9920
rect 8294 9868 8300 9920
rect 8352 9908 8358 9920
rect 8481 9911 8539 9917
rect 8481 9908 8493 9911
rect 8352 9880 8493 9908
rect 8352 9868 8358 9880
rect 8481 9877 8493 9880
rect 8527 9877 8539 9911
rect 8481 9871 8539 9877
rect 1104 9818 10488 9840
rect 1104 9766 4874 9818
rect 4926 9766 4938 9818
rect 4990 9766 5002 9818
rect 5054 9766 5066 9818
rect 5118 9766 5130 9818
rect 5182 9766 10488 9818
rect 1104 9744 10488 9766
rect 3786 9704 3792 9716
rect 2746 9676 3792 9704
rect 2133 9571 2191 9577
rect 2133 9537 2145 9571
rect 2179 9568 2191 9571
rect 2746 9568 2774 9676
rect 3786 9664 3792 9676
rect 3844 9664 3850 9716
rect 4430 9664 4436 9716
rect 4488 9704 4494 9716
rect 5074 9704 5080 9716
rect 4488 9676 5080 9704
rect 4488 9664 4494 9676
rect 5074 9664 5080 9676
rect 5132 9664 5138 9716
rect 5258 9674 5264 9686
rect 5184 9646 5264 9674
rect 3237 9639 3295 9645
rect 3237 9605 3249 9639
rect 3283 9636 3295 9639
rect 5184 9636 5212 9646
rect 3283 9608 4016 9636
rect 3283 9605 3295 9608
rect 3237 9599 3295 9605
rect 2179 9540 2774 9568
rect 3329 9571 3387 9577
rect 2179 9537 2191 9540
rect 2133 9531 2191 9537
rect 3329 9537 3341 9571
rect 3375 9537 3387 9571
rect 3329 9531 3387 9537
rect 3421 9571 3479 9577
rect 3421 9537 3433 9571
rect 3467 9568 3479 9571
rect 3510 9568 3516 9580
rect 3467 9540 3516 9568
rect 3467 9537 3479 9540
rect 3421 9531 3479 9537
rect 1762 9460 1768 9512
rect 1820 9460 1826 9512
rect 2225 9503 2283 9509
rect 2225 9469 2237 9503
rect 2271 9500 2283 9503
rect 2314 9500 2320 9512
rect 2271 9472 2320 9500
rect 2271 9469 2283 9472
rect 2225 9463 2283 9469
rect 2314 9460 2320 9472
rect 2372 9500 2378 9512
rect 2409 9503 2467 9509
rect 2409 9500 2421 9503
rect 2372 9472 2421 9500
rect 2372 9460 2378 9472
rect 2409 9469 2421 9472
rect 2455 9469 2467 9503
rect 3344 9500 3372 9531
rect 3510 9528 3516 9540
rect 3568 9528 3574 9580
rect 3988 9509 4016 9608
rect 4816 9608 5212 9636
rect 5258 9634 5264 9646
rect 5316 9634 5322 9686
rect 5534 9664 5540 9716
rect 5592 9704 5598 9716
rect 5592 9676 5672 9704
rect 5592 9664 5598 9676
rect 5644 9674 5672 9676
rect 5644 9646 5764 9674
rect 5810 9664 5816 9716
rect 5868 9704 5874 9716
rect 5868 9676 6316 9704
rect 5868 9664 5874 9676
rect 5736 9636 5764 9646
rect 6288 9636 6316 9676
rect 6454 9664 6460 9716
rect 6512 9704 6518 9716
rect 6549 9707 6607 9713
rect 6549 9704 6561 9707
rect 6512 9676 6561 9704
rect 6512 9664 6518 9676
rect 6549 9673 6561 9676
rect 6595 9673 6607 9707
rect 6549 9667 6607 9673
rect 6638 9664 6644 9716
rect 6696 9704 6702 9716
rect 6917 9707 6975 9713
rect 6917 9704 6929 9707
rect 6696 9676 6929 9704
rect 6696 9664 6702 9676
rect 6917 9673 6929 9676
rect 6963 9673 6975 9707
rect 6917 9667 6975 9673
rect 7374 9664 7380 9716
rect 7432 9664 7438 9716
rect 7484 9676 7906 9704
rect 7009 9639 7067 9645
rect 7009 9636 7021 9639
rect 5736 9608 5948 9636
rect 6288 9608 7021 9636
rect 4062 9528 4068 9580
rect 4120 9528 4126 9580
rect 4816 9577 4844 9608
rect 4801 9571 4859 9577
rect 4801 9537 4813 9571
rect 4847 9537 4859 9571
rect 4801 9531 4859 9537
rect 4982 9528 4988 9580
rect 5040 9528 5046 9580
rect 5166 9528 5172 9580
rect 5224 9528 5230 9580
rect 5350 9528 5356 9580
rect 5408 9566 5414 9580
rect 5408 9538 5451 9566
rect 5408 9528 5414 9538
rect 5626 9528 5632 9580
rect 5684 9528 5690 9580
rect 5813 9571 5871 9577
rect 5813 9537 5825 9571
rect 5859 9566 5871 9571
rect 5920 9566 5948 9608
rect 7009 9605 7021 9608
rect 7055 9636 7067 9639
rect 7484 9636 7512 9676
rect 7055 9608 7512 9636
rect 7055 9605 7067 9608
rect 7009 9599 7067 9605
rect 5859 9538 5948 9566
rect 5859 9537 5871 9538
rect 5813 9531 5871 9537
rect 5994 9528 6000 9580
rect 6052 9528 6058 9580
rect 6638 9528 6644 9580
rect 6696 9528 6702 9580
rect 7558 9550 7564 9602
rect 7616 9550 7622 9602
rect 7650 9596 7656 9648
rect 7708 9596 7714 9648
rect 7878 9645 7906 9676
rect 8018 9664 8024 9716
rect 8076 9704 8082 9716
rect 8076 9676 8432 9704
rect 8076 9664 8082 9676
rect 7863 9639 7921 9645
rect 7863 9605 7875 9639
rect 7909 9605 7921 9639
rect 7863 9599 7921 9605
rect 8110 9596 8116 9648
rect 8168 9636 8174 9648
rect 8297 9639 8355 9645
rect 8297 9636 8309 9639
rect 8168 9608 8309 9636
rect 8168 9596 8174 9608
rect 8297 9605 8309 9608
rect 8343 9605 8355 9639
rect 8404 9636 8432 9676
rect 8404 9608 8524 9636
rect 8297 9599 8355 9605
rect 7746 9571 7804 9577
rect 7746 9568 7758 9571
rect 7561 9537 7573 9550
rect 7607 9537 7619 9550
rect 7561 9531 7619 9537
rect 7679 9540 7758 9568
rect 3973 9503 4031 9509
rect 3344 9472 3464 9500
rect 2409 9463 2467 9469
rect 2682 9392 2688 9444
rect 2740 9392 2746 9444
rect 3436 9376 3464 9472
rect 3973 9469 3985 9503
rect 4019 9469 4031 9503
rect 3973 9463 4031 9469
rect 4433 9503 4491 9509
rect 4433 9469 4445 9503
rect 4479 9500 4491 9503
rect 4706 9500 4712 9512
rect 4479 9472 4712 9500
rect 4479 9469 4491 9472
rect 4433 9463 4491 9469
rect 3605 9435 3663 9441
rect 3605 9401 3617 9435
rect 3651 9401 3663 9435
rect 3988 9432 4016 9463
rect 4706 9460 4712 9472
rect 4764 9460 4770 9512
rect 5537 9503 5595 9509
rect 5537 9469 5549 9503
rect 5583 9500 5595 9503
rect 6012 9500 6040 9528
rect 5583 9472 6040 9500
rect 5583 9469 5595 9472
rect 5537 9463 5595 9469
rect 5166 9432 5172 9444
rect 3988 9404 5172 9432
rect 3605 9395 3663 9401
rect 2866 9324 2872 9376
rect 2924 9324 2930 9376
rect 3053 9367 3111 9373
rect 3053 9333 3065 9367
rect 3099 9364 3111 9367
rect 3234 9364 3240 9376
rect 3099 9336 3240 9364
rect 3099 9333 3111 9336
rect 3053 9327 3111 9333
rect 3234 9324 3240 9336
rect 3292 9324 3298 9376
rect 3418 9324 3424 9376
rect 3476 9324 3482 9376
rect 3620 9364 3648 9395
rect 5166 9392 5172 9404
rect 5224 9392 5230 9444
rect 5994 9392 6000 9444
rect 6052 9392 6058 9444
rect 6656 9432 6684 9528
rect 7193 9503 7251 9509
rect 7193 9469 7205 9503
rect 7239 9500 7251 9503
rect 7466 9500 7472 9512
rect 7239 9472 7472 9500
rect 7239 9469 7251 9472
rect 7193 9463 7251 9469
rect 7466 9460 7472 9472
rect 7524 9460 7530 9512
rect 7679 9432 7707 9540
rect 7746 9537 7758 9540
rect 7792 9537 7804 9571
rect 8202 9568 8208 9580
rect 7746 9531 7804 9537
rect 8036 9540 8208 9568
rect 8036 9509 8064 9540
rect 8202 9528 8208 9540
rect 8260 9528 8266 9580
rect 8386 9528 8392 9580
rect 8444 9528 8450 9580
rect 8496 9577 8524 9608
rect 8481 9571 8539 9577
rect 8481 9537 8493 9571
rect 8527 9568 8539 9571
rect 9122 9568 9128 9580
rect 8527 9540 9128 9568
rect 8527 9537 8539 9540
rect 8481 9531 8539 9537
rect 9122 9528 9128 9540
rect 9180 9528 9186 9580
rect 8021 9503 8079 9509
rect 8021 9469 8033 9503
rect 8067 9469 8079 9503
rect 8021 9463 8079 9469
rect 8665 9435 8723 9441
rect 6656 9404 8294 9432
rect 4062 9364 4068 9376
rect 3620 9336 4068 9364
rect 4062 9324 4068 9336
rect 4120 9324 4126 9376
rect 4525 9367 4583 9373
rect 4525 9333 4537 9367
rect 4571 9364 4583 9367
rect 4614 9364 4620 9376
rect 4571 9336 4620 9364
rect 4571 9333 4583 9336
rect 4525 9327 4583 9333
rect 4614 9324 4620 9336
rect 4672 9324 4678 9376
rect 4801 9367 4859 9373
rect 4801 9333 4813 9367
rect 4847 9364 4859 9367
rect 5258 9364 5264 9376
rect 4847 9336 5264 9364
rect 4847 9333 4859 9336
rect 4801 9327 4859 9333
rect 5258 9324 5264 9336
rect 5316 9324 5322 9376
rect 6638 9324 6644 9376
rect 6696 9364 6702 9376
rect 8113 9367 8171 9373
rect 8113 9364 8125 9367
rect 6696 9336 8125 9364
rect 6696 9324 6702 9336
rect 8113 9333 8125 9336
rect 8159 9333 8171 9367
rect 8266 9364 8294 9404
rect 8665 9401 8677 9435
rect 8711 9432 8723 9435
rect 8754 9432 8760 9444
rect 8711 9404 8760 9432
rect 8711 9401 8723 9404
rect 8665 9395 8723 9401
rect 8754 9392 8760 9404
rect 8812 9392 8818 9444
rect 8846 9364 8852 9376
rect 8266 9336 8852 9364
rect 8113 9327 8171 9333
rect 8846 9324 8852 9336
rect 8904 9324 8910 9376
rect 1104 9274 10488 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 10488 9274
rect 1104 9200 10488 9222
rect 2866 9120 2872 9172
rect 2924 9169 2930 9172
rect 2924 9163 2939 9169
rect 2927 9129 2939 9163
rect 2924 9123 2939 9129
rect 2924 9120 2930 9123
rect 4246 9120 4252 9172
rect 4304 9160 4310 9172
rect 4709 9163 4767 9169
rect 4709 9160 4721 9163
rect 4304 9132 4721 9160
rect 4304 9120 4310 9132
rect 4709 9129 4721 9132
rect 4755 9129 4767 9163
rect 4709 9123 4767 9129
rect 4982 9120 4988 9172
rect 5040 9160 5046 9172
rect 5442 9160 5448 9172
rect 5040 9132 5448 9160
rect 5040 9120 5046 9132
rect 5442 9120 5448 9132
rect 5500 9120 5506 9172
rect 5537 9163 5595 9169
rect 5537 9129 5549 9163
rect 5583 9160 5595 9163
rect 6086 9160 6092 9172
rect 5583 9132 6092 9160
rect 5583 9129 5595 9132
rect 5537 9123 5595 9129
rect 6086 9120 6092 9132
rect 6144 9160 6150 9172
rect 7006 9160 7012 9172
rect 6144 9132 7012 9160
rect 6144 9120 6150 9132
rect 7006 9120 7012 9132
rect 7064 9120 7070 9172
rect 7653 9163 7711 9169
rect 7653 9129 7665 9163
rect 7699 9160 7711 9163
rect 8386 9160 8392 9172
rect 7699 9132 8392 9160
rect 7699 9129 7711 9132
rect 7653 9123 7711 9129
rect 8386 9120 8392 9132
rect 8444 9120 8450 9172
rect 4338 9052 4344 9104
rect 4396 9092 4402 9104
rect 5626 9092 5632 9104
rect 4396 9064 5632 9092
rect 4396 9052 4402 9064
rect 5626 9052 5632 9064
rect 5684 9052 5690 9104
rect 5718 9052 5724 9104
rect 5776 9052 5782 9104
rect 5810 9052 5816 9104
rect 5868 9092 5874 9104
rect 5905 9095 5963 9101
rect 5905 9092 5917 9095
rect 5868 9064 5917 9092
rect 5868 9052 5874 9064
rect 5905 9061 5917 9064
rect 5951 9061 5963 9095
rect 5905 9055 5963 9061
rect 6362 9052 6368 9104
rect 6420 9052 6426 9104
rect 7558 9052 7564 9104
rect 7616 9092 7622 9104
rect 8478 9092 8484 9104
rect 7616 9064 8484 9092
rect 7616 9052 7622 9064
rect 8478 9052 8484 9064
rect 8536 9052 8542 9104
rect 2774 8984 2780 9036
rect 2832 9024 2838 9036
rect 3145 9027 3203 9033
rect 3145 9024 3157 9027
rect 2832 8996 3157 9024
rect 2832 8984 2838 8996
rect 3145 8993 3157 8996
rect 3191 8993 3203 9027
rect 3145 8987 3203 8993
rect 3973 9027 4031 9033
rect 3973 8993 3985 9027
rect 4019 9024 4031 9027
rect 4522 9024 4528 9036
rect 4019 8996 4528 9024
rect 4019 8993 4031 8996
rect 3973 8987 4031 8993
rect 4522 8984 4528 8996
rect 4580 9024 4586 9036
rect 5169 9027 5227 9033
rect 5169 9024 5181 9027
rect 4580 8996 5181 9024
rect 4580 8984 4586 8996
rect 5169 8993 5181 8996
rect 5215 9024 5227 9027
rect 6380 9024 6408 9052
rect 7009 9027 7067 9033
rect 5215 8996 6684 9024
rect 5215 8993 5227 8996
rect 5169 8987 5227 8993
rect 3605 8959 3663 8965
rect 3605 8925 3617 8959
rect 3651 8956 3663 8959
rect 4065 8959 4123 8965
rect 3651 8928 4016 8956
rect 3651 8925 3663 8928
rect 3605 8919 3663 8925
rect 3142 8888 3148 8900
rect 2438 8860 3148 8888
rect 3142 8848 3148 8860
rect 3200 8848 3206 8900
rect 1394 8780 1400 8832
rect 1452 8780 1458 8832
rect 3418 8780 3424 8832
rect 3476 8780 3482 8832
rect 3786 8780 3792 8832
rect 3844 8780 3850 8832
rect 3988 8820 4016 8928
rect 4065 8925 4077 8959
rect 4111 8925 4123 8959
rect 4065 8919 4123 8925
rect 4080 8888 4108 8919
rect 4430 8916 4436 8968
rect 4488 8916 4494 8968
rect 4709 8959 4767 8965
rect 4709 8958 4721 8959
rect 4632 8930 4721 8958
rect 4632 8888 4660 8930
rect 4709 8925 4721 8930
rect 4755 8925 4767 8959
rect 4709 8919 4767 8925
rect 5074 8916 5080 8968
rect 5132 8916 5138 8968
rect 5813 8959 5871 8965
rect 5813 8956 5825 8959
rect 5736 8928 5825 8956
rect 4080 8860 4660 8888
rect 4632 8832 4660 8860
rect 4154 8820 4160 8832
rect 3988 8792 4160 8820
rect 4154 8780 4160 8792
rect 4212 8780 4218 8832
rect 4246 8780 4252 8832
rect 4304 8780 4310 8832
rect 4338 8780 4344 8832
rect 4396 8780 4402 8832
rect 4430 8780 4436 8832
rect 4488 8820 4494 8832
rect 4525 8823 4583 8829
rect 4525 8820 4537 8823
rect 4488 8792 4537 8820
rect 4488 8780 4494 8792
rect 4525 8789 4537 8792
rect 4571 8789 4583 8823
rect 4525 8783 4583 8789
rect 4614 8780 4620 8832
rect 4672 8780 4678 8832
rect 5537 8823 5595 8829
rect 5537 8789 5549 8823
rect 5583 8820 5595 8823
rect 5736 8820 5764 8928
rect 5813 8925 5825 8928
rect 5859 8925 5871 8959
rect 5813 8919 5871 8925
rect 6086 8916 6092 8968
rect 6144 8916 6150 8968
rect 6656 8965 6684 8996
rect 7009 8993 7021 9027
rect 7055 9024 7067 9027
rect 8662 9024 8668 9036
rect 7055 8996 8668 9024
rect 7055 8993 7067 8996
rect 7009 8987 7067 8993
rect 8662 8984 8668 8996
rect 8720 8984 8726 9036
rect 6365 8959 6423 8965
rect 6365 8925 6377 8959
rect 6411 8925 6423 8959
rect 6549 8959 6607 8965
rect 6549 8956 6561 8959
rect 6365 8919 6423 8925
rect 6472 8928 6561 8956
rect 5810 8820 5816 8832
rect 5583 8792 5816 8820
rect 5583 8789 5595 8792
rect 5537 8783 5595 8789
rect 5810 8780 5816 8792
rect 5868 8820 5874 8832
rect 6380 8820 6408 8919
rect 6472 8832 6500 8928
rect 6549 8925 6561 8928
rect 6595 8925 6607 8959
rect 6549 8919 6607 8925
rect 6641 8959 6699 8965
rect 6641 8925 6653 8959
rect 6687 8925 6699 8959
rect 6641 8919 6699 8925
rect 6733 8959 6791 8965
rect 6733 8925 6745 8959
rect 6779 8956 6791 8959
rect 7285 8959 7343 8965
rect 7285 8956 7297 8959
rect 6779 8928 7297 8956
rect 6779 8925 6791 8928
rect 6733 8919 6791 8925
rect 7285 8925 7297 8928
rect 7331 8956 7343 8959
rect 7374 8956 7380 8968
rect 7331 8928 7380 8956
rect 7331 8925 7343 8928
rect 7285 8919 7343 8925
rect 7374 8916 7380 8928
rect 7432 8916 7438 8968
rect 7469 8959 7527 8965
rect 7469 8925 7481 8959
rect 7515 8925 7527 8959
rect 7469 8919 7527 8925
rect 7745 8959 7803 8965
rect 7745 8925 7757 8959
rect 7791 8956 7803 8959
rect 8021 8959 8079 8965
rect 8021 8956 8033 8959
rect 7791 8928 8033 8956
rect 7791 8925 7803 8928
rect 7745 8919 7803 8925
rect 8021 8925 8033 8928
rect 8067 8956 8079 8959
rect 8294 8956 8300 8968
rect 8067 8928 8300 8956
rect 8067 8925 8079 8928
rect 8021 8919 8079 8925
rect 7484 8888 7512 8919
rect 8294 8916 8300 8928
rect 8352 8956 8358 8968
rect 8754 8956 8760 8968
rect 8352 8928 8760 8956
rect 8352 8916 8358 8928
rect 8754 8916 8760 8928
rect 8812 8916 8818 8968
rect 7484 8860 8064 8888
rect 8036 8832 8064 8860
rect 5868 8792 6408 8820
rect 5868 8780 5874 8792
rect 6454 8780 6460 8832
rect 6512 8780 6518 8832
rect 6914 8780 6920 8832
rect 6972 8820 6978 8832
rect 7101 8823 7159 8829
rect 7101 8820 7113 8823
rect 6972 8792 7113 8820
rect 6972 8780 6978 8792
rect 7101 8789 7113 8792
rect 7147 8789 7159 8823
rect 7101 8783 7159 8789
rect 8018 8780 8024 8832
rect 8076 8780 8082 8832
rect 8570 8780 8576 8832
rect 8628 8780 8634 8832
rect 1104 8730 10488 8752
rect 1104 8678 4874 8730
rect 4926 8678 4938 8730
rect 4990 8678 5002 8730
rect 5054 8678 5066 8730
rect 5118 8678 5130 8730
rect 5182 8678 10488 8730
rect 1104 8656 10488 8678
rect 1394 8576 1400 8628
rect 1452 8576 1458 8628
rect 2682 8576 2688 8628
rect 2740 8576 2746 8628
rect 3053 8619 3111 8625
rect 3053 8585 3065 8619
rect 3099 8585 3111 8619
rect 3053 8579 3111 8585
rect 3237 8619 3295 8625
rect 3237 8585 3249 8619
rect 3283 8616 3295 8619
rect 3418 8616 3424 8628
rect 3283 8588 3424 8616
rect 3283 8585 3295 8588
rect 3237 8579 3295 8585
rect 1412 8480 1440 8576
rect 2866 8508 2872 8560
rect 2924 8548 2930 8560
rect 3068 8548 3096 8579
rect 3418 8576 3424 8588
rect 3476 8616 3482 8628
rect 3878 8616 3884 8628
rect 3476 8588 3884 8616
rect 3476 8576 3482 8588
rect 3878 8576 3884 8588
rect 3936 8576 3942 8628
rect 4338 8576 4344 8628
rect 4396 8576 4402 8628
rect 4433 8619 4491 8625
rect 4433 8585 4445 8619
rect 4479 8616 4491 8619
rect 4479 8588 4660 8616
rect 4479 8585 4491 8588
rect 4433 8579 4491 8585
rect 3510 8548 3516 8560
rect 2924 8520 3516 8548
rect 2924 8508 2930 8520
rect 3510 8508 3516 8520
rect 3568 8508 3574 8560
rect 3786 8508 3792 8560
rect 3844 8508 3850 8560
rect 4356 8548 4384 8576
rect 3896 8520 4384 8548
rect 1489 8483 1547 8489
rect 1489 8480 1501 8483
rect 1412 8452 1501 8480
rect 1489 8449 1501 8452
rect 1535 8449 1547 8483
rect 1489 8443 1547 8449
rect 1673 8483 1731 8489
rect 1673 8449 1685 8483
rect 1719 8480 1731 8483
rect 2406 8480 2412 8492
rect 1719 8452 2412 8480
rect 1719 8449 1731 8452
rect 1673 8443 1731 8449
rect 1504 8412 1532 8443
rect 2406 8440 2412 8452
rect 2464 8480 2470 8492
rect 2961 8483 3019 8489
rect 2961 8480 2973 8483
rect 2464 8452 2973 8480
rect 2464 8440 2470 8452
rect 2961 8449 2973 8452
rect 3007 8449 3019 8483
rect 2961 8443 3019 8449
rect 3329 8483 3387 8489
rect 3329 8449 3341 8483
rect 3375 8480 3387 8483
rect 3804 8480 3832 8508
rect 3896 8489 3924 8520
rect 3375 8452 3832 8480
rect 3881 8483 3939 8489
rect 3375 8449 3387 8452
rect 3329 8443 3387 8449
rect 3881 8449 3893 8483
rect 3927 8449 3939 8483
rect 3881 8443 3939 8449
rect 4249 8483 4307 8489
rect 4249 8449 4261 8483
rect 4295 8480 4307 8483
rect 4430 8480 4436 8492
rect 4295 8452 4436 8480
rect 4295 8449 4307 8452
rect 4249 8443 4307 8449
rect 4430 8440 4436 8452
rect 4488 8440 4494 8492
rect 4632 8480 4660 8588
rect 4706 8576 4712 8628
rect 4764 8576 4770 8628
rect 5534 8576 5540 8628
rect 5592 8616 5598 8628
rect 5592 8588 6132 8616
rect 5592 8576 5598 8588
rect 4724 8548 4752 8576
rect 4724 8520 5028 8548
rect 5000 8489 5028 8520
rect 5092 8520 5764 8548
rect 5092 8489 5120 8520
rect 5736 8492 5764 8520
rect 4985 8483 5043 8489
rect 4632 8452 4752 8480
rect 1949 8415 2007 8421
rect 1949 8412 1961 8415
rect 1504 8384 1961 8412
rect 1949 8381 1961 8384
rect 1995 8381 2007 8415
rect 1949 8375 2007 8381
rect 2593 8415 2651 8421
rect 2593 8381 2605 8415
rect 2639 8412 2651 8415
rect 2869 8415 2927 8421
rect 2869 8412 2881 8415
rect 2639 8384 2881 8412
rect 2639 8381 2651 8384
rect 2593 8375 2651 8381
rect 2869 8381 2881 8384
rect 2915 8381 2927 8415
rect 2869 8375 2927 8381
rect 3789 8415 3847 8421
rect 3789 8381 3801 8415
rect 3835 8381 3847 8415
rect 3789 8375 3847 8381
rect 1857 8347 1915 8353
rect 1857 8313 1869 8347
rect 1903 8344 1915 8347
rect 2682 8344 2688 8356
rect 1903 8316 2688 8344
rect 1903 8313 1915 8316
rect 1857 8307 1915 8313
rect 2682 8304 2688 8316
rect 2740 8344 2746 8356
rect 3804 8344 3832 8375
rect 4154 8372 4160 8424
rect 4212 8412 4218 8424
rect 4724 8412 4752 8452
rect 4985 8449 4997 8483
rect 5031 8449 5043 8483
rect 4985 8443 5043 8449
rect 5077 8483 5135 8489
rect 5077 8449 5089 8483
rect 5123 8449 5135 8483
rect 5077 8443 5135 8449
rect 5445 8483 5503 8489
rect 5445 8449 5457 8483
rect 5491 8480 5503 8483
rect 5626 8480 5632 8492
rect 5491 8452 5632 8480
rect 5491 8449 5503 8452
rect 5445 8443 5503 8449
rect 5626 8440 5632 8452
rect 5684 8440 5690 8492
rect 5718 8440 5724 8492
rect 5776 8440 5782 8492
rect 6104 8489 6132 8588
rect 6638 8576 6644 8628
rect 6696 8576 6702 8628
rect 6733 8619 6791 8625
rect 6733 8585 6745 8619
rect 6779 8616 6791 8619
rect 8294 8616 8300 8628
rect 6779 8588 8300 8616
rect 6779 8585 6791 8588
rect 6733 8579 6791 8585
rect 8294 8576 8300 8588
rect 8352 8576 8358 8628
rect 8570 8576 8576 8628
rect 8628 8576 8634 8628
rect 8662 8576 8668 8628
rect 8720 8576 8726 8628
rect 9030 8576 9036 8628
rect 9088 8576 9094 8628
rect 6089 8483 6147 8489
rect 6089 8449 6101 8483
rect 6135 8480 6147 8483
rect 6178 8480 6184 8492
rect 6135 8452 6184 8480
rect 6135 8449 6147 8452
rect 6089 8443 6147 8449
rect 6178 8440 6184 8452
rect 6236 8480 6242 8492
rect 6365 8483 6423 8489
rect 6365 8480 6377 8483
rect 6236 8452 6377 8480
rect 6236 8440 6242 8452
rect 6365 8449 6377 8452
rect 6411 8449 6423 8483
rect 6365 8443 6423 8449
rect 6549 8483 6607 8489
rect 6549 8449 6561 8483
rect 6595 8480 6607 8483
rect 6656 8480 6684 8576
rect 7190 8508 7196 8560
rect 7248 8508 7254 8560
rect 6595 8452 6684 8480
rect 6595 8449 6607 8452
rect 6549 8443 6607 8449
rect 5169 8415 5227 8421
rect 4212 8384 5120 8412
rect 4212 8372 4218 8384
rect 5092 8356 5120 8384
rect 5169 8381 5181 8415
rect 5215 8381 5227 8415
rect 5169 8375 5227 8381
rect 5261 8415 5319 8421
rect 5261 8381 5273 8415
rect 5307 8412 5319 8415
rect 5537 8415 5595 8421
rect 5537 8412 5549 8415
rect 5307 8384 5549 8412
rect 5307 8381 5319 8384
rect 5261 8375 5319 8381
rect 5537 8381 5549 8384
rect 5583 8381 5595 8415
rect 5537 8375 5595 8381
rect 2740 8316 3832 8344
rect 4356 8316 4936 8344
rect 2740 8304 2746 8316
rect 4249 8279 4307 8285
rect 4249 8245 4261 8279
rect 4295 8276 4307 8279
rect 4356 8276 4384 8316
rect 4295 8248 4384 8276
rect 4295 8245 4307 8248
rect 4249 8239 4307 8245
rect 4706 8236 4712 8288
rect 4764 8276 4770 8288
rect 4801 8279 4859 8285
rect 4801 8276 4813 8279
rect 4764 8248 4813 8276
rect 4764 8236 4770 8248
rect 4801 8245 4813 8248
rect 4847 8245 4859 8279
rect 4908 8276 4936 8316
rect 5074 8304 5080 8356
rect 5132 8304 5138 8356
rect 5184 8344 5212 8375
rect 5994 8372 6000 8424
rect 6052 8412 6058 8424
rect 6564 8412 6592 8443
rect 8478 8440 8484 8492
rect 8536 8440 8542 8492
rect 8588 8480 8616 8576
rect 8680 8548 8708 8576
rect 8680 8520 8800 8548
rect 8665 8483 8723 8489
rect 8665 8480 8677 8483
rect 8588 8452 8677 8480
rect 8665 8449 8677 8452
rect 8711 8449 8723 8483
rect 8665 8443 8723 8449
rect 6052 8384 6592 8412
rect 8205 8415 8263 8421
rect 6052 8372 6058 8384
rect 8205 8381 8217 8415
rect 8251 8412 8263 8415
rect 8573 8415 8631 8421
rect 8251 8384 8524 8412
rect 8251 8381 8263 8384
rect 8205 8375 8263 8381
rect 6457 8347 6515 8353
rect 6457 8344 6469 8347
rect 5184 8316 6469 8344
rect 6457 8313 6469 8316
rect 6503 8313 6515 8347
rect 8496 8344 8524 8384
rect 8573 8381 8585 8415
rect 8619 8412 8631 8415
rect 8772 8412 8800 8520
rect 8846 8440 8852 8492
rect 8904 8480 8910 8492
rect 9036 8483 9094 8489
rect 9036 8480 9048 8483
rect 8904 8452 9048 8480
rect 8904 8440 8910 8452
rect 9036 8449 9048 8452
rect 9082 8449 9094 8483
rect 9036 8443 9094 8449
rect 8619 8384 8800 8412
rect 8619 8381 8631 8384
rect 8573 8375 8631 8381
rect 9217 8347 9275 8353
rect 9217 8344 9229 8347
rect 6457 8307 6515 8313
rect 6656 8316 6960 8344
rect 8496 8316 9229 8344
rect 6656 8276 6684 8316
rect 6932 8288 6960 8316
rect 9217 8313 9229 8316
rect 9263 8313 9275 8347
rect 9217 8307 9275 8313
rect 4908 8248 6684 8276
rect 4801 8239 4859 8245
rect 6914 8236 6920 8288
rect 6972 8236 6978 8288
rect 1104 8186 10488 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 10488 8186
rect 1104 8112 10488 8134
rect 2314 8032 2320 8084
rect 2372 8032 2378 8084
rect 6270 8032 6276 8084
rect 6328 8032 6334 8084
rect 2958 7964 2964 8016
rect 3016 7964 3022 8016
rect 5074 7964 5080 8016
rect 5132 8004 5138 8016
rect 5534 8004 5540 8016
rect 5132 7976 5540 8004
rect 5132 7964 5138 7976
rect 5534 7964 5540 7976
rect 5592 7964 5598 8016
rect 1670 7896 1676 7948
rect 1728 7896 1734 7948
rect 2133 7939 2191 7945
rect 2133 7905 2145 7939
rect 2179 7936 2191 7939
rect 6288 7936 6316 8032
rect 8386 7964 8392 8016
rect 8444 8004 8450 8016
rect 8444 7976 9536 8004
rect 8444 7964 8450 7976
rect 6641 7939 6699 7945
rect 6641 7936 6653 7939
rect 2179 7908 4476 7936
rect 6288 7908 6653 7936
rect 2179 7905 2191 7908
rect 2133 7899 2191 7905
rect 1394 7828 1400 7880
rect 1452 7828 1458 7880
rect 2038 7828 2044 7880
rect 2096 7828 2102 7880
rect 2682 7828 2688 7880
rect 2740 7828 2746 7880
rect 3160 7877 3188 7908
rect 3145 7871 3203 7877
rect 2792 7840 3004 7868
rect 2501 7803 2559 7809
rect 2501 7769 2513 7803
rect 2547 7800 2559 7803
rect 2792 7800 2820 7840
rect 2547 7772 2820 7800
rect 2547 7769 2559 7772
rect 2501 7763 2559 7769
rect 2866 7760 2872 7812
rect 2924 7760 2930 7812
rect 2976 7800 3004 7840
rect 3145 7837 3157 7871
rect 3191 7837 3203 7871
rect 3145 7831 3203 7837
rect 3234 7828 3240 7880
rect 3292 7868 3298 7880
rect 3421 7871 3479 7877
rect 3421 7868 3433 7871
rect 3292 7840 3433 7868
rect 3292 7828 3298 7840
rect 3421 7837 3433 7840
rect 3467 7837 3479 7871
rect 3421 7831 3479 7837
rect 3605 7871 3663 7877
rect 3605 7837 3617 7871
rect 3651 7837 3663 7871
rect 3605 7831 3663 7837
rect 3620 7800 3648 7831
rect 3878 7828 3884 7880
rect 3936 7868 3942 7880
rect 3973 7871 4031 7877
rect 3973 7868 3985 7871
rect 3936 7840 3985 7868
rect 3936 7828 3942 7840
rect 3973 7837 3985 7840
rect 4019 7837 4031 7871
rect 3973 7831 4031 7837
rect 4448 7812 4476 7908
rect 6641 7905 6653 7908
rect 6687 7936 6699 7939
rect 8478 7936 8484 7948
rect 6687 7908 8484 7936
rect 6687 7905 6699 7908
rect 6641 7899 6699 7905
rect 8478 7896 8484 7908
rect 8536 7896 8542 7948
rect 9508 7945 9536 7976
rect 9493 7939 9551 7945
rect 9493 7905 9505 7939
rect 9539 7905 9551 7939
rect 9493 7899 9551 7905
rect 4614 7828 4620 7880
rect 4672 7828 4678 7880
rect 4798 7828 4804 7880
rect 4856 7828 4862 7880
rect 4065 7803 4123 7809
rect 4065 7800 4077 7803
rect 2976 7772 3556 7800
rect 3620 7772 4077 7800
rect 1578 7692 1584 7744
rect 1636 7692 1642 7744
rect 2593 7735 2651 7741
rect 2593 7701 2605 7735
rect 2639 7732 2651 7735
rect 3418 7732 3424 7744
rect 2639 7704 3424 7732
rect 2639 7701 2651 7704
rect 2593 7695 2651 7701
rect 3418 7692 3424 7704
rect 3476 7692 3482 7744
rect 3528 7732 3556 7772
rect 4065 7769 4077 7772
rect 4111 7769 4123 7803
rect 4065 7763 4123 7769
rect 4430 7760 4436 7812
rect 4488 7760 4494 7812
rect 6914 7760 6920 7812
rect 6972 7760 6978 7812
rect 7190 7760 7196 7812
rect 7248 7800 7254 7812
rect 7248 7772 7406 7800
rect 7248 7760 7254 7772
rect 3602 7732 3608 7744
rect 3528 7704 3608 7732
rect 3602 7692 3608 7704
rect 3660 7692 3666 7744
rect 3694 7692 3700 7744
rect 3752 7732 3758 7744
rect 3881 7735 3939 7741
rect 3881 7732 3893 7735
rect 3752 7704 3893 7732
rect 3752 7692 3758 7704
rect 3881 7701 3893 7704
rect 3927 7701 3939 7735
rect 3881 7695 3939 7701
rect 4338 7692 4344 7744
rect 4396 7732 4402 7744
rect 6086 7732 6092 7744
rect 4396 7704 6092 7732
rect 4396 7692 4402 7704
rect 6086 7692 6092 7704
rect 6144 7692 6150 7744
rect 6270 7692 6276 7744
rect 6328 7732 6334 7744
rect 6730 7732 6736 7744
rect 6328 7704 6736 7732
rect 6328 7692 6334 7704
rect 6730 7692 6736 7704
rect 6788 7692 6794 7744
rect 7300 7732 7328 7772
rect 7742 7732 7748 7744
rect 7300 7704 7748 7732
rect 7742 7692 7748 7704
rect 7800 7692 7806 7744
rect 8938 7692 8944 7744
rect 8996 7692 9002 7744
rect 1104 7642 10488 7664
rect 1104 7590 4874 7642
rect 4926 7590 4938 7642
rect 4990 7590 5002 7642
rect 5054 7590 5066 7642
rect 5118 7590 5130 7642
rect 5182 7590 10488 7642
rect 1104 7568 10488 7590
rect 1118 7488 1124 7540
rect 1176 7528 1182 7540
rect 1489 7531 1547 7537
rect 1489 7528 1501 7531
rect 1176 7500 1501 7528
rect 1176 7488 1182 7500
rect 1489 7497 1501 7500
rect 1535 7497 1547 7531
rect 1489 7491 1547 7497
rect 1857 7531 1915 7537
rect 1857 7497 1869 7531
rect 1903 7528 1915 7531
rect 2038 7528 2044 7540
rect 1903 7500 2044 7528
rect 1903 7497 1915 7500
rect 1857 7491 1915 7497
rect 2038 7488 2044 7500
rect 2096 7488 2102 7540
rect 2774 7488 2780 7540
rect 2832 7528 2838 7540
rect 2869 7531 2927 7537
rect 2869 7528 2881 7531
rect 2832 7500 2881 7528
rect 2832 7488 2838 7500
rect 2869 7497 2881 7500
rect 2915 7497 2927 7531
rect 2869 7491 2927 7497
rect 1673 7395 1731 7401
rect 1673 7361 1685 7395
rect 1719 7392 1731 7395
rect 2884 7392 2912 7491
rect 6086 7488 6092 7540
rect 6144 7488 6150 7540
rect 6178 7488 6184 7540
rect 6236 7488 6242 7540
rect 6733 7531 6791 7537
rect 6733 7497 6745 7531
rect 6779 7528 6791 7531
rect 6914 7528 6920 7540
rect 6779 7500 6920 7528
rect 6779 7497 6791 7500
rect 6733 7491 6791 7497
rect 6914 7488 6920 7500
rect 6972 7488 6978 7540
rect 8478 7488 8484 7540
rect 8536 7528 8542 7540
rect 9033 7531 9091 7537
rect 9033 7528 9045 7531
rect 8536 7500 9045 7528
rect 8536 7488 8542 7500
rect 9033 7497 9045 7500
rect 9079 7497 9091 7531
rect 9033 7491 9091 7497
rect 4338 7420 4344 7472
rect 4396 7420 4402 7472
rect 4706 7420 4712 7472
rect 4764 7420 4770 7472
rect 6104 7460 6132 7488
rect 7745 7463 7803 7469
rect 7745 7460 7757 7463
rect 6104 7432 7757 7460
rect 7745 7429 7757 7432
rect 7791 7429 7803 7463
rect 7745 7423 7803 7429
rect 8938 7420 8944 7472
rect 8996 7420 9002 7472
rect 4433 7395 4491 7401
rect 4433 7392 4445 7395
rect 1719 7364 2774 7392
rect 2884 7364 4445 7392
rect 1719 7361 1731 7364
rect 1673 7355 1731 7361
rect 2406 7284 2412 7336
rect 2464 7284 2470 7336
rect 2746 7324 2774 7364
rect 4433 7361 4445 7364
rect 4479 7361 4491 7395
rect 4433 7355 4491 7361
rect 5718 7352 5724 7404
rect 5776 7352 5782 7404
rect 6270 7392 6276 7404
rect 5842 7364 6276 7392
rect 6270 7352 6276 7364
rect 6328 7352 6334 7404
rect 6549 7395 6607 7401
rect 6549 7361 6561 7395
rect 6595 7392 6607 7395
rect 6822 7392 6828 7404
rect 6595 7364 6828 7392
rect 6595 7361 6607 7364
rect 6549 7355 6607 7361
rect 6822 7352 6828 7364
rect 6880 7352 6886 7404
rect 6917 7395 6975 7401
rect 6917 7361 6929 7395
rect 6963 7361 6975 7395
rect 6917 7355 6975 7361
rect 7193 7395 7251 7401
rect 7193 7361 7205 7395
rect 7239 7392 7251 7395
rect 7282 7392 7288 7404
rect 7239 7364 7288 7392
rect 7239 7361 7251 7364
rect 7193 7355 7251 7361
rect 2866 7324 2872 7336
rect 2746 7296 2872 7324
rect 2866 7284 2872 7296
rect 2924 7324 2930 7336
rect 3602 7324 3608 7336
rect 2924 7296 3608 7324
rect 2924 7284 2930 7296
rect 3602 7284 3608 7296
rect 3660 7284 3666 7336
rect 5736 7324 5764 7352
rect 6932 7324 6960 7355
rect 7282 7352 7288 7364
rect 7340 7352 7346 7404
rect 7377 7395 7435 7401
rect 7377 7361 7389 7395
rect 7423 7361 7435 7395
rect 7377 7355 7435 7361
rect 7653 7395 7711 7401
rect 7653 7361 7665 7395
rect 7699 7392 7711 7395
rect 7926 7392 7932 7404
rect 7699 7364 7932 7392
rect 7699 7361 7711 7364
rect 7653 7355 7711 7361
rect 5736 7296 6960 7324
rect 7392 7324 7420 7355
rect 7926 7352 7932 7364
rect 7984 7352 7990 7404
rect 8956 7324 8984 7420
rect 7392 7296 8984 7324
rect 6270 7216 6276 7268
rect 6328 7256 6334 7268
rect 7006 7256 7012 7268
rect 6328 7228 7012 7256
rect 6328 7216 6334 7228
rect 7006 7216 7012 7228
rect 7064 7256 7070 7268
rect 7064 7228 7972 7256
rect 7064 7216 7070 7228
rect 7944 7200 7972 7228
rect 4430 7148 4436 7200
rect 4488 7188 4494 7200
rect 4798 7188 4804 7200
rect 4488 7160 4804 7188
rect 4488 7148 4494 7160
rect 4798 7148 4804 7160
rect 4856 7148 4862 7200
rect 6362 7148 6368 7200
rect 6420 7188 6426 7200
rect 6457 7191 6515 7197
rect 6457 7188 6469 7191
rect 6420 7160 6469 7188
rect 6420 7148 6426 7160
rect 6457 7157 6469 7160
rect 6503 7157 6515 7191
rect 6457 7151 6515 7157
rect 6822 7148 6828 7200
rect 6880 7188 6886 7200
rect 7466 7188 7472 7200
rect 6880 7160 7472 7188
rect 6880 7148 6886 7160
rect 7466 7148 7472 7160
rect 7524 7148 7530 7200
rect 7558 7148 7564 7200
rect 7616 7148 7622 7200
rect 7926 7148 7932 7200
rect 7984 7148 7990 7200
rect 1104 7098 10488 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 10488 7098
rect 1104 7024 10488 7046
rect 1670 6993 1676 6996
rect 1660 6987 1676 6993
rect 1660 6953 1672 6987
rect 1660 6947 1676 6953
rect 1670 6944 1676 6947
rect 1728 6944 1734 6996
rect 2774 6984 2780 6996
rect 2746 6944 2780 6984
rect 2832 6944 2838 6996
rect 3786 6944 3792 6996
rect 3844 6984 3850 6996
rect 4430 6984 4436 6996
rect 3844 6956 4436 6984
rect 3844 6944 3850 6956
rect 4430 6944 4436 6956
rect 4488 6944 4494 6996
rect 5350 6944 5356 6996
rect 5408 6984 5414 6996
rect 5537 6987 5595 6993
rect 5537 6984 5549 6987
rect 5408 6956 5549 6984
rect 5408 6944 5414 6956
rect 5537 6953 5549 6956
rect 5583 6953 5595 6987
rect 5537 6947 5595 6953
rect 5626 6944 5632 6996
rect 5684 6944 5690 6996
rect 6196 6956 6500 6984
rect 1397 6851 1455 6857
rect 1397 6817 1409 6851
rect 1443 6848 1455 6851
rect 2746 6848 2774 6944
rect 3789 6851 3847 6857
rect 3789 6848 3801 6851
rect 1443 6820 3801 6848
rect 1443 6817 1455 6820
rect 1397 6811 1455 6817
rect 3789 6817 3801 6820
rect 3835 6817 3847 6851
rect 3789 6811 3847 6817
rect 4065 6851 4123 6857
rect 4065 6817 4077 6851
rect 4111 6848 4123 6851
rect 4614 6848 4620 6860
rect 4111 6820 4620 6848
rect 4111 6817 4123 6820
rect 4065 6811 4123 6817
rect 4614 6808 4620 6820
rect 4672 6808 4678 6860
rect 5534 6808 5540 6860
rect 5592 6848 5598 6860
rect 5592 6820 6132 6848
rect 5592 6808 5598 6820
rect 3142 6780 3148 6792
rect 2806 6752 3148 6780
rect 3142 6740 3148 6752
rect 3200 6740 3206 6792
rect 3513 6783 3571 6789
rect 3513 6749 3525 6783
rect 3559 6780 3571 6783
rect 3694 6780 3700 6792
rect 3559 6752 3700 6780
rect 3559 6749 3571 6752
rect 3513 6743 3571 6749
rect 3694 6740 3700 6752
rect 3752 6740 3758 6792
rect 5905 6783 5963 6789
rect 5905 6749 5917 6783
rect 5951 6749 5963 6783
rect 5905 6743 5963 6749
rect 3160 6712 3188 6740
rect 4154 6712 4160 6724
rect 3160 6684 4160 6712
rect 4154 6672 4160 6684
rect 4212 6712 4218 6724
rect 4212 6684 4554 6712
rect 4212 6672 4218 6684
rect 5442 6672 5448 6724
rect 5500 6712 5506 6724
rect 5920 6712 5948 6743
rect 5994 6740 6000 6792
rect 6052 6740 6058 6792
rect 6104 6789 6132 6820
rect 6089 6783 6147 6789
rect 6089 6749 6101 6783
rect 6135 6749 6147 6783
rect 6089 6743 6147 6749
rect 6196 6712 6224 6956
rect 6365 6919 6423 6925
rect 6365 6916 6377 6919
rect 6288 6888 6377 6916
rect 6288 6848 6316 6888
rect 6365 6885 6377 6888
rect 6411 6885 6423 6919
rect 6472 6916 6500 6956
rect 6546 6944 6552 6996
rect 6604 6944 6610 6996
rect 6914 6944 6920 6996
rect 6972 6984 6978 6996
rect 7193 6987 7251 6993
rect 7193 6984 7205 6987
rect 6972 6956 7205 6984
rect 6972 6944 6978 6956
rect 7193 6953 7205 6956
rect 7239 6953 7251 6987
rect 7193 6947 7251 6953
rect 7282 6944 7288 6996
rect 7340 6984 7346 6996
rect 7469 6987 7527 6993
rect 7469 6984 7481 6987
rect 7340 6956 7481 6984
rect 7340 6944 7346 6956
rect 7469 6953 7481 6956
rect 7515 6953 7527 6987
rect 7469 6947 7527 6953
rect 6822 6916 6828 6928
rect 6472 6888 6828 6916
rect 6365 6879 6423 6885
rect 6822 6876 6828 6888
rect 6880 6876 6886 6928
rect 8018 6876 8024 6928
rect 8076 6876 8082 6928
rect 8294 6876 8300 6928
rect 8352 6876 8358 6928
rect 6454 6848 6460 6860
rect 6288 6820 6460 6848
rect 6288 6789 6316 6820
rect 6454 6808 6460 6820
rect 6512 6848 6518 6860
rect 7834 6848 7840 6860
rect 6512 6820 7840 6848
rect 6512 6808 6518 6820
rect 7834 6808 7840 6820
rect 7892 6808 7898 6860
rect 8754 6808 8760 6860
rect 8812 6848 8818 6860
rect 8941 6851 8999 6857
rect 8941 6848 8953 6851
rect 8812 6820 8953 6848
rect 8812 6808 8818 6820
rect 8941 6817 8953 6820
rect 8987 6817 8999 6851
rect 8941 6811 8999 6817
rect 6273 6783 6331 6789
rect 6273 6749 6285 6783
rect 6319 6749 6331 6783
rect 6273 6743 6331 6749
rect 6472 6752 6684 6780
rect 5500 6684 5672 6712
rect 5920 6684 6224 6712
rect 5500 6672 5506 6684
rect 2406 6604 2412 6656
rect 2464 6644 2470 6656
rect 3145 6647 3203 6653
rect 3145 6644 3157 6647
rect 2464 6616 3157 6644
rect 2464 6604 2470 6616
rect 3145 6613 3157 6616
rect 3191 6613 3203 6647
rect 3145 6607 3203 6613
rect 3326 6604 3332 6656
rect 3384 6604 3390 6656
rect 5644 6644 5672 6684
rect 6472 6644 6500 6752
rect 6656 6712 6684 6752
rect 6822 6740 6828 6792
rect 6880 6780 6886 6792
rect 6917 6783 6975 6789
rect 6917 6780 6929 6783
rect 6880 6752 6929 6780
rect 6880 6740 6886 6752
rect 6917 6749 6929 6752
rect 6963 6749 6975 6783
rect 6917 6743 6975 6749
rect 7282 6740 7288 6792
rect 7340 6780 7346 6792
rect 8573 6783 8631 6789
rect 8573 6780 8585 6783
rect 7340 6752 8585 6780
rect 7340 6740 7346 6752
rect 8573 6749 8585 6752
rect 8619 6749 8631 6783
rect 8573 6743 8631 6749
rect 9122 6740 9128 6792
rect 9180 6740 9186 6792
rect 7009 6715 7067 6721
rect 7009 6712 7021 6715
rect 6656 6684 7021 6712
rect 7009 6681 7021 6684
rect 7055 6681 7067 6715
rect 7653 6715 7711 6721
rect 7009 6675 7067 6681
rect 7116 6684 7512 6712
rect 6549 6647 6607 6653
rect 6549 6644 6561 6647
rect 5644 6616 6561 6644
rect 6549 6613 6561 6616
rect 6595 6613 6607 6647
rect 6549 6607 6607 6613
rect 6730 6604 6736 6656
rect 6788 6644 6794 6656
rect 7116 6644 7144 6684
rect 6788 6616 7144 6644
rect 6788 6604 6794 6616
rect 7190 6604 7196 6656
rect 7248 6653 7254 6656
rect 7248 6647 7267 6653
rect 7255 6613 7267 6647
rect 7248 6607 7267 6613
rect 7248 6604 7254 6607
rect 7374 6604 7380 6656
rect 7432 6604 7438 6656
rect 7484 6644 7512 6684
rect 7653 6681 7665 6715
rect 7699 6712 7711 6715
rect 9030 6712 9036 6724
rect 7699 6684 9036 6712
rect 7699 6681 7711 6684
rect 7653 6675 7711 6681
rect 9030 6672 9036 6684
rect 9088 6712 9094 6724
rect 9309 6715 9367 6721
rect 9309 6712 9321 6715
rect 9088 6684 9321 6712
rect 9088 6672 9094 6684
rect 9309 6681 9321 6684
rect 9355 6681 9367 6715
rect 9309 6675 9367 6681
rect 7745 6647 7803 6653
rect 7745 6644 7757 6647
rect 7484 6616 7757 6644
rect 7745 6613 7757 6616
rect 7791 6613 7803 6647
rect 7745 6607 7803 6613
rect 7834 6604 7840 6656
rect 7892 6604 7898 6656
rect 8110 6604 8116 6656
rect 8168 6604 8174 6656
rect 1104 6554 10488 6576
rect 1104 6502 4874 6554
rect 4926 6502 4938 6554
rect 4990 6502 5002 6554
rect 5054 6502 5066 6554
rect 5118 6502 5130 6554
rect 5182 6502 10488 6554
rect 1104 6480 10488 6502
rect 2774 6400 2780 6452
rect 2832 6400 2838 6452
rect 2958 6400 2964 6452
rect 3016 6440 3022 6452
rect 4617 6443 4675 6449
rect 3016 6412 3188 6440
rect 3016 6400 3022 6412
rect 2314 6372 2320 6384
rect 1688 6344 2320 6372
rect 1578 6264 1584 6316
rect 1636 6264 1642 6316
rect 1688 6313 1716 6344
rect 2314 6332 2320 6344
rect 2372 6332 2378 6384
rect 2792 6372 2820 6400
rect 3160 6381 3188 6412
rect 4617 6409 4629 6443
rect 4663 6440 4675 6443
rect 4706 6440 4712 6452
rect 4663 6412 4712 6440
rect 4663 6409 4675 6412
rect 4617 6403 4675 6409
rect 4706 6400 4712 6412
rect 4764 6400 4770 6452
rect 6270 6440 6276 6452
rect 5092 6412 6276 6440
rect 3145 6375 3203 6381
rect 2792 6344 2912 6372
rect 2884 6313 2912 6344
rect 3145 6341 3157 6375
rect 3191 6341 3203 6375
rect 3145 6335 3203 6341
rect 4154 6332 4160 6384
rect 4212 6332 4218 6384
rect 4430 6332 4436 6384
rect 4488 6372 4494 6384
rect 5092 6381 5120 6412
rect 6270 6400 6276 6412
rect 6328 6400 6334 6452
rect 6365 6443 6423 6449
rect 6365 6409 6377 6443
rect 6411 6440 6423 6443
rect 6546 6440 6552 6452
rect 6411 6412 6552 6440
rect 6411 6409 6423 6412
rect 6365 6403 6423 6409
rect 6546 6400 6552 6412
rect 6604 6400 6610 6452
rect 6638 6400 6644 6452
rect 6696 6440 6702 6452
rect 6696 6412 7696 6440
rect 6696 6400 6702 6412
rect 4861 6375 4919 6381
rect 4861 6372 4873 6375
rect 4488 6344 4873 6372
rect 4488 6332 4494 6344
rect 4861 6341 4873 6344
rect 4907 6341 4919 6375
rect 4861 6335 4919 6341
rect 5077 6375 5135 6381
rect 5077 6341 5089 6375
rect 5123 6341 5135 6375
rect 5902 6372 5908 6384
rect 5077 6335 5135 6341
rect 5184 6344 5908 6372
rect 1673 6307 1731 6313
rect 1673 6273 1685 6307
rect 1719 6273 1731 6307
rect 1673 6267 1731 6273
rect 1857 6307 1915 6313
rect 1857 6273 1869 6307
rect 1903 6304 1915 6307
rect 2869 6307 2927 6313
rect 1903 6276 2636 6304
rect 1903 6273 1915 6276
rect 1857 6267 1915 6273
rect 1762 6196 1768 6248
rect 1820 6196 1826 6248
rect 1854 6128 1860 6180
rect 1912 6168 1918 6180
rect 2133 6171 2191 6177
rect 2133 6168 2145 6171
rect 1912 6140 2145 6168
rect 1912 6128 1918 6140
rect 2133 6137 2145 6140
rect 2179 6137 2191 6171
rect 2133 6131 2191 6137
rect 2038 6060 2044 6112
rect 2096 6060 2102 6112
rect 2608 6100 2636 6276
rect 2869 6273 2881 6307
rect 2915 6273 2927 6307
rect 2869 6267 2927 6273
rect 2777 6239 2835 6245
rect 2777 6205 2789 6239
rect 2823 6236 2835 6239
rect 3142 6236 3148 6248
rect 2823 6208 3148 6236
rect 2823 6205 2835 6208
rect 2777 6199 2835 6205
rect 3142 6196 3148 6208
rect 3200 6196 3206 6248
rect 3786 6196 3792 6248
rect 3844 6236 3850 6248
rect 5092 6236 5120 6335
rect 3844 6208 5120 6236
rect 3844 6196 3850 6208
rect 4709 6171 4767 6177
rect 4709 6137 4721 6171
rect 4755 6168 4767 6171
rect 4798 6168 4804 6180
rect 4755 6140 4804 6168
rect 4755 6137 4767 6140
rect 4709 6131 4767 6137
rect 4798 6128 4804 6140
rect 4856 6128 4862 6180
rect 3878 6100 3884 6112
rect 2608 6072 3884 6100
rect 3878 6060 3884 6072
rect 3936 6100 3942 6112
rect 4893 6103 4951 6109
rect 4893 6100 4905 6103
rect 3936 6072 4905 6100
rect 3936 6060 3942 6072
rect 4893 6069 4905 6072
rect 4939 6100 4951 6103
rect 5184 6100 5212 6344
rect 5902 6332 5908 6344
rect 5960 6372 5966 6384
rect 6730 6372 6736 6384
rect 5960 6344 6736 6372
rect 5960 6332 5966 6344
rect 6730 6332 6736 6344
rect 6788 6332 6794 6384
rect 7101 6375 7159 6381
rect 7101 6341 7113 6375
rect 7147 6372 7159 6375
rect 7147 6344 7328 6372
rect 7147 6341 7159 6344
rect 7101 6335 7159 6341
rect 7300 6316 7328 6344
rect 5350 6264 5356 6316
rect 5408 6304 5414 6316
rect 5813 6307 5871 6313
rect 5813 6304 5825 6307
rect 5408 6276 5825 6304
rect 5408 6264 5414 6276
rect 5813 6273 5825 6276
rect 5859 6273 5871 6307
rect 5813 6267 5871 6273
rect 5828 6168 5856 6267
rect 6178 6264 6184 6316
rect 6236 6304 6242 6316
rect 6549 6307 6607 6313
rect 6549 6304 6561 6307
rect 6236 6276 6561 6304
rect 6236 6264 6242 6276
rect 6549 6273 6561 6276
rect 6595 6304 6607 6307
rect 7190 6304 7196 6316
rect 6595 6276 7196 6304
rect 6595 6273 6607 6276
rect 6549 6267 6607 6273
rect 7190 6264 7196 6276
rect 7248 6264 7254 6316
rect 7282 6264 7288 6316
rect 7340 6264 7346 6316
rect 7668 6313 7696 6412
rect 8110 6400 8116 6452
rect 8168 6400 8174 6452
rect 7469 6307 7527 6313
rect 7469 6273 7481 6307
rect 7515 6273 7527 6307
rect 7469 6267 7527 6273
rect 7561 6307 7619 6313
rect 7561 6273 7573 6307
rect 7607 6273 7619 6307
rect 7561 6267 7619 6273
rect 7653 6307 7711 6313
rect 7653 6273 7665 6307
rect 7699 6273 7711 6307
rect 8021 6307 8079 6313
rect 8021 6304 8033 6307
rect 7653 6267 7711 6273
rect 7944 6276 8033 6304
rect 6641 6239 6699 6245
rect 6641 6205 6653 6239
rect 6687 6236 6699 6239
rect 6914 6236 6920 6248
rect 6687 6208 6920 6236
rect 6687 6205 6699 6208
rect 6641 6199 6699 6205
rect 6914 6196 6920 6208
rect 6972 6196 6978 6248
rect 7484 6236 7512 6267
rect 7116 6208 7512 6236
rect 7116 6180 7144 6208
rect 6822 6168 6828 6180
rect 5828 6140 6828 6168
rect 6822 6128 6828 6140
rect 6880 6128 6886 6180
rect 7098 6128 7104 6180
rect 7156 6128 7162 6180
rect 7374 6168 7380 6180
rect 7208 6140 7380 6168
rect 4939 6072 5212 6100
rect 4939 6069 4951 6072
rect 4893 6063 4951 6069
rect 5258 6060 5264 6112
rect 5316 6060 5322 6112
rect 6730 6060 6736 6112
rect 6788 6100 6794 6112
rect 7208 6100 7236 6140
rect 7374 6128 7380 6140
rect 7432 6168 7438 6180
rect 7576 6168 7604 6267
rect 7432 6140 7604 6168
rect 7432 6128 7438 6140
rect 6788 6072 7236 6100
rect 6788 6060 6794 6072
rect 7282 6060 7288 6112
rect 7340 6100 7346 6112
rect 7944 6109 7972 6276
rect 8021 6273 8033 6276
rect 8067 6273 8079 6307
rect 8128 6304 8156 6400
rect 8205 6307 8263 6313
rect 8205 6304 8217 6307
rect 8128 6276 8217 6304
rect 8021 6267 8079 6273
rect 8205 6273 8217 6276
rect 8251 6273 8263 6307
rect 8205 6267 8263 6273
rect 7929 6103 7987 6109
rect 7929 6100 7941 6103
rect 7340 6072 7941 6100
rect 7340 6060 7346 6072
rect 7929 6069 7941 6072
rect 7975 6069 7987 6103
rect 7929 6063 7987 6069
rect 8205 6103 8263 6109
rect 8205 6069 8217 6103
rect 8251 6100 8263 6103
rect 8386 6100 8392 6112
rect 8251 6072 8392 6100
rect 8251 6069 8263 6072
rect 8205 6063 8263 6069
rect 8386 6060 8392 6072
rect 8444 6060 8450 6112
rect 1104 6010 10488 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 10488 6010
rect 1104 5936 10488 5958
rect 1660 5899 1718 5905
rect 1660 5865 1672 5899
rect 1706 5896 1718 5899
rect 1854 5896 1860 5908
rect 1706 5868 1860 5896
rect 1706 5865 1718 5868
rect 1660 5859 1718 5865
rect 1854 5856 1860 5868
rect 1912 5856 1918 5908
rect 2038 5856 2044 5908
rect 2096 5896 2102 5908
rect 2096 5868 3280 5896
rect 2096 5856 2102 5868
rect 2774 5828 2780 5840
rect 2746 5788 2780 5828
rect 2832 5788 2838 5840
rect 1397 5763 1455 5769
rect 1397 5729 1409 5763
rect 1443 5760 1455 5763
rect 2746 5760 2774 5788
rect 1443 5732 2774 5760
rect 1443 5729 1455 5732
rect 1397 5723 1455 5729
rect 3252 5701 3280 5868
rect 3418 5856 3424 5908
rect 3476 5856 3482 5908
rect 3786 5856 3792 5908
rect 3844 5896 3850 5908
rect 3970 5896 3976 5908
rect 3844 5868 3976 5896
rect 3844 5856 3850 5868
rect 3970 5856 3976 5868
rect 4028 5856 4034 5908
rect 4341 5899 4399 5905
rect 4341 5865 4353 5899
rect 4387 5896 4399 5899
rect 4614 5896 4620 5908
rect 4387 5868 4620 5896
rect 4387 5865 4399 5868
rect 4341 5859 4399 5865
rect 4614 5856 4620 5868
rect 4672 5856 4678 5908
rect 5258 5856 5264 5908
rect 5316 5856 5322 5908
rect 5442 5856 5448 5908
rect 5500 5856 5506 5908
rect 7009 5899 7067 5905
rect 7009 5865 7021 5899
rect 7055 5896 7067 5899
rect 7190 5896 7196 5908
rect 7055 5868 7196 5896
rect 7055 5865 7067 5868
rect 7009 5859 7067 5865
rect 7190 5856 7196 5868
rect 7248 5856 7254 5908
rect 8386 5856 8392 5908
rect 8444 5896 8450 5908
rect 8493 5899 8551 5905
rect 8493 5896 8505 5899
rect 8444 5868 8505 5896
rect 8444 5856 8450 5868
rect 8493 5865 8505 5868
rect 8539 5865 8551 5899
rect 8493 5859 8551 5865
rect 3712 5800 5212 5828
rect 3237 5695 3295 5701
rect 3237 5661 3249 5695
rect 3283 5661 3295 5695
rect 3712 5692 3740 5800
rect 5184 5772 5212 5800
rect 3789 5763 3847 5769
rect 3789 5729 3801 5763
rect 3835 5760 3847 5763
rect 4893 5763 4951 5769
rect 4893 5760 4905 5763
rect 3835 5732 4905 5760
rect 3835 5729 3847 5732
rect 3789 5723 3847 5729
rect 4893 5729 4905 5732
rect 4939 5729 4951 5763
rect 4893 5723 4951 5729
rect 5166 5720 5172 5772
rect 5224 5720 5230 5772
rect 3881 5695 3939 5701
rect 3881 5692 3893 5695
rect 3712 5664 3893 5692
rect 3237 5655 3295 5661
rect 3881 5661 3893 5664
rect 3927 5661 3939 5695
rect 3881 5655 3939 5661
rect 4249 5695 4307 5701
rect 4249 5661 4261 5695
rect 4295 5692 4307 5695
rect 5276 5692 5304 5856
rect 5460 5692 5488 5856
rect 6928 5763 6986 5769
rect 6928 5729 6940 5763
rect 6974 5760 6986 5763
rect 8478 5760 8484 5772
rect 6974 5732 8484 5760
rect 6974 5729 6986 5732
rect 6928 5723 6986 5729
rect 8478 5720 8484 5732
rect 8536 5760 8542 5772
rect 8757 5763 8815 5769
rect 8757 5760 8769 5763
rect 8536 5732 8769 5760
rect 8536 5720 8542 5732
rect 8757 5729 8769 5732
rect 8803 5729 8815 5763
rect 8757 5723 8815 5729
rect 4295 5664 5304 5692
rect 5368 5664 5488 5692
rect 10137 5695 10195 5701
rect 4295 5661 4307 5664
rect 4249 5655 4307 5661
rect 2314 5584 2320 5636
rect 2372 5584 2378 5636
rect 4614 5624 4620 5636
rect 3160 5596 4620 5624
rect 3160 5565 3188 5596
rect 4614 5584 4620 5596
rect 4672 5584 4678 5636
rect 5368 5624 5396 5664
rect 10137 5661 10149 5695
rect 10183 5661 10195 5695
rect 10137 5655 10195 5661
rect 5092 5596 5396 5624
rect 3145 5559 3203 5565
rect 3145 5525 3157 5559
rect 3191 5525 3203 5559
rect 3145 5519 3203 5525
rect 4157 5559 4215 5565
rect 4157 5525 4169 5559
rect 4203 5556 4215 5559
rect 4338 5556 4344 5568
rect 4203 5528 4344 5556
rect 4203 5525 4215 5528
rect 4157 5519 4215 5525
rect 4338 5516 4344 5528
rect 4396 5556 4402 5568
rect 4798 5556 4804 5568
rect 4396 5528 4804 5556
rect 4396 5516 4402 5528
rect 4798 5516 4804 5528
rect 4856 5556 4862 5568
rect 5092 5556 5120 5596
rect 6086 5584 6092 5636
rect 6144 5584 6150 5636
rect 6638 5584 6644 5636
rect 6696 5584 6702 5636
rect 7742 5584 7748 5636
rect 7800 5584 7806 5636
rect 10152 5624 10180 5655
rect 10502 5624 10508 5636
rect 10152 5596 10508 5624
rect 10502 5584 10508 5596
rect 10560 5584 10566 5636
rect 4856 5528 5120 5556
rect 5169 5559 5227 5565
rect 4856 5516 4862 5528
rect 5169 5525 5181 5559
rect 5215 5556 5227 5559
rect 6270 5556 6276 5568
rect 5215 5528 6276 5556
rect 5215 5525 5227 5528
rect 5169 5519 5227 5525
rect 6270 5516 6276 5528
rect 6328 5556 6334 5568
rect 7098 5556 7104 5568
rect 6328 5528 7104 5556
rect 6328 5516 6334 5528
rect 7098 5516 7104 5528
rect 7156 5516 7162 5568
rect 7466 5516 7472 5568
rect 7524 5556 7530 5568
rect 9953 5559 10011 5565
rect 9953 5556 9965 5559
rect 7524 5528 9965 5556
rect 7524 5516 7530 5528
rect 9953 5525 9965 5528
rect 9999 5525 10011 5559
rect 9953 5519 10011 5525
rect 1104 5466 10488 5488
rect 1104 5414 4874 5466
rect 4926 5414 4938 5466
rect 4990 5414 5002 5466
rect 5054 5414 5066 5466
rect 5118 5414 5130 5466
rect 5182 5414 10488 5466
rect 1104 5392 10488 5414
rect 1762 5312 1768 5364
rect 1820 5352 1826 5364
rect 1949 5355 2007 5361
rect 1949 5352 1961 5355
rect 1820 5324 1961 5352
rect 1820 5312 1826 5324
rect 1949 5321 1961 5324
rect 1995 5321 2007 5355
rect 2774 5352 2780 5364
rect 1949 5315 2007 5321
rect 2608 5324 2780 5352
rect 1118 5244 1124 5296
rect 1176 5284 1182 5296
rect 1176 5256 2176 5284
rect 1176 5244 1182 5256
rect 1394 5176 1400 5228
rect 1452 5176 1458 5228
rect 2148 5225 2176 5256
rect 2608 5225 2636 5324
rect 2774 5312 2780 5324
rect 2832 5352 2838 5364
rect 2832 5324 4476 5352
rect 2832 5312 2838 5324
rect 4448 5225 4476 5324
rect 6178 5312 6184 5364
rect 6236 5312 6242 5364
rect 6270 5312 6276 5364
rect 6328 5312 6334 5364
rect 6365 5355 6423 5361
rect 6365 5321 6377 5355
rect 6411 5352 6423 5355
rect 6638 5352 6644 5364
rect 6411 5324 6644 5352
rect 6411 5321 6423 5324
rect 6365 5315 6423 5321
rect 6638 5312 6644 5324
rect 6696 5312 6702 5364
rect 7558 5352 7564 5364
rect 7024 5324 7564 5352
rect 1857 5219 1915 5225
rect 1857 5216 1869 5219
rect 1596 5188 1869 5216
rect 1596 5089 1624 5188
rect 1857 5185 1869 5188
rect 1903 5185 1915 5219
rect 1857 5179 1915 5185
rect 2133 5219 2191 5225
rect 2133 5185 2145 5219
rect 2179 5185 2191 5219
rect 2133 5179 2191 5185
rect 2593 5219 2651 5225
rect 2593 5185 2605 5219
rect 2639 5185 2651 5219
rect 4433 5219 4491 5225
rect 2593 5179 2651 5185
rect 2869 5151 2927 5157
rect 2869 5117 2881 5151
rect 2915 5148 2927 5151
rect 3326 5148 3332 5160
rect 2915 5120 3332 5148
rect 2915 5117 2927 5120
rect 2869 5111 2927 5117
rect 3326 5108 3332 5120
rect 3384 5108 3390 5160
rect 3988 5148 4016 5202
rect 4433 5185 4445 5219
rect 4479 5185 4491 5219
rect 6288 5216 6316 5312
rect 7024 5225 7052 5324
rect 7558 5312 7564 5324
rect 7616 5312 7622 5364
rect 7742 5312 7748 5364
rect 7800 5352 7806 5364
rect 7800 5324 8248 5352
rect 7800 5312 7806 5324
rect 8220 5284 8248 5324
rect 8478 5312 8484 5364
rect 8536 5312 8542 5364
rect 8142 5256 8248 5284
rect 8496 5284 8524 5312
rect 8496 5256 8892 5284
rect 8864 5225 8892 5256
rect 6549 5219 6607 5225
rect 6549 5216 6561 5219
rect 4433 5179 4491 5185
rect 4062 5148 4068 5160
rect 3988 5120 4068 5148
rect 4062 5108 4068 5120
rect 4120 5108 4126 5160
rect 4706 5108 4712 5160
rect 4764 5108 4770 5160
rect 5828 5148 5856 5202
rect 6288 5188 6561 5216
rect 6549 5185 6561 5188
rect 6595 5185 6607 5219
rect 6549 5179 6607 5185
rect 6825 5219 6883 5225
rect 6825 5185 6837 5219
rect 6871 5185 6883 5219
rect 6825 5179 6883 5185
rect 7009 5219 7067 5225
rect 7009 5185 7021 5219
rect 7055 5185 7067 5219
rect 7009 5179 7067 5185
rect 8849 5219 8907 5225
rect 8849 5185 8861 5219
rect 8895 5185 8907 5219
rect 8849 5179 8907 5185
rect 6086 5148 6092 5160
rect 5828 5120 6092 5148
rect 6086 5108 6092 5120
rect 6144 5108 6150 5160
rect 1581 5083 1639 5089
rect 1581 5049 1593 5083
rect 1627 5049 1639 5083
rect 1581 5043 1639 5049
rect 4338 5040 4344 5092
rect 4396 5040 4402 5092
rect 2314 4972 2320 5024
rect 2372 4972 2378 5024
rect 6104 5012 6132 5108
rect 6840 5092 6868 5179
rect 6914 5108 6920 5160
rect 6972 5148 6978 5160
rect 7101 5151 7159 5157
rect 7101 5148 7113 5151
rect 6972 5120 7113 5148
rect 6972 5108 6978 5120
rect 7101 5117 7113 5120
rect 7147 5117 7159 5151
rect 8202 5148 8208 5160
rect 7101 5111 7159 5117
rect 7208 5120 8208 5148
rect 6362 5040 6368 5092
rect 6420 5080 6426 5092
rect 6638 5080 6644 5092
rect 6420 5052 6644 5080
rect 6420 5040 6426 5052
rect 6638 5040 6644 5052
rect 6696 5040 6702 5092
rect 6730 5040 6736 5092
rect 6788 5040 6794 5092
rect 6822 5040 6828 5092
rect 6880 5080 6886 5092
rect 7208 5080 7236 5120
rect 8202 5108 8208 5120
rect 8260 5108 8266 5160
rect 8570 5108 8576 5160
rect 8628 5108 8634 5160
rect 6880 5052 7236 5080
rect 6880 5040 6886 5052
rect 7558 5040 7564 5092
rect 7616 5040 7622 5092
rect 7576 5012 7604 5040
rect 6104 4984 7604 5012
rect 1104 4922 10488 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 10488 4922
rect 1104 4848 10488 4870
rect 2774 4808 2780 4820
rect 2746 4768 2780 4808
rect 2832 4768 2838 4820
rect 3142 4768 3148 4820
rect 3200 4768 3206 4820
rect 3326 4768 3332 4820
rect 3384 4808 3390 4820
rect 3789 4811 3847 4817
rect 3789 4808 3801 4811
rect 3384 4780 3801 4808
rect 3384 4768 3390 4780
rect 3789 4777 3801 4780
rect 3835 4777 3847 4811
rect 3789 4771 3847 4777
rect 3970 4768 3976 4820
rect 4028 4768 4034 4820
rect 4706 4768 4712 4820
rect 4764 4808 4770 4820
rect 5445 4811 5503 4817
rect 5445 4808 5457 4811
rect 4764 4780 5457 4808
rect 4764 4768 4770 4780
rect 5445 4777 5457 4780
rect 5491 4777 5503 4811
rect 5445 4771 5503 4777
rect 6822 4768 6828 4820
rect 6880 4768 6886 4820
rect 6914 4768 6920 4820
rect 6972 4768 6978 4820
rect 7926 4768 7932 4820
rect 7984 4808 7990 4820
rect 8021 4811 8079 4817
rect 8021 4808 8033 4811
rect 7984 4780 8033 4808
rect 7984 4768 7990 4780
rect 8021 4777 8033 4780
rect 8067 4777 8079 4811
rect 8021 4771 8079 4777
rect 1397 4675 1455 4681
rect 1397 4641 1409 4675
rect 1443 4672 1455 4675
rect 2746 4672 2774 4768
rect 4798 4700 4804 4752
rect 4856 4700 4862 4752
rect 6730 4740 6736 4752
rect 5460 4712 6736 4740
rect 1443 4644 2774 4672
rect 4525 4675 4583 4681
rect 1443 4641 1455 4644
rect 1397 4635 1455 4641
rect 4525 4641 4537 4675
rect 4571 4672 4583 4675
rect 4614 4672 4620 4684
rect 4571 4644 4620 4672
rect 4571 4641 4583 4644
rect 4525 4635 4583 4641
rect 4614 4632 4620 4644
rect 4672 4632 4678 4684
rect 4065 4607 4123 4613
rect 4065 4573 4077 4607
rect 4111 4573 4123 4607
rect 4065 4567 4123 4573
rect 4341 4607 4399 4613
rect 4341 4573 4353 4607
rect 4387 4604 4399 4607
rect 4816 4604 4844 4700
rect 5460 4613 5488 4712
rect 6730 4700 6736 4712
rect 6788 4700 6794 4752
rect 6932 4740 6960 4768
rect 6932 4712 7696 4740
rect 6178 4632 6184 4684
rect 6236 4672 6242 4684
rect 6457 4675 6515 4681
rect 6457 4672 6469 4675
rect 6236 4644 6469 4672
rect 6236 4632 6242 4644
rect 6457 4641 6469 4644
rect 6503 4641 6515 4675
rect 6457 4635 6515 4641
rect 6917 4675 6975 4681
rect 6917 4641 6929 4675
rect 6963 4672 6975 4675
rect 7098 4672 7104 4684
rect 6963 4644 7104 4672
rect 6963 4641 6975 4644
rect 6917 4635 6975 4641
rect 7098 4632 7104 4644
rect 7156 4632 7162 4684
rect 7668 4681 7696 4712
rect 7653 4675 7711 4681
rect 7653 4641 7665 4675
rect 7699 4641 7711 4675
rect 7653 4635 7711 4641
rect 4387 4576 4844 4604
rect 5169 4607 5227 4613
rect 4387 4573 4399 4576
rect 4341 4567 4399 4573
rect 5169 4573 5181 4607
rect 5215 4573 5227 4607
rect 5169 4567 5227 4573
rect 5445 4607 5503 4613
rect 5445 4573 5457 4607
rect 5491 4573 5503 4607
rect 5445 4567 5503 4573
rect 1670 4496 1676 4548
rect 1728 4496 1734 4548
rect 2314 4496 2320 4548
rect 2372 4496 2378 4548
rect 4080 4536 4108 4567
rect 5184 4536 5212 4567
rect 5534 4564 5540 4616
rect 5592 4604 5598 4616
rect 5629 4607 5687 4613
rect 5629 4604 5641 4607
rect 5592 4576 5641 4604
rect 5592 4564 5598 4576
rect 5629 4573 5641 4576
rect 5675 4573 5687 4607
rect 5629 4567 5687 4573
rect 6638 4564 6644 4616
rect 6696 4564 6702 4616
rect 7834 4564 7840 4616
rect 7892 4564 7898 4616
rect 6656 4536 6684 4564
rect 4080 4508 6684 4536
rect 4430 4428 4436 4480
rect 4488 4468 4494 4480
rect 5077 4471 5135 4477
rect 5077 4468 5089 4471
rect 4488 4440 5089 4468
rect 4488 4428 4494 4440
rect 5077 4437 5089 4440
rect 5123 4437 5135 4471
rect 5077 4431 5135 4437
rect 5902 4428 5908 4480
rect 5960 4428 5966 4480
rect 7098 4428 7104 4480
rect 7156 4428 7162 4480
rect 1104 4378 10488 4400
rect 1104 4326 4874 4378
rect 4926 4326 4938 4378
rect 4990 4326 5002 4378
rect 5054 4326 5066 4378
rect 5118 4326 5130 4378
rect 5182 4326 10488 4378
rect 1104 4304 10488 4326
rect 1670 4224 1676 4276
rect 1728 4264 1734 4276
rect 1765 4267 1823 4273
rect 1765 4264 1777 4267
rect 1728 4236 1777 4264
rect 1728 4224 1734 4236
rect 1765 4233 1777 4236
rect 1811 4233 1823 4267
rect 1765 4227 1823 4233
rect 4062 4224 4068 4276
rect 4120 4264 4126 4276
rect 4157 4267 4215 4273
rect 4157 4264 4169 4267
rect 4120 4236 4169 4264
rect 4120 4224 4126 4236
rect 4157 4233 4169 4236
rect 4203 4233 4215 4267
rect 4157 4227 4215 4233
rect 4798 4224 4804 4276
rect 4856 4264 4862 4276
rect 5261 4267 5319 4273
rect 5261 4264 5273 4267
rect 4856 4236 5273 4264
rect 4856 4224 4862 4236
rect 5261 4233 5273 4236
rect 5307 4233 5319 4267
rect 5261 4227 5319 4233
rect 5902 4224 5908 4276
rect 5960 4224 5966 4276
rect 7098 4224 7104 4276
rect 7156 4224 7162 4276
rect 4430 4156 4436 4208
rect 4488 4196 4494 4208
rect 5445 4199 5503 4205
rect 4488 4168 5396 4196
rect 4488 4156 4494 4168
rect 1673 4131 1731 4137
rect 1673 4097 1685 4131
rect 1719 4097 1731 4131
rect 1673 4091 1731 4097
rect 1688 4060 1716 4091
rect 2038 4088 2044 4140
rect 2096 4088 2102 4140
rect 5169 4131 5227 4137
rect 5169 4097 5181 4131
rect 5215 4097 5227 4131
rect 5368 4128 5396 4168
rect 5445 4165 5457 4199
rect 5491 4196 5503 4199
rect 5920 4196 5948 4224
rect 5491 4168 5948 4196
rect 5491 4165 5503 4168
rect 5445 4159 5503 4165
rect 5629 4131 5687 4137
rect 5629 4128 5641 4131
rect 5368 4100 5641 4128
rect 5169 4091 5227 4097
rect 5629 4097 5641 4100
rect 5675 4097 5687 4131
rect 5629 4091 5687 4097
rect 7009 4131 7067 4137
rect 7009 4097 7021 4131
rect 7055 4128 7067 4131
rect 7116 4128 7144 4224
rect 7055 4100 7144 4128
rect 7055 4097 7067 4100
rect 7009 4091 7067 4097
rect 2133 4063 2191 4069
rect 2133 4060 2145 4063
rect 1688 4032 2145 4060
rect 2133 4029 2145 4032
rect 2179 4029 2191 4063
rect 5184 4060 5212 4091
rect 5350 4060 5356 4072
rect 5184 4032 5356 4060
rect 2133 4023 2191 4029
rect 5350 4020 5356 4032
rect 5408 4020 5414 4072
rect 6086 4060 6092 4072
rect 5828 4032 6092 4060
rect 1486 3952 1492 4004
rect 1544 3952 1550 4004
rect 5445 3995 5503 4001
rect 5445 3961 5457 3995
rect 5491 3992 5503 3995
rect 5534 3992 5540 4004
rect 5491 3964 5540 3992
rect 5491 3961 5503 3964
rect 5445 3955 5503 3961
rect 5534 3952 5540 3964
rect 5592 3952 5598 4004
rect 5828 4001 5856 4032
rect 6086 4020 6092 4032
rect 6144 4020 6150 4072
rect 7101 4063 7159 4069
rect 7101 4029 7113 4063
rect 7147 4060 7159 4063
rect 7282 4060 7288 4072
rect 7147 4032 7288 4060
rect 7147 4029 7159 4032
rect 7101 4023 7159 4029
rect 7282 4020 7288 4032
rect 7340 4020 7346 4072
rect 7377 4063 7435 4069
rect 7377 4029 7389 4063
rect 7423 4060 7435 4063
rect 8570 4060 8576 4072
rect 7423 4032 8576 4060
rect 7423 4029 7435 4032
rect 7377 4023 7435 4029
rect 8570 4020 8576 4032
rect 8628 4020 8634 4072
rect 5813 3995 5871 4001
rect 5813 3961 5825 3995
rect 5859 3961 5871 3995
rect 5813 3955 5871 3961
rect 1104 3834 10488 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 10488 3834
rect 1104 3760 10488 3782
rect 1581 3723 1639 3729
rect 1581 3689 1593 3723
rect 1627 3720 1639 3723
rect 2038 3720 2044 3732
rect 1627 3692 2044 3720
rect 1627 3689 1639 3692
rect 1581 3683 1639 3689
rect 2038 3680 2044 3692
rect 2096 3680 2102 3732
rect 5537 3723 5595 3729
rect 5537 3689 5549 3723
rect 5583 3720 5595 3723
rect 5583 3692 5764 3720
rect 5583 3689 5595 3692
rect 5537 3683 5595 3689
rect 5736 3596 5764 3692
rect 5718 3544 5724 3596
rect 5776 3584 5782 3596
rect 5997 3587 6055 3593
rect 5997 3584 6009 3587
rect 5776 3556 6009 3584
rect 5776 3544 5782 3556
rect 5997 3553 6009 3556
rect 6043 3553 6055 3587
rect 5997 3547 6055 3553
rect 934 3476 940 3528
rect 992 3516 998 3528
rect 1397 3519 1455 3525
rect 1397 3516 1409 3519
rect 992 3488 1409 3516
rect 992 3476 998 3488
rect 1397 3485 1409 3488
rect 1443 3485 1455 3519
rect 1397 3479 1455 3485
rect 3970 3476 3976 3528
rect 4028 3476 4034 3528
rect 4614 3476 4620 3528
rect 4672 3476 4678 3528
rect 5902 3516 5908 3528
rect 5536 3491 5908 3516
rect 5491 3488 5908 3491
rect 5491 3485 5564 3488
rect 5491 3451 5503 3485
rect 5537 3454 5564 3485
rect 5902 3476 5908 3488
rect 5960 3516 5966 3528
rect 6089 3519 6147 3525
rect 6089 3516 6101 3519
rect 5960 3488 6101 3516
rect 5960 3476 5966 3488
rect 6089 3485 6101 3488
rect 6135 3485 6147 3519
rect 6089 3479 6147 3485
rect 5537 3451 5549 3454
rect 5491 3445 5549 3451
rect 5721 3451 5779 3457
rect 5721 3417 5733 3451
rect 5767 3448 5779 3451
rect 5813 3451 5871 3457
rect 5813 3448 5825 3451
rect 5767 3420 5825 3448
rect 5767 3417 5779 3420
rect 5721 3411 5779 3417
rect 5813 3417 5825 3420
rect 5859 3448 5871 3451
rect 5994 3448 6000 3460
rect 5859 3420 6000 3448
rect 5859 3417 5871 3420
rect 5813 3411 5871 3417
rect 5994 3408 6000 3420
rect 6052 3408 6058 3460
rect 3878 3340 3884 3392
rect 3936 3380 3942 3392
rect 4157 3383 4215 3389
rect 4157 3380 4169 3383
rect 3936 3352 4169 3380
rect 3936 3340 3942 3352
rect 4157 3349 4169 3352
rect 4203 3349 4215 3383
rect 4157 3343 4215 3349
rect 4798 3340 4804 3392
rect 4856 3340 4862 3392
rect 5350 3340 5356 3392
rect 5408 3340 5414 3392
rect 6086 3340 6092 3392
rect 6144 3340 6150 3392
rect 1104 3290 10488 3312
rect 1104 3238 4874 3290
rect 4926 3238 4938 3290
rect 4990 3238 5002 3290
rect 5054 3238 5066 3290
rect 5118 3238 5130 3290
rect 5182 3238 10488 3290
rect 1104 3216 10488 3238
rect 3697 3179 3755 3185
rect 3697 3145 3709 3179
rect 3743 3176 3755 3179
rect 3970 3176 3976 3188
rect 3743 3148 3976 3176
rect 3743 3145 3755 3148
rect 3697 3139 3755 3145
rect 3970 3136 3976 3148
rect 4028 3136 4034 3188
rect 4614 3136 4620 3188
rect 4672 3176 4678 3188
rect 4709 3179 4767 3185
rect 4709 3176 4721 3179
rect 4672 3148 4721 3176
rect 4672 3136 4678 3148
rect 4709 3145 4721 3148
rect 4755 3145 4767 3179
rect 4709 3139 4767 3145
rect 5902 3136 5908 3188
rect 5960 3176 5966 3188
rect 6181 3179 6239 3185
rect 5960 3148 6132 3176
rect 5960 3136 5966 3148
rect 4356 3080 4568 3108
rect 4065 3043 4123 3049
rect 4065 3009 4077 3043
rect 4111 3040 4123 3043
rect 4356 3040 4384 3080
rect 4111 3012 4384 3040
rect 4111 3009 4123 3012
rect 4065 3003 4123 3009
rect 4430 3000 4436 3052
rect 4488 3000 4494 3052
rect 4540 3049 4568 3080
rect 4525 3043 4583 3049
rect 4525 3009 4537 3043
rect 4571 3040 4583 3043
rect 4985 3043 5043 3049
rect 4985 3040 4997 3043
rect 4571 3012 4997 3040
rect 4571 3009 4583 3012
rect 4525 3003 4583 3009
rect 4985 3009 4997 3012
rect 5031 3040 5043 3043
rect 5920 3040 5948 3136
rect 5994 3068 6000 3120
rect 6052 3068 6058 3120
rect 6104 3108 6132 3148
rect 6181 3145 6193 3179
rect 6227 3176 6239 3179
rect 7282 3176 7288 3188
rect 6227 3148 7288 3176
rect 6227 3145 6239 3148
rect 6181 3139 6239 3145
rect 7282 3136 7288 3148
rect 7340 3136 7346 3188
rect 6733 3111 6791 3117
rect 6733 3108 6745 3111
rect 6104 3080 6745 3108
rect 6733 3077 6745 3080
rect 6779 3108 6791 3111
rect 9398 3108 9404 3120
rect 6779 3080 9404 3108
rect 6779 3077 6791 3080
rect 6733 3071 6791 3077
rect 9398 3068 9404 3080
rect 9456 3068 9462 3120
rect 5031 3012 5948 3040
rect 6012 3040 6040 3068
rect 6365 3043 6423 3049
rect 6365 3040 6377 3043
rect 6012 3012 6377 3040
rect 5031 3009 5043 3012
rect 4985 3003 5043 3009
rect 6365 3009 6377 3012
rect 6411 3009 6423 3043
rect 6365 3003 6423 3009
rect 2958 2932 2964 2984
rect 3016 2972 3022 2984
rect 3881 2975 3939 2981
rect 3881 2972 3893 2975
rect 3016 2944 3893 2972
rect 3016 2932 3022 2944
rect 3881 2941 3893 2944
rect 3927 2941 3939 2975
rect 3881 2935 3939 2941
rect 3896 2904 3924 2935
rect 3970 2932 3976 2984
rect 4028 2972 4034 2984
rect 4341 2975 4399 2981
rect 4341 2972 4353 2975
rect 4028 2944 4353 2972
rect 4028 2932 4034 2944
rect 4341 2941 4353 2944
rect 4387 2972 4399 2975
rect 5077 2975 5135 2981
rect 5077 2972 5089 2975
rect 4387 2944 5089 2972
rect 4387 2941 4399 2944
rect 4341 2935 4399 2941
rect 5077 2941 5089 2944
rect 5123 2941 5135 2975
rect 5077 2935 5135 2941
rect 5169 2975 5227 2981
rect 5169 2941 5181 2975
rect 5215 2972 5227 2975
rect 5629 2975 5687 2981
rect 5629 2972 5641 2975
rect 5215 2944 5641 2972
rect 5215 2941 5227 2944
rect 5169 2935 5227 2941
rect 5629 2941 5641 2944
rect 5675 2972 5687 2975
rect 5718 2972 5724 2984
rect 5675 2944 5724 2972
rect 5675 2941 5687 2944
rect 5629 2935 5687 2941
rect 4430 2904 4436 2916
rect 3896 2876 4436 2904
rect 4430 2864 4436 2876
rect 4488 2904 4494 2916
rect 5184 2904 5212 2935
rect 5718 2932 5724 2944
rect 5776 2972 5782 2984
rect 5776 2944 6224 2972
rect 5776 2932 5782 2944
rect 4488 2876 5212 2904
rect 4488 2864 4494 2876
rect 4798 2796 4804 2848
rect 4856 2796 4862 2848
rect 5902 2796 5908 2848
rect 5960 2836 5966 2848
rect 5997 2839 6055 2845
rect 5997 2836 6009 2839
rect 5960 2808 6009 2836
rect 5960 2796 5966 2808
rect 5997 2805 6009 2808
rect 6043 2805 6055 2839
rect 6196 2836 6224 2944
rect 6733 2839 6791 2845
rect 6733 2836 6745 2839
rect 6196 2808 6745 2836
rect 5997 2799 6055 2805
rect 6733 2805 6745 2808
rect 6779 2805 6791 2839
rect 6733 2799 6791 2805
rect 6914 2796 6920 2848
rect 6972 2796 6978 2848
rect 1104 2746 10488 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 10488 2746
rect 1104 2672 10488 2694
rect 5718 2592 5724 2644
rect 5776 2632 5782 2644
rect 5997 2635 6055 2641
rect 5997 2632 6009 2635
rect 5776 2604 6009 2632
rect 5776 2592 5782 2604
rect 5997 2601 6009 2604
rect 6043 2601 6055 2635
rect 5997 2595 6055 2601
rect 5629 2567 5687 2573
rect 5629 2533 5641 2567
rect 5675 2564 5687 2567
rect 5902 2564 5908 2576
rect 5675 2536 5908 2564
rect 5675 2533 5687 2536
rect 5629 2527 5687 2533
rect 5902 2524 5908 2536
rect 5960 2524 5966 2576
rect 2958 2456 2964 2508
rect 3016 2456 3022 2508
rect 3970 2456 3976 2508
rect 4028 2496 4034 2508
rect 4065 2499 4123 2505
rect 4065 2496 4077 2499
rect 4028 2468 4077 2496
rect 4028 2456 4034 2468
rect 4065 2465 4077 2468
rect 4111 2465 4123 2499
rect 4065 2459 4123 2465
rect 2682 2388 2688 2440
rect 2740 2388 2746 2440
rect 3234 2388 3240 2440
rect 3292 2428 3298 2440
rect 3789 2431 3847 2437
rect 3789 2428 3801 2431
rect 3292 2400 3801 2428
rect 3292 2388 3298 2400
rect 3789 2397 3801 2400
rect 3835 2397 3847 2431
rect 3789 2391 3847 2397
rect 4080 2360 4108 2459
rect 9398 2456 9404 2508
rect 9456 2456 9462 2508
rect 4798 2388 4804 2440
rect 4856 2428 4862 2440
rect 4893 2431 4951 2437
rect 4893 2428 4905 2431
rect 4856 2400 4905 2428
rect 4856 2388 4862 2400
rect 4893 2397 4905 2400
rect 4939 2397 4951 2431
rect 4893 2391 4951 2397
rect 5261 2431 5319 2437
rect 5261 2397 5273 2431
rect 5307 2428 5319 2431
rect 5350 2428 5356 2440
rect 5307 2400 5356 2428
rect 5307 2397 5319 2400
rect 5261 2391 5319 2397
rect 5350 2388 5356 2400
rect 5408 2388 5414 2440
rect 6086 2388 6092 2440
rect 6144 2428 6150 2440
rect 6549 2431 6607 2437
rect 6549 2428 6561 2431
rect 6144 2400 6561 2428
rect 6144 2388 6150 2400
rect 6549 2397 6561 2400
rect 6595 2397 6607 2431
rect 6549 2391 6607 2397
rect 6914 2388 6920 2440
rect 6972 2428 6978 2440
rect 7193 2431 7251 2437
rect 7193 2428 7205 2431
rect 6972 2400 7205 2428
rect 6972 2388 6978 2400
rect 7193 2397 7205 2400
rect 7239 2397 7251 2431
rect 7193 2391 7251 2397
rect 7282 2388 7288 2440
rect 7340 2428 7346 2440
rect 7837 2431 7895 2437
rect 7837 2428 7849 2431
rect 7340 2400 7849 2428
rect 7340 2388 7346 2400
rect 7837 2397 7849 2400
rect 7883 2397 7895 2431
rect 7837 2391 7895 2397
rect 8481 2431 8539 2437
rect 8481 2397 8493 2431
rect 8527 2397 8539 2431
rect 8481 2391 8539 2397
rect 5994 2360 6000 2372
rect 4080 2332 6000 2360
rect 5994 2320 6000 2332
rect 6052 2320 6058 2372
rect 8496 2360 8524 2391
rect 9122 2388 9128 2440
rect 9180 2388 9186 2440
rect 6196 2332 8524 2360
rect 5074 2252 5080 2304
rect 5132 2252 5138 2304
rect 5445 2295 5503 2301
rect 5445 2261 5457 2295
rect 5491 2292 5503 2295
rect 5810 2292 5816 2304
rect 5491 2264 5816 2292
rect 5491 2261 5503 2264
rect 5445 2255 5503 2261
rect 5810 2252 5816 2264
rect 5868 2252 5874 2304
rect 6196 2301 6224 2332
rect 6181 2295 6239 2301
rect 6181 2261 6193 2295
rect 6227 2261 6239 2295
rect 6181 2255 6239 2261
rect 6454 2252 6460 2304
rect 6512 2292 6518 2304
rect 6733 2295 6791 2301
rect 6733 2292 6745 2295
rect 6512 2264 6745 2292
rect 6512 2252 6518 2264
rect 6733 2261 6745 2264
rect 6779 2261 6791 2295
rect 6733 2255 6791 2261
rect 7098 2252 7104 2304
rect 7156 2292 7162 2304
rect 7377 2295 7435 2301
rect 7377 2292 7389 2295
rect 7156 2264 7389 2292
rect 7156 2252 7162 2264
rect 7377 2261 7389 2264
rect 7423 2261 7435 2295
rect 7377 2255 7435 2261
rect 7742 2252 7748 2304
rect 7800 2292 7806 2304
rect 8021 2295 8079 2301
rect 8021 2292 8033 2295
rect 7800 2264 8033 2292
rect 7800 2252 7806 2264
rect 8021 2261 8033 2264
rect 8067 2261 8079 2295
rect 8021 2255 8079 2261
rect 8386 2252 8392 2304
rect 8444 2292 8450 2304
rect 8665 2295 8723 2301
rect 8665 2292 8677 2295
rect 8444 2264 8677 2292
rect 8444 2252 8450 2264
rect 8665 2261 8677 2264
rect 8711 2261 8723 2295
rect 8665 2255 8723 2261
rect 1104 2202 10488 2224
rect 1104 2150 4874 2202
rect 4926 2150 4938 2202
rect 4990 2150 5002 2202
rect 5054 2150 5066 2202
rect 5118 2150 5130 2202
rect 5182 2150 10488 2202
rect 1104 2128 10488 2150
<< via1 >>
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 5816 11296 5868 11348
rect 5632 11271 5684 11280
rect 5632 11237 5641 11271
rect 5641 11237 5675 11271
rect 5675 11237 5684 11271
rect 5632 11228 5684 11237
rect 4712 11135 4764 11144
rect 4712 11101 4721 11135
rect 4721 11101 4755 11135
rect 4755 11101 4764 11135
rect 4712 11092 4764 11101
rect 5816 11160 5868 11212
rect 4252 11024 4304 11076
rect 5540 11092 5592 11144
rect 6092 11092 6144 11144
rect 4896 11067 4948 11076
rect 4896 11033 4905 11067
rect 4905 11033 4939 11067
rect 4939 11033 4948 11067
rect 4896 11024 4948 11033
rect 5448 11067 5500 11076
rect 5448 11033 5457 11067
rect 5457 11033 5491 11067
rect 5491 11033 5500 11067
rect 5448 11024 5500 11033
rect 6000 11024 6052 11076
rect 4160 10956 4212 11008
rect 5908 10956 5960 11008
rect 4874 10854 4926 10906
rect 4938 10854 4990 10906
rect 5002 10854 5054 10906
rect 5066 10854 5118 10906
rect 5130 10854 5182 10906
rect 2780 10752 2832 10804
rect 3700 10616 3752 10668
rect 3976 10752 4028 10804
rect 4804 10548 4856 10600
rect 6000 10752 6052 10804
rect 5816 10684 5868 10736
rect 7196 10684 7248 10736
rect 4160 10480 4212 10532
rect 4068 10455 4120 10464
rect 4068 10421 4077 10455
rect 4077 10421 4111 10455
rect 4111 10421 4120 10455
rect 4068 10412 4120 10421
rect 4252 10412 4304 10464
rect 6092 10455 6144 10464
rect 6092 10421 6101 10455
rect 6101 10421 6135 10455
rect 6135 10421 6144 10455
rect 6092 10412 6144 10421
rect 6276 10548 6328 10600
rect 7380 10548 7432 10600
rect 6736 10412 6788 10464
rect 8116 10455 8168 10464
rect 8116 10421 8125 10455
rect 8125 10421 8159 10455
rect 8159 10421 8168 10455
rect 8116 10412 8168 10421
rect 8208 10455 8260 10464
rect 8208 10421 8217 10455
rect 8217 10421 8251 10455
rect 8251 10421 8260 10455
rect 8208 10412 8260 10421
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 4804 10251 4856 10260
rect 4804 10217 4813 10251
rect 4813 10217 4847 10251
rect 4847 10217 4856 10251
rect 4804 10208 4856 10217
rect 6092 10208 6144 10260
rect 6276 10208 6328 10260
rect 2780 10072 2832 10124
rect 5908 10072 5960 10124
rect 7656 10072 7708 10124
rect 3240 10004 3292 10056
rect 3700 10004 3752 10056
rect 4436 10047 4488 10056
rect 4436 10013 4445 10047
rect 4445 10013 4479 10047
rect 4479 10013 4488 10047
rect 4436 10004 4488 10013
rect 4896 10047 4948 10056
rect 4896 10013 4938 10047
rect 4938 10013 4948 10047
rect 4896 10004 4948 10013
rect 1768 9936 1820 9988
rect 5632 10004 5684 10056
rect 5908 9979 5960 9988
rect 5908 9945 5917 9979
rect 5917 9945 5951 9979
rect 5951 9945 5960 9979
rect 5908 9936 5960 9945
rect 6460 9979 6512 9988
rect 6460 9945 6469 9979
rect 6469 9945 6503 9979
rect 6503 9945 6512 9979
rect 6460 9936 6512 9945
rect 6736 9936 6788 9988
rect 8116 9936 8168 9988
rect 9036 9936 9088 9988
rect 3792 9911 3844 9920
rect 3792 9877 3801 9911
rect 3801 9877 3835 9911
rect 3835 9877 3844 9911
rect 3792 9868 3844 9877
rect 5724 9868 5776 9920
rect 6644 9868 6696 9920
rect 7472 9868 7524 9920
rect 8024 9868 8076 9920
rect 8300 9868 8352 9920
rect 4874 9766 4926 9818
rect 4938 9766 4990 9818
rect 5002 9766 5054 9818
rect 5066 9766 5118 9818
rect 5130 9766 5182 9818
rect 3792 9664 3844 9716
rect 4436 9664 4488 9716
rect 5080 9664 5132 9716
rect 1768 9503 1820 9512
rect 1768 9469 1777 9503
rect 1777 9469 1811 9503
rect 1811 9469 1820 9503
rect 1768 9460 1820 9469
rect 2320 9460 2372 9512
rect 3516 9528 3568 9580
rect 5264 9634 5316 9686
rect 5540 9664 5592 9716
rect 5816 9664 5868 9716
rect 6460 9664 6512 9716
rect 6644 9664 6696 9716
rect 7380 9707 7432 9716
rect 7380 9673 7389 9707
rect 7389 9673 7423 9707
rect 7423 9673 7432 9707
rect 7380 9664 7432 9673
rect 4068 9571 4120 9580
rect 4068 9537 4077 9571
rect 4077 9537 4111 9571
rect 4111 9537 4120 9571
rect 4068 9528 4120 9537
rect 4988 9571 5040 9580
rect 4988 9537 4997 9571
rect 4997 9537 5031 9571
rect 5031 9537 5040 9571
rect 4988 9528 5040 9537
rect 5172 9571 5224 9580
rect 5172 9537 5181 9571
rect 5181 9537 5215 9571
rect 5215 9537 5224 9571
rect 5172 9528 5224 9537
rect 5356 9569 5408 9580
rect 5356 9535 5365 9569
rect 5365 9535 5399 9569
rect 5399 9535 5408 9569
rect 5356 9528 5408 9535
rect 5632 9571 5684 9580
rect 5632 9537 5641 9571
rect 5641 9537 5675 9571
rect 5675 9537 5684 9571
rect 5632 9528 5684 9537
rect 6000 9528 6052 9580
rect 6644 9528 6696 9580
rect 7564 9571 7616 9602
rect 7564 9550 7573 9571
rect 7573 9550 7607 9571
rect 7607 9550 7616 9571
rect 7656 9639 7708 9648
rect 7656 9605 7665 9639
rect 7665 9605 7699 9639
rect 7699 9605 7708 9639
rect 7656 9596 7708 9605
rect 8024 9664 8076 9716
rect 8116 9596 8168 9648
rect 2688 9435 2740 9444
rect 2688 9401 2697 9435
rect 2697 9401 2731 9435
rect 2731 9401 2740 9435
rect 2688 9392 2740 9401
rect 4712 9460 4764 9512
rect 2872 9367 2924 9376
rect 2872 9333 2881 9367
rect 2881 9333 2915 9367
rect 2915 9333 2924 9367
rect 2872 9324 2924 9333
rect 3240 9324 3292 9376
rect 3424 9324 3476 9376
rect 5172 9392 5224 9444
rect 6000 9435 6052 9444
rect 6000 9401 6009 9435
rect 6009 9401 6043 9435
rect 6043 9401 6052 9435
rect 6000 9392 6052 9401
rect 7472 9460 7524 9512
rect 8208 9528 8260 9580
rect 8392 9571 8444 9580
rect 8392 9537 8401 9571
rect 8401 9537 8435 9571
rect 8435 9537 8444 9571
rect 8392 9528 8444 9537
rect 9128 9528 9180 9580
rect 4068 9324 4120 9376
rect 4620 9324 4672 9376
rect 5264 9324 5316 9376
rect 6644 9324 6696 9376
rect 8760 9392 8812 9444
rect 8852 9324 8904 9376
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 2872 9163 2924 9172
rect 2872 9129 2893 9163
rect 2893 9129 2924 9163
rect 2872 9120 2924 9129
rect 4252 9120 4304 9172
rect 4988 9120 5040 9172
rect 5448 9120 5500 9172
rect 6092 9120 6144 9172
rect 7012 9120 7064 9172
rect 8392 9120 8444 9172
rect 4344 9052 4396 9104
rect 5632 9052 5684 9104
rect 5724 9095 5776 9104
rect 5724 9061 5733 9095
rect 5733 9061 5767 9095
rect 5767 9061 5776 9095
rect 5724 9052 5776 9061
rect 5816 9052 5868 9104
rect 6368 9052 6420 9104
rect 7564 9052 7616 9104
rect 8484 9052 8536 9104
rect 2780 8984 2832 9036
rect 4528 8984 4580 9036
rect 3148 8848 3200 8900
rect 1400 8823 1452 8832
rect 1400 8789 1409 8823
rect 1409 8789 1443 8823
rect 1443 8789 1452 8823
rect 1400 8780 1452 8789
rect 3424 8823 3476 8832
rect 3424 8789 3433 8823
rect 3433 8789 3467 8823
rect 3467 8789 3476 8823
rect 3424 8780 3476 8789
rect 3792 8823 3844 8832
rect 3792 8789 3801 8823
rect 3801 8789 3835 8823
rect 3835 8789 3844 8823
rect 3792 8780 3844 8789
rect 4436 8959 4488 8968
rect 4436 8925 4445 8959
rect 4445 8925 4479 8959
rect 4479 8925 4488 8959
rect 4436 8916 4488 8925
rect 5080 8959 5132 8968
rect 5080 8925 5089 8959
rect 5089 8925 5123 8959
rect 5123 8925 5132 8959
rect 5080 8916 5132 8925
rect 4160 8780 4212 8832
rect 4252 8823 4304 8832
rect 4252 8789 4261 8823
rect 4261 8789 4295 8823
rect 4295 8789 4304 8823
rect 4252 8780 4304 8789
rect 4344 8823 4396 8832
rect 4344 8789 4353 8823
rect 4353 8789 4387 8823
rect 4387 8789 4396 8823
rect 4344 8780 4396 8789
rect 4436 8780 4488 8832
rect 4620 8780 4672 8832
rect 6092 8959 6144 8968
rect 6092 8925 6101 8959
rect 6101 8925 6135 8959
rect 6135 8925 6144 8959
rect 6092 8916 6144 8925
rect 8668 8984 8720 9036
rect 5816 8780 5868 8832
rect 7380 8916 7432 8968
rect 8300 8916 8352 8968
rect 8760 8916 8812 8968
rect 6460 8780 6512 8832
rect 6920 8780 6972 8832
rect 8024 8780 8076 8832
rect 8576 8823 8628 8832
rect 8576 8789 8585 8823
rect 8585 8789 8619 8823
rect 8619 8789 8628 8823
rect 8576 8780 8628 8789
rect 4874 8678 4926 8730
rect 4938 8678 4990 8730
rect 5002 8678 5054 8730
rect 5066 8678 5118 8730
rect 5130 8678 5182 8730
rect 1400 8576 1452 8628
rect 2688 8619 2740 8628
rect 2688 8585 2697 8619
rect 2697 8585 2731 8619
rect 2731 8585 2740 8619
rect 2688 8576 2740 8585
rect 2872 8508 2924 8560
rect 3424 8576 3476 8628
rect 3884 8576 3936 8628
rect 4344 8576 4396 8628
rect 3516 8508 3568 8560
rect 3792 8508 3844 8560
rect 2412 8440 2464 8492
rect 4436 8440 4488 8492
rect 4712 8576 4764 8628
rect 5540 8576 5592 8628
rect 2688 8304 2740 8356
rect 4160 8372 4212 8424
rect 5632 8440 5684 8492
rect 5724 8440 5776 8492
rect 6644 8576 6696 8628
rect 8300 8576 8352 8628
rect 8576 8576 8628 8628
rect 8668 8576 8720 8628
rect 9036 8619 9088 8628
rect 9036 8585 9045 8619
rect 9045 8585 9079 8619
rect 9079 8585 9088 8619
rect 9036 8576 9088 8585
rect 6184 8440 6236 8492
rect 7196 8508 7248 8560
rect 4712 8236 4764 8288
rect 5080 8304 5132 8356
rect 6000 8372 6052 8424
rect 8484 8483 8536 8492
rect 8484 8449 8493 8483
rect 8493 8449 8527 8483
rect 8527 8449 8536 8483
rect 8484 8440 8536 8449
rect 8852 8440 8904 8492
rect 6920 8236 6972 8288
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 2320 8075 2372 8084
rect 2320 8041 2329 8075
rect 2329 8041 2363 8075
rect 2363 8041 2372 8075
rect 2320 8032 2372 8041
rect 6276 8032 6328 8084
rect 2964 8007 3016 8016
rect 2964 7973 2973 8007
rect 2973 7973 3007 8007
rect 3007 7973 3016 8007
rect 2964 7964 3016 7973
rect 5080 7964 5132 8016
rect 5540 7964 5592 8016
rect 1676 7939 1728 7948
rect 1676 7905 1685 7939
rect 1685 7905 1719 7939
rect 1719 7905 1728 7939
rect 1676 7896 1728 7905
rect 8392 8007 8444 8016
rect 8392 7973 8401 8007
rect 8401 7973 8435 8007
rect 8435 7973 8444 8007
rect 8392 7964 8444 7973
rect 1400 7871 1452 7880
rect 1400 7837 1409 7871
rect 1409 7837 1443 7871
rect 1443 7837 1452 7871
rect 1400 7828 1452 7837
rect 2044 7871 2096 7880
rect 2044 7837 2053 7871
rect 2053 7837 2087 7871
rect 2087 7837 2096 7871
rect 2044 7828 2096 7837
rect 2688 7871 2740 7880
rect 2688 7837 2697 7871
rect 2697 7837 2731 7871
rect 2731 7837 2740 7871
rect 2688 7828 2740 7837
rect 2872 7803 2924 7812
rect 2872 7769 2881 7803
rect 2881 7769 2915 7803
rect 2915 7769 2924 7803
rect 2872 7760 2924 7769
rect 3240 7828 3292 7880
rect 3884 7828 3936 7880
rect 8484 7896 8536 7948
rect 4620 7871 4672 7880
rect 4620 7837 4629 7871
rect 4629 7837 4663 7871
rect 4663 7837 4672 7871
rect 4620 7828 4672 7837
rect 4804 7871 4856 7880
rect 4804 7837 4813 7871
rect 4813 7837 4847 7871
rect 4847 7837 4856 7871
rect 4804 7828 4856 7837
rect 1584 7735 1636 7744
rect 1584 7701 1593 7735
rect 1593 7701 1627 7735
rect 1627 7701 1636 7735
rect 1584 7692 1636 7701
rect 3424 7692 3476 7744
rect 4436 7760 4488 7812
rect 6920 7803 6972 7812
rect 6920 7769 6929 7803
rect 6929 7769 6963 7803
rect 6963 7769 6972 7803
rect 6920 7760 6972 7769
rect 7196 7760 7248 7812
rect 3608 7692 3660 7744
rect 3700 7692 3752 7744
rect 4344 7692 4396 7744
rect 6092 7735 6144 7744
rect 6092 7701 6101 7735
rect 6101 7701 6135 7735
rect 6135 7701 6144 7735
rect 6092 7692 6144 7701
rect 6276 7692 6328 7744
rect 6736 7692 6788 7744
rect 7748 7692 7800 7744
rect 8944 7735 8996 7744
rect 8944 7701 8953 7735
rect 8953 7701 8987 7735
rect 8987 7701 8996 7735
rect 8944 7692 8996 7701
rect 4874 7590 4926 7642
rect 4938 7590 4990 7642
rect 5002 7590 5054 7642
rect 5066 7590 5118 7642
rect 5130 7590 5182 7642
rect 1124 7488 1176 7540
rect 2044 7488 2096 7540
rect 2780 7488 2832 7540
rect 6092 7488 6144 7540
rect 6184 7531 6236 7540
rect 6184 7497 6193 7531
rect 6193 7497 6227 7531
rect 6227 7497 6236 7531
rect 6184 7488 6236 7497
rect 6920 7488 6972 7540
rect 8484 7488 8536 7540
rect 4344 7463 4396 7472
rect 4344 7429 4353 7463
rect 4353 7429 4387 7463
rect 4387 7429 4396 7463
rect 4344 7420 4396 7429
rect 4712 7463 4764 7472
rect 4712 7429 4721 7463
rect 4721 7429 4755 7463
rect 4755 7429 4764 7463
rect 4712 7420 4764 7429
rect 8944 7420 8996 7472
rect 2412 7327 2464 7336
rect 2412 7293 2421 7327
rect 2421 7293 2455 7327
rect 2455 7293 2464 7327
rect 2412 7284 2464 7293
rect 5724 7352 5776 7404
rect 6276 7352 6328 7404
rect 6828 7352 6880 7404
rect 2872 7284 2924 7336
rect 3608 7284 3660 7336
rect 7288 7352 7340 7404
rect 7932 7352 7984 7404
rect 6276 7216 6328 7268
rect 7012 7216 7064 7268
rect 4436 7148 4488 7200
rect 4804 7148 4856 7200
rect 6368 7148 6420 7200
rect 6828 7148 6880 7200
rect 7472 7148 7524 7200
rect 7564 7191 7616 7200
rect 7564 7157 7573 7191
rect 7573 7157 7607 7191
rect 7607 7157 7616 7191
rect 7564 7148 7616 7157
rect 7932 7148 7984 7200
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 1676 6987 1728 6996
rect 1676 6953 1706 6987
rect 1706 6953 1728 6987
rect 1676 6944 1728 6953
rect 2780 6944 2832 6996
rect 3792 6944 3844 6996
rect 4436 6944 4488 6996
rect 5356 6944 5408 6996
rect 5632 6987 5684 6996
rect 5632 6953 5641 6987
rect 5641 6953 5675 6987
rect 5675 6953 5684 6987
rect 5632 6944 5684 6953
rect 4620 6808 4672 6860
rect 5540 6808 5592 6860
rect 3148 6740 3200 6792
rect 3700 6740 3752 6792
rect 4160 6672 4212 6724
rect 5448 6672 5500 6724
rect 6000 6783 6052 6792
rect 6000 6749 6009 6783
rect 6009 6749 6043 6783
rect 6043 6749 6052 6783
rect 6000 6740 6052 6749
rect 6552 6987 6604 6996
rect 6552 6953 6561 6987
rect 6561 6953 6595 6987
rect 6595 6953 6604 6987
rect 6552 6944 6604 6953
rect 6920 6944 6972 6996
rect 7288 6944 7340 6996
rect 6828 6876 6880 6928
rect 8024 6919 8076 6928
rect 8024 6885 8033 6919
rect 8033 6885 8067 6919
rect 8067 6885 8076 6919
rect 8024 6876 8076 6885
rect 8300 6919 8352 6928
rect 8300 6885 8309 6919
rect 8309 6885 8343 6919
rect 8343 6885 8352 6919
rect 8300 6876 8352 6885
rect 6460 6808 6512 6860
rect 7840 6808 7892 6860
rect 8760 6808 8812 6860
rect 2412 6604 2464 6656
rect 3332 6647 3384 6656
rect 3332 6613 3341 6647
rect 3341 6613 3375 6647
rect 3375 6613 3384 6647
rect 3332 6604 3384 6613
rect 6828 6740 6880 6792
rect 7288 6740 7340 6792
rect 9128 6783 9180 6792
rect 9128 6749 9137 6783
rect 9137 6749 9171 6783
rect 9171 6749 9180 6783
rect 9128 6740 9180 6749
rect 6736 6604 6788 6656
rect 7196 6647 7248 6656
rect 7196 6613 7221 6647
rect 7221 6613 7248 6647
rect 7196 6604 7248 6613
rect 7380 6647 7432 6656
rect 7380 6613 7389 6647
rect 7389 6613 7423 6647
rect 7423 6613 7432 6647
rect 7380 6604 7432 6613
rect 9036 6672 9088 6724
rect 7840 6647 7892 6656
rect 7840 6613 7849 6647
rect 7849 6613 7883 6647
rect 7883 6613 7892 6647
rect 7840 6604 7892 6613
rect 8116 6647 8168 6656
rect 8116 6613 8125 6647
rect 8125 6613 8159 6647
rect 8159 6613 8168 6647
rect 8116 6604 8168 6613
rect 4874 6502 4926 6554
rect 4938 6502 4990 6554
rect 5002 6502 5054 6554
rect 5066 6502 5118 6554
rect 5130 6502 5182 6554
rect 2780 6400 2832 6452
rect 2964 6400 3016 6452
rect 1584 6307 1636 6316
rect 1584 6273 1593 6307
rect 1593 6273 1627 6307
rect 1627 6273 1636 6307
rect 1584 6264 1636 6273
rect 2320 6332 2372 6384
rect 4712 6400 4764 6452
rect 4160 6332 4212 6384
rect 4436 6332 4488 6384
rect 6276 6400 6328 6452
rect 6552 6400 6604 6452
rect 6644 6400 6696 6452
rect 1768 6239 1820 6248
rect 1768 6205 1777 6239
rect 1777 6205 1811 6239
rect 1811 6205 1820 6239
rect 1768 6196 1820 6205
rect 1860 6128 1912 6180
rect 2044 6103 2096 6112
rect 2044 6069 2053 6103
rect 2053 6069 2087 6103
rect 2087 6069 2096 6103
rect 2044 6060 2096 6069
rect 3148 6196 3200 6248
rect 3792 6196 3844 6248
rect 4804 6128 4856 6180
rect 3884 6060 3936 6112
rect 5908 6332 5960 6384
rect 6736 6332 6788 6384
rect 5356 6264 5408 6316
rect 6184 6264 6236 6316
rect 7196 6264 7248 6316
rect 7288 6307 7340 6316
rect 7288 6273 7297 6307
rect 7297 6273 7331 6307
rect 7331 6273 7340 6307
rect 7288 6264 7340 6273
rect 8116 6400 8168 6452
rect 6920 6196 6972 6248
rect 6828 6128 6880 6180
rect 7104 6171 7156 6180
rect 7104 6137 7113 6171
rect 7113 6137 7147 6171
rect 7147 6137 7156 6171
rect 7104 6128 7156 6137
rect 5264 6103 5316 6112
rect 5264 6069 5273 6103
rect 5273 6069 5307 6103
rect 5307 6069 5316 6103
rect 5264 6060 5316 6069
rect 6736 6060 6788 6112
rect 7380 6128 7432 6180
rect 7288 6060 7340 6112
rect 8392 6060 8444 6112
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 1860 5856 1912 5908
rect 2044 5856 2096 5908
rect 2780 5788 2832 5840
rect 3424 5899 3476 5908
rect 3424 5865 3433 5899
rect 3433 5865 3467 5899
rect 3467 5865 3476 5899
rect 3424 5856 3476 5865
rect 3792 5856 3844 5908
rect 3976 5899 4028 5908
rect 3976 5865 3985 5899
rect 3985 5865 4019 5899
rect 4019 5865 4028 5899
rect 3976 5856 4028 5865
rect 4620 5856 4672 5908
rect 5264 5856 5316 5908
rect 5448 5856 5500 5908
rect 7196 5856 7248 5908
rect 8392 5856 8444 5908
rect 5172 5720 5224 5772
rect 8484 5720 8536 5772
rect 2320 5584 2372 5636
rect 4620 5584 4672 5636
rect 4344 5516 4396 5568
rect 4804 5516 4856 5568
rect 6092 5584 6144 5636
rect 6644 5627 6696 5636
rect 6644 5593 6653 5627
rect 6653 5593 6687 5627
rect 6687 5593 6696 5627
rect 6644 5584 6696 5593
rect 7748 5584 7800 5636
rect 10508 5584 10560 5636
rect 6276 5516 6328 5568
rect 7104 5516 7156 5568
rect 7472 5516 7524 5568
rect 4874 5414 4926 5466
rect 4938 5414 4990 5466
rect 5002 5414 5054 5466
rect 5066 5414 5118 5466
rect 5130 5414 5182 5466
rect 1768 5312 1820 5364
rect 1124 5244 1176 5296
rect 1400 5219 1452 5228
rect 1400 5185 1409 5219
rect 1409 5185 1443 5219
rect 1443 5185 1452 5219
rect 1400 5176 1452 5185
rect 2780 5312 2832 5364
rect 6184 5355 6236 5364
rect 6184 5321 6193 5355
rect 6193 5321 6227 5355
rect 6227 5321 6236 5355
rect 6184 5312 6236 5321
rect 6276 5312 6328 5364
rect 6644 5312 6696 5364
rect 3332 5108 3384 5160
rect 7564 5312 7616 5364
rect 7748 5312 7800 5364
rect 8484 5312 8536 5364
rect 4068 5108 4120 5160
rect 4712 5151 4764 5160
rect 4712 5117 4721 5151
rect 4721 5117 4755 5151
rect 4755 5117 4764 5151
rect 4712 5108 4764 5117
rect 6092 5108 6144 5160
rect 4344 5083 4396 5092
rect 4344 5049 4353 5083
rect 4353 5049 4387 5083
rect 4387 5049 4396 5083
rect 4344 5040 4396 5049
rect 2320 5015 2372 5024
rect 2320 4981 2329 5015
rect 2329 4981 2363 5015
rect 2363 4981 2372 5015
rect 2320 4972 2372 4981
rect 6920 5108 6972 5160
rect 6368 5040 6420 5092
rect 6644 5083 6696 5092
rect 6644 5049 6653 5083
rect 6653 5049 6687 5083
rect 6687 5049 6696 5083
rect 6644 5040 6696 5049
rect 6736 5083 6788 5092
rect 6736 5049 6745 5083
rect 6745 5049 6779 5083
rect 6779 5049 6788 5083
rect 6736 5040 6788 5049
rect 6828 5040 6880 5092
rect 8208 5108 8260 5160
rect 8576 5151 8628 5160
rect 8576 5117 8585 5151
rect 8585 5117 8619 5151
rect 8619 5117 8628 5151
rect 8576 5108 8628 5117
rect 7564 5040 7616 5092
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 2780 4768 2832 4820
rect 3148 4811 3200 4820
rect 3148 4777 3157 4811
rect 3157 4777 3191 4811
rect 3191 4777 3200 4811
rect 3148 4768 3200 4777
rect 3332 4768 3384 4820
rect 3976 4811 4028 4820
rect 3976 4777 3985 4811
rect 3985 4777 4019 4811
rect 4019 4777 4028 4811
rect 3976 4768 4028 4777
rect 4712 4768 4764 4820
rect 6828 4811 6880 4820
rect 6828 4777 6837 4811
rect 6837 4777 6871 4811
rect 6871 4777 6880 4811
rect 6828 4768 6880 4777
rect 6920 4768 6972 4820
rect 7932 4768 7984 4820
rect 4804 4700 4856 4752
rect 6736 4743 6788 4752
rect 4620 4632 4672 4684
rect 6736 4709 6745 4743
rect 6745 4709 6779 4743
rect 6779 4709 6788 4743
rect 6736 4700 6788 4709
rect 6184 4632 6236 4684
rect 7104 4632 7156 4684
rect 1676 4539 1728 4548
rect 1676 4505 1685 4539
rect 1685 4505 1719 4539
rect 1719 4505 1728 4539
rect 1676 4496 1728 4505
rect 2320 4496 2372 4548
rect 5540 4564 5592 4616
rect 6644 4607 6696 4616
rect 6644 4573 6653 4607
rect 6653 4573 6687 4607
rect 6687 4573 6696 4607
rect 6644 4564 6696 4573
rect 7840 4607 7892 4616
rect 7840 4573 7849 4607
rect 7849 4573 7883 4607
rect 7883 4573 7892 4607
rect 7840 4564 7892 4573
rect 4436 4428 4488 4480
rect 5908 4471 5960 4480
rect 5908 4437 5917 4471
rect 5917 4437 5951 4471
rect 5951 4437 5960 4471
rect 5908 4428 5960 4437
rect 7104 4471 7156 4480
rect 7104 4437 7113 4471
rect 7113 4437 7147 4471
rect 7147 4437 7156 4471
rect 7104 4428 7156 4437
rect 4874 4326 4926 4378
rect 4938 4326 4990 4378
rect 5002 4326 5054 4378
rect 5066 4326 5118 4378
rect 5130 4326 5182 4378
rect 1676 4224 1728 4276
rect 4068 4224 4120 4276
rect 4804 4224 4856 4276
rect 5908 4224 5960 4276
rect 7104 4224 7156 4276
rect 4436 4199 4488 4208
rect 4436 4165 4445 4199
rect 4445 4165 4479 4199
rect 4479 4165 4488 4199
rect 4436 4156 4488 4165
rect 2044 4131 2096 4140
rect 2044 4097 2053 4131
rect 2053 4097 2087 4131
rect 2087 4097 2096 4131
rect 2044 4088 2096 4097
rect 5356 4020 5408 4072
rect 1492 3995 1544 4004
rect 1492 3961 1501 3995
rect 1501 3961 1535 3995
rect 1535 3961 1544 3995
rect 1492 3952 1544 3961
rect 5540 3952 5592 4004
rect 6092 4020 6144 4072
rect 7288 4020 7340 4072
rect 8576 4020 8628 4072
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 2044 3680 2096 3732
rect 5724 3544 5776 3596
rect 940 3476 992 3528
rect 3976 3519 4028 3528
rect 3976 3485 3985 3519
rect 3985 3485 4019 3519
rect 4019 3485 4028 3519
rect 3976 3476 4028 3485
rect 4620 3519 4672 3528
rect 4620 3485 4629 3519
rect 4629 3485 4663 3519
rect 4663 3485 4672 3519
rect 4620 3476 4672 3485
rect 5908 3476 5960 3528
rect 6000 3408 6052 3460
rect 3884 3340 3936 3392
rect 4804 3383 4856 3392
rect 4804 3349 4813 3383
rect 4813 3349 4847 3383
rect 4847 3349 4856 3383
rect 4804 3340 4856 3349
rect 5356 3383 5408 3392
rect 5356 3349 5365 3383
rect 5365 3349 5399 3383
rect 5399 3349 5408 3383
rect 5356 3340 5408 3349
rect 6092 3383 6144 3392
rect 6092 3349 6101 3383
rect 6101 3349 6135 3383
rect 6135 3349 6144 3383
rect 6092 3340 6144 3349
rect 4874 3238 4926 3290
rect 4938 3238 4990 3290
rect 5002 3238 5054 3290
rect 5066 3238 5118 3290
rect 5130 3238 5182 3290
rect 3976 3136 4028 3188
rect 4620 3136 4672 3188
rect 5908 3136 5960 3188
rect 4436 3043 4488 3052
rect 4436 3009 4445 3043
rect 4445 3009 4479 3043
rect 4479 3009 4488 3043
rect 4436 3000 4488 3009
rect 6000 3111 6052 3120
rect 6000 3077 6009 3111
rect 6009 3077 6043 3111
rect 6043 3077 6052 3111
rect 6000 3068 6052 3077
rect 7288 3136 7340 3188
rect 9404 3068 9456 3120
rect 2964 2932 3016 2984
rect 3976 2975 4028 2984
rect 3976 2941 3985 2975
rect 3985 2941 4019 2975
rect 4019 2941 4028 2975
rect 3976 2932 4028 2941
rect 4436 2864 4488 2916
rect 5724 2932 5776 2984
rect 4804 2839 4856 2848
rect 4804 2805 4813 2839
rect 4813 2805 4847 2839
rect 4847 2805 4856 2839
rect 4804 2796 4856 2805
rect 5908 2796 5960 2848
rect 6920 2839 6972 2848
rect 6920 2805 6929 2839
rect 6929 2805 6963 2839
rect 6963 2805 6972 2839
rect 6920 2796 6972 2805
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 5724 2592 5776 2644
rect 5908 2524 5960 2576
rect 2964 2499 3016 2508
rect 2964 2465 2973 2499
rect 2973 2465 3007 2499
rect 3007 2465 3016 2499
rect 2964 2456 3016 2465
rect 3976 2456 4028 2508
rect 2688 2431 2740 2440
rect 2688 2397 2697 2431
rect 2697 2397 2731 2431
rect 2731 2397 2740 2431
rect 2688 2388 2740 2397
rect 3240 2388 3292 2440
rect 9404 2499 9456 2508
rect 9404 2465 9413 2499
rect 9413 2465 9447 2499
rect 9447 2465 9456 2499
rect 9404 2456 9456 2465
rect 4804 2388 4856 2440
rect 5356 2388 5408 2440
rect 6092 2388 6144 2440
rect 6920 2388 6972 2440
rect 7288 2388 7340 2440
rect 6000 2363 6052 2372
rect 6000 2329 6009 2363
rect 6009 2329 6043 2363
rect 6043 2329 6052 2363
rect 6000 2320 6052 2329
rect 9128 2431 9180 2440
rect 9128 2397 9137 2431
rect 9137 2397 9171 2431
rect 9171 2397 9180 2431
rect 9128 2388 9180 2397
rect 5080 2295 5132 2304
rect 5080 2261 5089 2295
rect 5089 2261 5123 2295
rect 5123 2261 5132 2295
rect 5080 2252 5132 2261
rect 5816 2252 5868 2304
rect 6460 2252 6512 2304
rect 7104 2252 7156 2304
rect 7748 2252 7800 2304
rect 8392 2252 8444 2304
rect 4874 2150 4926 2202
rect 4938 2150 4990 2202
rect 5002 2150 5054 2202
rect 5066 2150 5118 2202
rect 5130 2150 5182 2202
<< metal2 >>
rect 5814 12937 5870 13737
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 5828 11354 5856 12937
rect 5816 11348 5868 11354
rect 5816 11290 5868 11296
rect 5632 11280 5684 11286
rect 5632 11222 5684 11228
rect 4712 11144 4764 11150
rect 4712 11086 4764 11092
rect 5540 11144 5592 11150
rect 5540 11086 5592 11092
rect 4252 11076 4304 11082
rect 4252 11018 4304 11024
rect 4160 11008 4212 11014
rect 4160 10950 4212 10956
rect 2780 10804 2832 10810
rect 3976 10804 4028 10810
rect 2780 10746 2832 10752
rect 3712 10764 3976 10792
rect 2792 10130 2820 10746
rect 3712 10674 3740 10764
rect 3976 10746 4028 10752
rect 3700 10668 3752 10674
rect 3700 10610 3752 10616
rect 2780 10124 2832 10130
rect 2780 10066 2832 10072
rect 1768 9988 1820 9994
rect 1768 9930 1820 9936
rect 1780 9518 1808 9930
rect 1768 9512 1820 9518
rect 1768 9454 1820 9460
rect 2320 9512 2372 9518
rect 2320 9454 2372 9460
rect 1400 8832 1452 8838
rect 1400 8774 1452 8780
rect 1412 8634 1440 8774
rect 1400 8628 1452 8634
rect 1400 8570 1452 8576
rect 1122 8256 1178 8265
rect 1122 8191 1178 8200
rect 1136 7546 1164 8191
rect 2332 8090 2360 9454
rect 2688 9444 2740 9450
rect 2688 9386 2740 9392
rect 2700 8634 2728 9386
rect 2792 9042 2820 10066
rect 3712 10062 3740 10610
rect 4172 10538 4200 10950
rect 4160 10532 4212 10538
rect 4160 10474 4212 10480
rect 4264 10470 4292 11018
rect 4068 10464 4120 10470
rect 4068 10406 4120 10412
rect 4252 10464 4304 10470
rect 4252 10406 4304 10412
rect 4080 10146 4108 10406
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 4080 10118 4200 10146
rect 3240 10056 3292 10062
rect 3240 9998 3292 10004
rect 3700 10056 3752 10062
rect 3700 9998 3752 10004
rect 3252 9674 3280 9998
rect 3792 9920 3844 9926
rect 3792 9862 3844 9868
rect 3804 9722 3832 9862
rect 3160 9646 3280 9674
rect 3792 9716 3844 9722
rect 4172 9674 4200 10118
rect 4436 10056 4488 10062
rect 4436 9998 4488 10004
rect 4448 9722 4476 9998
rect 3792 9658 3844 9664
rect 4080 9646 4200 9674
rect 4436 9716 4488 9722
rect 4436 9658 4488 9664
rect 2872 9376 2924 9382
rect 2872 9318 2924 9324
rect 2884 9178 2912 9318
rect 2872 9172 2924 9178
rect 2872 9114 2924 9120
rect 2780 9036 2832 9042
rect 2780 8978 2832 8984
rect 2688 8628 2740 8634
rect 2688 8570 2740 8576
rect 2412 8492 2464 8498
rect 2412 8434 2464 8440
rect 2320 8084 2372 8090
rect 2320 8026 2372 8032
rect 1676 7948 1728 7954
rect 1676 7890 1728 7896
rect 1400 7880 1452 7886
rect 1400 7822 1452 7828
rect 1412 7585 1440 7822
rect 1584 7744 1636 7750
rect 1584 7686 1636 7692
rect 1398 7576 1454 7585
rect 1124 7540 1176 7546
rect 1398 7511 1454 7520
rect 1124 7482 1176 7488
rect 1596 6322 1624 7686
rect 1688 7002 1716 7890
rect 2044 7880 2096 7886
rect 2044 7822 2096 7828
rect 2056 7546 2084 7822
rect 2044 7540 2096 7546
rect 2044 7482 2096 7488
rect 2424 7342 2452 8434
rect 2688 8356 2740 8362
rect 2688 8298 2740 8304
rect 2700 7886 2728 8298
rect 2688 7880 2740 7886
rect 2688 7822 2740 7828
rect 2792 7546 2820 8978
rect 3160 8906 3188 9646
rect 4080 9586 4108 9646
rect 3516 9580 3568 9586
rect 3516 9522 3568 9528
rect 4068 9580 4120 9586
rect 4068 9522 4120 9528
rect 3240 9376 3292 9382
rect 3240 9318 3292 9324
rect 3424 9376 3476 9382
rect 3424 9318 3476 9324
rect 3148 8900 3200 8906
rect 3148 8842 3200 8848
rect 2872 8560 2924 8566
rect 2872 8502 2924 8508
rect 2884 7818 2912 8502
rect 2964 8016 3016 8022
rect 2964 7958 3016 7964
rect 2872 7812 2924 7818
rect 2872 7754 2924 7760
rect 2780 7540 2832 7546
rect 2780 7482 2832 7488
rect 2412 7336 2464 7342
rect 2412 7278 2464 7284
rect 1676 6996 1728 7002
rect 1676 6938 1728 6944
rect 2424 6662 2452 7278
rect 2792 7002 2820 7482
rect 2884 7342 2912 7754
rect 2872 7336 2924 7342
rect 2872 7278 2924 7284
rect 2780 6996 2832 7002
rect 2780 6938 2832 6944
rect 2412 6656 2464 6662
rect 2412 6598 2464 6604
rect 2792 6458 2820 6938
rect 2976 6458 3004 7958
rect 3160 6798 3188 8842
rect 3252 7886 3280 9318
rect 3436 8838 3464 9318
rect 3424 8832 3476 8838
rect 3424 8774 3476 8780
rect 3436 8634 3464 8774
rect 3424 8628 3476 8634
rect 3424 8570 3476 8576
rect 3240 7880 3292 7886
rect 3240 7822 3292 7828
rect 3436 7750 3464 8570
rect 3528 8566 3556 9522
rect 4080 9382 4108 9522
rect 4724 9518 4752 11086
rect 4896 11076 4948 11082
rect 4816 11036 4896 11064
rect 4816 10690 4844 11036
rect 4896 11018 4948 11024
rect 5448 11076 5500 11082
rect 5448 11018 5500 11024
rect 4874 10908 5182 10917
rect 4874 10906 4880 10908
rect 4936 10906 4960 10908
rect 5016 10906 5040 10908
rect 5096 10906 5120 10908
rect 5176 10906 5182 10908
rect 4936 10854 4938 10906
rect 5118 10854 5120 10906
rect 4874 10852 4880 10854
rect 4936 10852 4960 10854
rect 5016 10852 5040 10854
rect 5096 10852 5120 10854
rect 5176 10852 5182 10854
rect 4874 10843 5182 10852
rect 4816 10662 4936 10690
rect 4804 10600 4856 10606
rect 4804 10542 4856 10548
rect 4816 10266 4844 10542
rect 4804 10260 4856 10266
rect 4804 10202 4856 10208
rect 4908 10062 4936 10662
rect 4896 10056 4948 10062
rect 4802 10024 4858 10033
rect 4896 9998 4948 10004
rect 4802 9959 4858 9968
rect 4712 9512 4764 9518
rect 4712 9454 4764 9460
rect 4068 9376 4120 9382
rect 4068 9318 4120 9324
rect 4620 9376 4672 9382
rect 4620 9318 4672 9324
rect 4080 9160 4108 9318
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 4252 9172 4304 9178
rect 4080 9132 4252 9160
rect 4252 9114 4304 9120
rect 4264 8838 4292 9114
rect 4344 9104 4396 9110
rect 4344 9046 4396 9052
rect 4434 9072 4490 9081
rect 4356 8838 4384 9046
rect 4434 9007 4490 9016
rect 4528 9036 4580 9042
rect 4448 8974 4476 9007
rect 4528 8978 4580 8984
rect 4436 8968 4488 8974
rect 4436 8910 4488 8916
rect 4540 8922 4568 8978
rect 4632 8922 4660 9318
rect 4540 8894 4752 8922
rect 3792 8832 3844 8838
rect 3792 8774 3844 8780
rect 4160 8832 4212 8838
rect 4160 8774 4212 8780
rect 4252 8832 4304 8838
rect 4252 8774 4304 8780
rect 4344 8832 4396 8838
rect 4344 8774 4396 8780
rect 4436 8832 4488 8838
rect 4436 8774 4488 8780
rect 4620 8832 4672 8838
rect 4620 8774 4672 8780
rect 3804 8566 3832 8774
rect 3884 8628 3936 8634
rect 3884 8570 3936 8576
rect 3516 8560 3568 8566
rect 3516 8502 3568 8508
rect 3792 8560 3844 8566
rect 3792 8502 3844 8508
rect 3804 7834 3832 8502
rect 3896 7886 3924 8570
rect 4172 8430 4200 8774
rect 4356 8634 4384 8774
rect 4344 8628 4396 8634
rect 4344 8570 4396 8576
rect 4448 8498 4476 8774
rect 4436 8492 4488 8498
rect 4436 8434 4488 8440
rect 4160 8424 4212 8430
rect 4160 8366 4212 8372
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 4632 7886 4660 8774
rect 4724 8634 4752 8894
rect 4712 8628 4764 8634
rect 4712 8570 4764 8576
rect 4712 8288 4764 8294
rect 4712 8230 4764 8236
rect 3620 7806 3832 7834
rect 3884 7880 3936 7886
rect 3884 7822 3936 7828
rect 4620 7880 4672 7886
rect 4620 7822 4672 7828
rect 3620 7750 3648 7806
rect 3424 7744 3476 7750
rect 3424 7686 3476 7692
rect 3608 7744 3660 7750
rect 3608 7686 3660 7692
rect 3700 7744 3752 7750
rect 3700 7686 3752 7692
rect 3608 7336 3660 7342
rect 3608 7278 3660 7284
rect 3330 6896 3386 6905
rect 3330 6831 3386 6840
rect 3148 6792 3200 6798
rect 3148 6734 3200 6740
rect 3344 6662 3372 6831
rect 3332 6656 3384 6662
rect 3620 6644 3648 7278
rect 3712 6798 3740 7686
rect 3804 7002 3832 7806
rect 3792 6996 3844 7002
rect 3792 6938 3844 6944
rect 3700 6792 3752 6798
rect 3700 6734 3752 6740
rect 3620 6616 3832 6644
rect 3332 6598 3384 6604
rect 2780 6452 2832 6458
rect 2780 6394 2832 6400
rect 2964 6452 3016 6458
rect 2964 6394 3016 6400
rect 2320 6384 2372 6390
rect 2320 6326 2372 6332
rect 1584 6316 1636 6322
rect 1584 6258 1636 6264
rect 1768 6248 1820 6254
rect 1768 6190 1820 6196
rect 1398 5536 1454 5545
rect 1398 5471 1454 5480
rect 1124 5296 1176 5302
rect 1124 5238 1176 5244
rect 1136 4865 1164 5238
rect 1412 5234 1440 5471
rect 1780 5370 1808 6190
rect 1860 6180 1912 6186
rect 1860 6122 1912 6128
rect 1872 5914 1900 6122
rect 2044 6112 2096 6118
rect 2044 6054 2096 6060
rect 2056 5914 2084 6054
rect 1860 5908 1912 5914
rect 1860 5850 1912 5856
rect 2044 5908 2096 5914
rect 2044 5850 2096 5856
rect 2332 5642 2360 6326
rect 2792 5846 2820 6394
rect 3804 6254 3832 6616
rect 3148 6248 3200 6254
rect 3792 6248 3844 6254
rect 3148 6190 3200 6196
rect 3422 6216 3478 6225
rect 2780 5840 2832 5846
rect 2780 5782 2832 5788
rect 2320 5636 2372 5642
rect 2320 5578 2372 5584
rect 1768 5364 1820 5370
rect 1768 5306 1820 5312
rect 1400 5228 1452 5234
rect 1400 5170 1452 5176
rect 2332 5030 2360 5578
rect 2792 5370 2820 5782
rect 2780 5364 2832 5370
rect 2780 5306 2832 5312
rect 2320 5024 2372 5030
rect 2320 4966 2372 4972
rect 1122 4856 1178 4865
rect 1122 4791 1178 4800
rect 2332 4554 2360 4966
rect 2792 4826 2820 5306
rect 3160 4826 3188 6190
rect 3792 6190 3844 6196
rect 3422 6151 3478 6160
rect 3436 5914 3464 6151
rect 3804 5914 3832 6190
rect 3896 6118 3924 7822
rect 4436 7812 4488 7818
rect 4436 7754 4488 7760
rect 4344 7744 4396 7750
rect 4344 7686 4396 7692
rect 4356 7478 4384 7686
rect 4344 7472 4396 7478
rect 4344 7414 4396 7420
rect 4448 7206 4476 7754
rect 4632 7324 4660 7822
rect 4724 7478 4752 8230
rect 4816 7886 4844 9959
rect 4874 9820 5182 9829
rect 4874 9818 4880 9820
rect 4936 9818 4960 9820
rect 5016 9818 5040 9820
rect 5096 9818 5120 9820
rect 5176 9818 5182 9820
rect 4936 9766 4938 9818
rect 5118 9766 5120 9818
rect 4874 9764 4880 9766
rect 4936 9764 4960 9766
rect 5016 9764 5040 9766
rect 5096 9764 5120 9766
rect 5176 9764 5182 9766
rect 4874 9755 5182 9764
rect 5080 9716 5132 9722
rect 5080 9658 5132 9664
rect 5264 9686 5316 9692
rect 4988 9580 5040 9586
rect 4988 9522 5040 9528
rect 5000 9178 5028 9522
rect 4988 9172 5040 9178
rect 4988 9114 5040 9120
rect 5092 8974 5120 9658
rect 5460 9674 5488 11018
rect 5552 9722 5580 11086
rect 5644 10062 5672 11222
rect 5816 11212 5868 11218
rect 5816 11154 5868 11160
rect 5828 10742 5856 11154
rect 6092 11144 6144 11150
rect 6092 11086 6144 11092
rect 6000 11076 6052 11082
rect 6000 11018 6052 11024
rect 5908 11008 5960 11014
rect 5908 10950 5960 10956
rect 5816 10736 5868 10742
rect 5816 10678 5868 10684
rect 5632 10056 5684 10062
rect 5632 9998 5684 10004
rect 5724 9920 5776 9926
rect 5724 9862 5776 9868
rect 5264 9628 5316 9634
rect 5368 9646 5488 9674
rect 5540 9716 5592 9722
rect 5540 9658 5592 9664
rect 5170 9616 5226 9625
rect 5170 9551 5172 9560
rect 5224 9551 5226 9560
rect 5172 9522 5224 9528
rect 5276 9466 5304 9628
rect 5368 9586 5396 9646
rect 5356 9580 5408 9586
rect 5356 9522 5408 9528
rect 5172 9444 5224 9450
rect 5276 9438 5396 9466
rect 5172 9386 5224 9392
rect 5184 9353 5212 9386
rect 5264 9376 5316 9382
rect 5170 9344 5226 9353
rect 5264 9318 5316 9324
rect 5170 9279 5226 9288
rect 5080 8968 5132 8974
rect 5080 8910 5132 8916
rect 4874 8732 5182 8741
rect 4874 8730 4880 8732
rect 4936 8730 4960 8732
rect 5016 8730 5040 8732
rect 5096 8730 5120 8732
rect 5176 8730 5182 8732
rect 4936 8678 4938 8730
rect 5118 8678 5120 8730
rect 4874 8676 4880 8678
rect 4936 8676 4960 8678
rect 5016 8676 5040 8678
rect 5096 8676 5120 8678
rect 5176 8676 5182 8678
rect 4874 8667 5182 8676
rect 5080 8356 5132 8362
rect 5080 8298 5132 8304
rect 5092 8022 5120 8298
rect 5080 8016 5132 8022
rect 5080 7958 5132 7964
rect 4804 7880 4856 7886
rect 4804 7822 4856 7828
rect 4874 7644 5182 7653
rect 4874 7642 4880 7644
rect 4936 7642 4960 7644
rect 5016 7642 5040 7644
rect 5096 7642 5120 7644
rect 5176 7642 5182 7644
rect 4936 7590 4938 7642
rect 5118 7590 5120 7642
rect 4874 7588 4880 7590
rect 4936 7588 4960 7590
rect 5016 7588 5040 7590
rect 5096 7588 5120 7590
rect 5176 7588 5182 7590
rect 4874 7579 5182 7588
rect 4712 7472 4764 7478
rect 4712 7414 4764 7420
rect 4632 7296 4752 7324
rect 4436 7200 4488 7206
rect 4436 7142 4488 7148
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 4436 6996 4488 7002
rect 4436 6938 4488 6944
rect 4160 6724 4212 6730
rect 4160 6666 4212 6672
rect 4172 6390 4200 6666
rect 4448 6390 4476 6938
rect 4620 6860 4672 6866
rect 4620 6802 4672 6808
rect 4160 6384 4212 6390
rect 4080 6344 4160 6372
rect 3884 6112 3936 6118
rect 3884 6054 3936 6060
rect 3424 5908 3476 5914
rect 3424 5850 3476 5856
rect 3792 5908 3844 5914
rect 3792 5850 3844 5856
rect 3976 5908 4028 5914
rect 3976 5850 4028 5856
rect 3332 5160 3384 5166
rect 3332 5102 3384 5108
rect 3344 4826 3372 5102
rect 3988 4826 4016 5850
rect 4080 5166 4108 6344
rect 4160 6326 4212 6332
rect 4436 6384 4488 6390
rect 4436 6326 4488 6332
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 4632 5914 4660 6802
rect 4724 6458 4752 7296
rect 4804 7200 4856 7206
rect 4804 7142 4856 7148
rect 4712 6452 4764 6458
rect 4712 6394 4764 6400
rect 4816 6186 4844 7142
rect 4874 6556 5182 6565
rect 4874 6554 4880 6556
rect 4936 6554 4960 6556
rect 5016 6554 5040 6556
rect 5096 6554 5120 6556
rect 5176 6554 5182 6556
rect 4936 6502 4938 6554
rect 5118 6502 5120 6554
rect 4874 6500 4880 6502
rect 4936 6500 4960 6502
rect 5016 6500 5040 6502
rect 5096 6500 5120 6502
rect 5176 6500 5182 6502
rect 4874 6491 5182 6500
rect 5276 6202 5304 9318
rect 5368 7002 5396 9438
rect 5460 9330 5488 9646
rect 5552 9489 5580 9658
rect 5630 9616 5686 9625
rect 5630 9551 5632 9560
rect 5684 9551 5686 9560
rect 5632 9522 5684 9528
rect 5538 9480 5594 9489
rect 5538 9415 5594 9424
rect 5460 9302 5580 9330
rect 5448 9172 5500 9178
rect 5448 9114 5500 9120
rect 5356 6996 5408 7002
rect 5356 6938 5408 6944
rect 5368 6322 5396 6938
rect 5460 6730 5488 9114
rect 5552 8634 5580 9302
rect 5644 9110 5672 9522
rect 5736 9110 5764 9862
rect 5828 9722 5856 10678
rect 5920 10130 5948 10950
rect 6012 10810 6040 11018
rect 6000 10804 6052 10810
rect 6000 10746 6052 10752
rect 5908 10124 5960 10130
rect 5908 10066 5960 10072
rect 5908 9988 5960 9994
rect 5908 9930 5960 9936
rect 5816 9716 5868 9722
rect 5816 9658 5868 9664
rect 5828 9110 5856 9658
rect 5920 9432 5948 9930
rect 6012 9586 6040 10746
rect 6104 10470 6132 11086
rect 7196 10736 7248 10742
rect 7196 10678 7248 10684
rect 6276 10600 6328 10606
rect 6276 10542 6328 10548
rect 6092 10464 6144 10470
rect 6092 10406 6144 10412
rect 6104 10266 6132 10406
rect 6288 10266 6316 10542
rect 6736 10464 6788 10470
rect 6736 10406 6788 10412
rect 6092 10260 6144 10266
rect 6092 10202 6144 10208
rect 6276 10260 6328 10266
rect 6276 10202 6328 10208
rect 6000 9580 6052 9586
rect 6000 9522 6052 9528
rect 6000 9444 6052 9450
rect 5920 9404 6000 9432
rect 6000 9386 6052 9392
rect 6012 9353 6040 9386
rect 5998 9344 6054 9353
rect 5998 9279 6054 9288
rect 6092 9172 6144 9178
rect 6092 9114 6144 9120
rect 5632 9104 5684 9110
rect 5632 9046 5684 9052
rect 5724 9104 5776 9110
rect 5724 9046 5776 9052
rect 5816 9104 5868 9110
rect 5816 9046 5868 9052
rect 5828 8922 5856 9046
rect 6104 8974 6132 9114
rect 5736 8894 5856 8922
rect 6092 8968 6144 8974
rect 6092 8910 6144 8916
rect 5540 8628 5592 8634
rect 5540 8570 5592 8576
rect 5736 8498 5764 8894
rect 5816 8832 5868 8838
rect 5816 8774 5868 8780
rect 5632 8492 5684 8498
rect 5632 8434 5684 8440
rect 5724 8492 5776 8498
rect 5724 8434 5776 8440
rect 5540 8016 5592 8022
rect 5540 7958 5592 7964
rect 5552 6866 5580 7958
rect 5644 7426 5672 8434
rect 5644 7410 5764 7426
rect 5644 7404 5776 7410
rect 5644 7398 5724 7404
rect 5644 7002 5672 7398
rect 5724 7346 5776 7352
rect 5632 6996 5684 7002
rect 5632 6938 5684 6944
rect 5540 6860 5592 6866
rect 5540 6802 5592 6808
rect 5448 6724 5500 6730
rect 5448 6666 5500 6672
rect 5356 6316 5408 6322
rect 5356 6258 5408 6264
rect 4804 6180 4856 6186
rect 4804 6122 4856 6128
rect 5184 6174 5304 6202
rect 4620 5908 4672 5914
rect 4620 5850 4672 5856
rect 5184 5778 5212 6174
rect 5264 6112 5316 6118
rect 5264 6054 5316 6060
rect 5276 5914 5304 6054
rect 5264 5908 5316 5914
rect 5264 5850 5316 5856
rect 5172 5772 5224 5778
rect 5172 5714 5224 5720
rect 4620 5636 4672 5642
rect 4620 5578 4672 5584
rect 4344 5568 4396 5574
rect 4344 5510 4396 5516
rect 4068 5160 4120 5166
rect 4068 5102 4120 5108
rect 2780 4820 2832 4826
rect 2780 4762 2832 4768
rect 3148 4820 3200 4826
rect 3148 4762 3200 4768
rect 3332 4820 3384 4826
rect 3332 4762 3384 4768
rect 3976 4820 4028 4826
rect 3976 4762 4028 4768
rect 1676 4548 1728 4554
rect 1676 4490 1728 4496
rect 2320 4548 2372 4554
rect 2320 4490 2372 4496
rect 1688 4282 1716 4490
rect 4080 4282 4108 5102
rect 4356 5098 4384 5510
rect 4344 5092 4396 5098
rect 4344 5034 4396 5040
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 4632 4690 4660 5578
rect 4804 5568 4856 5574
rect 4804 5510 4856 5516
rect 4712 5160 4764 5166
rect 4712 5102 4764 5108
rect 4724 4826 4752 5102
rect 4712 4820 4764 4826
rect 4712 4762 4764 4768
rect 4816 4758 4844 5510
rect 4874 5468 5182 5477
rect 4874 5466 4880 5468
rect 4936 5466 4960 5468
rect 5016 5466 5040 5468
rect 5096 5466 5120 5468
rect 5176 5466 5182 5468
rect 4936 5414 4938 5466
rect 5118 5414 5120 5466
rect 4874 5412 4880 5414
rect 4936 5412 4960 5414
rect 5016 5412 5040 5414
rect 5096 5412 5120 5414
rect 5176 5412 5182 5414
rect 4874 5403 5182 5412
rect 4804 4752 4856 4758
rect 4804 4694 4856 4700
rect 4620 4684 4672 4690
rect 4620 4626 4672 4632
rect 4436 4480 4488 4486
rect 4436 4422 4488 4428
rect 1676 4276 1728 4282
rect 1676 4218 1728 4224
rect 4068 4276 4120 4282
rect 4068 4218 4120 4224
rect 4448 4214 4476 4422
rect 4816 4282 4844 4694
rect 4874 4380 5182 4389
rect 4874 4378 4880 4380
rect 4936 4378 4960 4380
rect 5016 4378 5040 4380
rect 5096 4378 5120 4380
rect 5176 4378 5182 4380
rect 4936 4326 4938 4378
rect 5118 4326 5120 4378
rect 4874 4324 4880 4326
rect 4936 4324 4960 4326
rect 5016 4324 5040 4326
rect 5096 4324 5120 4326
rect 5176 4324 5182 4326
rect 4874 4315 5182 4324
rect 4804 4276 4856 4282
rect 4804 4218 4856 4224
rect 4436 4208 4488 4214
rect 1490 4176 1546 4185
rect 4436 4150 4488 4156
rect 1490 4111 1546 4120
rect 2044 4140 2096 4146
rect 1504 4010 1532 4111
rect 2044 4082 2096 4088
rect 1492 4004 1544 4010
rect 1492 3946 1544 3952
rect 2056 3738 2084 4082
rect 5368 4078 5396 6258
rect 5460 5914 5488 6666
rect 5828 6372 5856 8774
rect 6184 8492 6236 8498
rect 6184 8434 6236 8440
rect 6000 8424 6052 8430
rect 6000 8366 6052 8372
rect 6012 6798 6040 8366
rect 6092 7744 6144 7750
rect 6092 7686 6144 7692
rect 6104 7546 6132 7686
rect 6196 7546 6224 8434
rect 6288 8090 6316 10202
rect 6748 9994 6776 10406
rect 6460 9988 6512 9994
rect 6460 9930 6512 9936
rect 6736 9988 6788 9994
rect 6736 9930 6788 9936
rect 6472 9722 6500 9930
rect 6644 9920 6696 9926
rect 6644 9862 6696 9868
rect 6656 9722 6684 9862
rect 6460 9716 6512 9722
rect 6460 9658 6512 9664
rect 6644 9716 6696 9722
rect 6644 9658 6696 9664
rect 6656 9586 6684 9658
rect 6644 9580 6696 9586
rect 6644 9522 6696 9528
rect 6642 9480 6698 9489
rect 6642 9415 6698 9424
rect 6656 9382 6684 9415
rect 6644 9376 6696 9382
rect 6644 9318 6696 9324
rect 6368 9104 6420 9110
rect 6368 9046 6420 9052
rect 6276 8084 6328 8090
rect 6276 8026 6328 8032
rect 6276 7744 6328 7750
rect 6276 7686 6328 7692
rect 6092 7540 6144 7546
rect 6092 7482 6144 7488
rect 6184 7540 6236 7546
rect 6184 7482 6236 7488
rect 6288 7410 6316 7686
rect 6276 7404 6328 7410
rect 6276 7346 6328 7352
rect 6276 7268 6328 7274
rect 6276 7210 6328 7216
rect 6000 6792 6052 6798
rect 6000 6734 6052 6740
rect 6288 6458 6316 7210
rect 6380 7206 6408 9046
rect 6460 8832 6512 8838
rect 6460 8774 6512 8780
rect 6368 7200 6420 7206
rect 6368 7142 6420 7148
rect 6276 6452 6328 6458
rect 6276 6394 6328 6400
rect 5908 6384 5960 6390
rect 5828 6344 5908 6372
rect 5908 6326 5960 6332
rect 6380 6338 6408 7142
rect 6472 6866 6500 8774
rect 6656 8634 6684 9318
rect 6644 8628 6696 8634
rect 6644 8570 6696 8576
rect 6748 7750 6776 9930
rect 7012 9172 7064 9178
rect 7012 9114 7064 9120
rect 6920 8832 6972 8838
rect 6920 8774 6972 8780
rect 6932 8294 6960 8774
rect 6920 8288 6972 8294
rect 6920 8230 6972 8236
rect 6920 7812 6972 7818
rect 6920 7754 6972 7760
rect 6736 7744 6788 7750
rect 6736 7686 6788 7692
rect 6932 7546 6960 7754
rect 6920 7540 6972 7546
rect 6920 7482 6972 7488
rect 6828 7404 6880 7410
rect 6828 7346 6880 7352
rect 6840 7206 6868 7346
rect 7024 7274 7052 9114
rect 7208 8566 7236 10678
rect 7380 10600 7432 10606
rect 7380 10542 7432 10548
rect 7392 9722 7420 10542
rect 8116 10464 8168 10470
rect 8116 10406 8168 10412
rect 8208 10464 8260 10470
rect 8208 10406 8260 10412
rect 7656 10124 7708 10130
rect 7656 10066 7708 10072
rect 7472 9920 7524 9926
rect 7472 9862 7524 9868
rect 7380 9716 7432 9722
rect 7380 9658 7432 9664
rect 7484 9518 7512 9862
rect 7668 9654 7696 10066
rect 8128 9994 8156 10406
rect 8116 9988 8168 9994
rect 8116 9930 8168 9936
rect 8024 9920 8076 9926
rect 8024 9862 8076 9868
rect 8036 9722 8064 9862
rect 8024 9716 8076 9722
rect 8128 9697 8156 9930
rect 8024 9658 8076 9664
rect 8114 9688 8170 9697
rect 7656 9648 7708 9654
rect 7564 9602 7616 9608
rect 8114 9623 8116 9632
rect 7656 9590 7708 9596
rect 8168 9623 8170 9632
rect 8116 9590 8168 9596
rect 8220 9586 8248 10406
rect 9036 9988 9088 9994
rect 9036 9930 9088 9936
rect 8300 9920 8352 9926
rect 8300 9862 8352 9868
rect 8312 9674 8340 9862
rect 8312 9646 8524 9674
rect 7564 9544 7616 9550
rect 8208 9580 8260 9586
rect 7472 9512 7524 9518
rect 7392 9472 7472 9500
rect 7392 8974 7420 9472
rect 7472 9454 7524 9460
rect 7576 9110 7604 9544
rect 8208 9522 8260 9528
rect 8392 9580 8444 9586
rect 8392 9522 8444 9528
rect 8022 9480 8078 9489
rect 8022 9415 8078 9424
rect 7564 9104 7616 9110
rect 7564 9046 7616 9052
rect 7380 8968 7432 8974
rect 7380 8910 7432 8916
rect 8036 8838 8064 9415
rect 8404 9178 8432 9522
rect 8392 9172 8444 9178
rect 8392 9114 8444 9120
rect 8300 8968 8352 8974
rect 8300 8910 8352 8916
rect 8024 8832 8076 8838
rect 8024 8774 8076 8780
rect 7196 8560 7248 8566
rect 7196 8502 7248 8508
rect 7208 7818 7236 8502
rect 7196 7812 7248 7818
rect 7196 7754 7248 7760
rect 7748 7744 7800 7750
rect 7748 7686 7800 7692
rect 7288 7404 7340 7410
rect 7288 7346 7340 7352
rect 7012 7268 7064 7274
rect 7012 7210 7064 7216
rect 6828 7200 6880 7206
rect 6828 7142 6880 7148
rect 6552 6996 6604 7002
rect 6552 6938 6604 6944
rect 6460 6860 6512 6866
rect 6460 6802 6512 6808
rect 6564 6458 6592 6938
rect 6840 6934 6868 7142
rect 7300 7002 7328 7346
rect 7472 7200 7524 7206
rect 7472 7142 7524 7148
rect 7564 7200 7616 7206
rect 7564 7142 7616 7148
rect 6920 6996 6972 7002
rect 6920 6938 6972 6944
rect 7288 6996 7340 7002
rect 7288 6938 7340 6944
rect 6828 6928 6880 6934
rect 6828 6870 6880 6876
rect 6828 6792 6880 6798
rect 6932 6780 6960 6938
rect 6880 6752 6960 6780
rect 7288 6792 7340 6798
rect 6828 6734 6880 6740
rect 7288 6734 7340 6740
rect 6736 6656 6788 6662
rect 6736 6598 6788 6604
rect 6552 6452 6604 6458
rect 6552 6394 6604 6400
rect 6644 6452 6696 6458
rect 6644 6394 6696 6400
rect 6656 6338 6684 6394
rect 6748 6390 6776 6598
rect 6184 6316 6236 6322
rect 6184 6258 6236 6264
rect 6380 6310 6684 6338
rect 6736 6384 6788 6390
rect 6736 6326 6788 6332
rect 5448 5908 5500 5914
rect 5448 5850 5500 5856
rect 6092 5636 6144 5642
rect 6092 5578 6144 5584
rect 6104 5166 6132 5578
rect 6196 5370 6224 6258
rect 6276 5568 6328 5574
rect 6276 5510 6328 5516
rect 6288 5370 6316 5510
rect 6184 5364 6236 5370
rect 6184 5306 6236 5312
rect 6276 5364 6328 5370
rect 6276 5306 6328 5312
rect 6092 5160 6144 5166
rect 6092 5102 6144 5108
rect 5540 4616 5592 4622
rect 5540 4558 5592 4564
rect 5356 4072 5408 4078
rect 5356 4014 5408 4020
rect 5552 4010 5580 4558
rect 5908 4480 5960 4486
rect 5908 4422 5960 4428
rect 5920 4282 5948 4422
rect 5908 4276 5960 4282
rect 5908 4218 5960 4224
rect 6104 4078 6132 5102
rect 6196 4690 6224 5306
rect 6380 5098 6408 6310
rect 6840 6186 6868 6734
rect 7196 6656 7248 6662
rect 7196 6598 7248 6604
rect 7208 6322 7236 6598
rect 7300 6322 7328 6734
rect 7380 6656 7432 6662
rect 7380 6598 7432 6604
rect 7196 6316 7248 6322
rect 7196 6258 7248 6264
rect 7288 6316 7340 6322
rect 7288 6258 7340 6264
rect 6920 6248 6972 6254
rect 7300 6202 7328 6258
rect 6920 6190 6972 6196
rect 6828 6180 6880 6186
rect 6828 6122 6880 6128
rect 6736 6112 6788 6118
rect 6736 6054 6788 6060
rect 6644 5636 6696 5642
rect 6644 5578 6696 5584
rect 6656 5370 6684 5578
rect 6644 5364 6696 5370
rect 6644 5306 6696 5312
rect 6748 5098 6776 6054
rect 6932 5166 6960 6190
rect 7104 6180 7156 6186
rect 7104 6122 7156 6128
rect 7208 6174 7328 6202
rect 7392 6186 7420 6598
rect 7380 6180 7432 6186
rect 7116 5574 7144 6122
rect 7208 5914 7236 6174
rect 7380 6122 7432 6128
rect 7288 6112 7340 6118
rect 7288 6054 7340 6060
rect 7196 5908 7248 5914
rect 7196 5850 7248 5856
rect 7104 5568 7156 5574
rect 7104 5510 7156 5516
rect 6920 5160 6972 5166
rect 6920 5102 6972 5108
rect 6368 5092 6420 5098
rect 6368 5034 6420 5040
rect 6644 5092 6696 5098
rect 6644 5034 6696 5040
rect 6736 5092 6788 5098
rect 6736 5034 6788 5040
rect 6828 5092 6880 5098
rect 6828 5034 6880 5040
rect 6184 4684 6236 4690
rect 6184 4626 6236 4632
rect 6656 4622 6684 5034
rect 6748 4758 6776 5034
rect 6840 4826 6868 5034
rect 6932 4826 6960 5102
rect 6828 4820 6880 4826
rect 6828 4762 6880 4768
rect 6920 4820 6972 4826
rect 6920 4762 6972 4768
rect 6736 4752 6788 4758
rect 6736 4694 6788 4700
rect 7116 4690 7144 5510
rect 7104 4684 7156 4690
rect 7104 4626 7156 4632
rect 6644 4616 6696 4622
rect 6644 4558 6696 4564
rect 7104 4480 7156 4486
rect 7104 4422 7156 4428
rect 7116 4282 7144 4422
rect 7104 4276 7156 4282
rect 7104 4218 7156 4224
rect 7300 4078 7328 6054
rect 7484 5574 7512 7142
rect 7472 5568 7524 5574
rect 7472 5510 7524 5516
rect 7576 5370 7604 7142
rect 7760 5642 7788 7686
rect 7932 7404 7984 7410
rect 7932 7346 7984 7352
rect 7944 7206 7972 7346
rect 7932 7200 7984 7206
rect 7932 7142 7984 7148
rect 7840 6860 7892 6866
rect 7840 6802 7892 6808
rect 7852 6662 7880 6802
rect 7840 6656 7892 6662
rect 7840 6598 7892 6604
rect 7748 5636 7800 5642
rect 7748 5578 7800 5584
rect 7760 5370 7788 5578
rect 7564 5364 7616 5370
rect 7564 5306 7616 5312
rect 7748 5364 7800 5370
rect 7748 5306 7800 5312
rect 7760 5114 7788 5306
rect 7576 5098 7788 5114
rect 7564 5092 7788 5098
rect 7616 5086 7788 5092
rect 7564 5034 7616 5040
rect 7852 4622 7880 6598
rect 7944 4826 7972 7142
rect 8036 6934 8064 8774
rect 8312 8634 8340 8910
rect 8300 8628 8352 8634
rect 8300 8570 8352 8576
rect 8404 8022 8432 9114
rect 8496 9110 8524 9646
rect 8760 9444 8812 9450
rect 8760 9386 8812 9392
rect 8484 9104 8536 9110
rect 8484 9046 8536 9052
rect 8668 9036 8720 9042
rect 8668 8978 8720 8984
rect 8576 8832 8628 8838
rect 8576 8774 8628 8780
rect 8588 8634 8616 8774
rect 8680 8634 8708 8978
rect 8772 8974 8800 9386
rect 8852 9376 8904 9382
rect 8852 9318 8904 9324
rect 8760 8968 8812 8974
rect 8760 8910 8812 8916
rect 8576 8628 8628 8634
rect 8576 8570 8628 8576
rect 8668 8628 8720 8634
rect 8668 8570 8720 8576
rect 8484 8492 8536 8498
rect 8484 8434 8536 8440
rect 8392 8016 8444 8022
rect 8392 7958 8444 7964
rect 8496 7954 8524 8434
rect 8484 7948 8536 7954
rect 8484 7890 8536 7896
rect 8496 7546 8524 7890
rect 8484 7540 8536 7546
rect 8484 7482 8536 7488
rect 8024 6928 8076 6934
rect 8024 6870 8076 6876
rect 8300 6928 8352 6934
rect 8300 6870 8352 6876
rect 8116 6656 8168 6662
rect 8116 6598 8168 6604
rect 8128 6458 8156 6598
rect 8116 6452 8168 6458
rect 8116 6394 8168 6400
rect 8312 5250 8340 6870
rect 8392 6112 8444 6118
rect 8392 6054 8444 6060
rect 8404 5914 8432 6054
rect 8392 5908 8444 5914
rect 8392 5850 8444 5856
rect 8496 5778 8524 7482
rect 8772 6866 8800 8910
rect 8864 8498 8892 9318
rect 9048 8634 9076 9930
rect 9128 9580 9180 9586
rect 9128 9522 9180 9528
rect 9036 8628 9088 8634
rect 9036 8570 9088 8576
rect 8852 8492 8904 8498
rect 8852 8434 8904 8440
rect 8944 7744 8996 7750
rect 8944 7686 8996 7692
rect 8956 7478 8984 7686
rect 8944 7472 8996 7478
rect 8944 7414 8996 7420
rect 8760 6860 8812 6866
rect 8760 6802 8812 6808
rect 9048 6730 9076 8570
rect 9140 6798 9168 9522
rect 9128 6792 9180 6798
rect 9128 6734 9180 6740
rect 9036 6724 9088 6730
rect 9036 6666 9088 6672
rect 8484 5772 8536 5778
rect 8484 5714 8536 5720
rect 8496 5370 8524 5714
rect 10508 5636 10560 5642
rect 10508 5578 10560 5584
rect 10520 5545 10548 5578
rect 10506 5536 10562 5545
rect 10506 5471 10562 5480
rect 8484 5364 8536 5370
rect 8484 5306 8536 5312
rect 8220 5222 8340 5250
rect 8220 5166 8248 5222
rect 8208 5160 8260 5166
rect 8208 5102 8260 5108
rect 8576 5160 8628 5166
rect 8576 5102 8628 5108
rect 7932 4820 7984 4826
rect 7932 4762 7984 4768
rect 7840 4616 7892 4622
rect 7840 4558 7892 4564
rect 8588 4078 8616 5102
rect 6092 4072 6144 4078
rect 6092 4014 6144 4020
rect 7288 4072 7340 4078
rect 7288 4014 7340 4020
rect 8576 4072 8628 4078
rect 8576 4014 8628 4020
rect 5540 4004 5592 4010
rect 5540 3946 5592 3952
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 2044 3732 2096 3738
rect 2044 3674 2096 3680
rect 5724 3596 5776 3602
rect 5724 3538 5776 3544
rect 940 3528 992 3534
rect 938 3496 940 3505
rect 3976 3528 4028 3534
rect 992 3496 994 3505
rect 3976 3470 4028 3476
rect 4620 3528 4672 3534
rect 4620 3470 4672 3476
rect 938 3431 994 3440
rect 3884 3392 3936 3398
rect 3884 3334 3936 3340
rect 2964 2984 3016 2990
rect 2964 2926 3016 2932
rect 2976 2514 3004 2926
rect 2964 2508 3016 2514
rect 2964 2450 3016 2456
rect 2688 2440 2740 2446
rect 2608 2400 2688 2428
rect 2608 800 2636 2400
rect 2688 2382 2740 2388
rect 3240 2440 3292 2446
rect 3240 2382 3292 2388
rect 3252 800 3280 2382
rect 3896 800 3924 3334
rect 3988 3194 4016 3470
rect 4632 3194 4660 3470
rect 4804 3392 4856 3398
rect 4804 3334 4856 3340
rect 5356 3392 5408 3398
rect 5356 3334 5408 3340
rect 3976 3188 4028 3194
rect 3976 3130 4028 3136
rect 4620 3188 4672 3194
rect 4620 3130 4672 3136
rect 4816 3074 4844 3334
rect 4874 3292 5182 3301
rect 4874 3290 4880 3292
rect 4936 3290 4960 3292
rect 5016 3290 5040 3292
rect 5096 3290 5120 3292
rect 5176 3290 5182 3292
rect 4936 3238 4938 3290
rect 5118 3238 5120 3290
rect 4874 3236 4880 3238
rect 4936 3236 4960 3238
rect 5016 3236 5040 3238
rect 5096 3236 5120 3238
rect 5176 3236 5182 3238
rect 4874 3227 5182 3236
rect 4436 3052 4488 3058
rect 4436 2994 4488 3000
rect 4632 3046 4844 3074
rect 3976 2984 4028 2990
rect 3976 2926 4028 2932
rect 3988 2514 4016 2926
rect 4448 2922 4476 2994
rect 4436 2916 4488 2922
rect 4436 2858 4488 2864
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 3976 2508 4028 2514
rect 3976 2450 4028 2456
rect 4632 1714 4660 3046
rect 4804 2848 4856 2854
rect 4804 2790 4856 2796
rect 4816 2446 4844 2790
rect 5368 2446 5396 3334
rect 5736 2990 5764 3538
rect 5908 3528 5960 3534
rect 5908 3470 5960 3476
rect 5920 3194 5948 3470
rect 6000 3460 6052 3466
rect 6000 3402 6052 3408
rect 5908 3188 5960 3194
rect 5908 3130 5960 3136
rect 5724 2984 5776 2990
rect 5724 2926 5776 2932
rect 5736 2650 5764 2926
rect 5920 2854 5948 3130
rect 6012 3126 6040 3402
rect 6092 3392 6144 3398
rect 6092 3334 6144 3340
rect 6000 3120 6052 3126
rect 6000 3062 6052 3068
rect 5908 2848 5960 2854
rect 5908 2790 5960 2796
rect 5724 2644 5776 2650
rect 5724 2586 5776 2592
rect 5920 2582 5948 2790
rect 5908 2576 5960 2582
rect 5908 2518 5960 2524
rect 4804 2440 4856 2446
rect 4804 2382 4856 2388
rect 5356 2440 5408 2446
rect 5356 2382 5408 2388
rect 6012 2378 6040 3062
rect 6104 2446 6132 3334
rect 7288 3188 7340 3194
rect 7288 3130 7340 3136
rect 6920 2848 6972 2854
rect 6920 2790 6972 2796
rect 6932 2446 6960 2790
rect 7300 2446 7328 3130
rect 9404 3120 9456 3126
rect 9404 3062 9456 3068
rect 9416 2514 9444 3062
rect 9404 2508 9456 2514
rect 9404 2450 9456 2456
rect 6092 2440 6144 2446
rect 6092 2382 6144 2388
rect 6920 2440 6972 2446
rect 6920 2382 6972 2388
rect 7288 2440 7340 2446
rect 7288 2382 7340 2388
rect 9128 2440 9180 2446
rect 9128 2382 9180 2388
rect 6000 2372 6052 2378
rect 6000 2314 6052 2320
rect 5080 2304 5132 2310
rect 5816 2304 5868 2310
rect 5132 2264 5304 2292
rect 5080 2246 5132 2252
rect 4874 2204 5182 2213
rect 4874 2202 4880 2204
rect 4936 2202 4960 2204
rect 5016 2202 5040 2204
rect 5096 2202 5120 2204
rect 5176 2202 5182 2204
rect 4936 2150 4938 2202
rect 5118 2150 5120 2202
rect 4874 2148 4880 2150
rect 4936 2148 4960 2150
rect 5016 2148 5040 2150
rect 5096 2148 5120 2150
rect 5176 2148 5182 2150
rect 4874 2139 5182 2148
rect 4540 1686 4660 1714
rect 4540 800 4568 1686
rect 5276 1170 5304 2264
rect 5816 2246 5868 2252
rect 6460 2304 6512 2310
rect 6460 2246 6512 2252
rect 7104 2304 7156 2310
rect 7104 2246 7156 2252
rect 7748 2304 7800 2310
rect 7748 2246 7800 2252
rect 8392 2304 8444 2310
rect 8392 2246 8444 2252
rect 5184 1142 5304 1170
rect 5184 800 5212 1142
rect 5828 800 5856 2246
rect 6472 800 6500 2246
rect 7116 800 7144 2246
rect 7760 800 7788 2246
rect 8404 800 8432 2246
rect 9140 1306 9168 2382
rect 9048 1278 9168 1306
rect 9048 800 9076 1278
rect 2594 0 2650 800
rect 3238 0 3294 800
rect 3882 0 3938 800
rect 4526 0 4582 800
rect 5170 0 5226 800
rect 5814 0 5870 800
rect 6458 0 6514 800
rect 7102 0 7158 800
rect 7746 0 7802 800
rect 8390 0 8446 800
rect 9034 0 9090 800
<< via2 >>
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 1122 8200 1178 8256
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 1398 7520 1454 7576
rect 4880 10906 4936 10908
rect 4960 10906 5016 10908
rect 5040 10906 5096 10908
rect 5120 10906 5176 10908
rect 4880 10854 4926 10906
rect 4926 10854 4936 10906
rect 4960 10854 4990 10906
rect 4990 10854 5002 10906
rect 5002 10854 5016 10906
rect 5040 10854 5054 10906
rect 5054 10854 5066 10906
rect 5066 10854 5096 10906
rect 5120 10854 5130 10906
rect 5130 10854 5176 10906
rect 4880 10852 4936 10854
rect 4960 10852 5016 10854
rect 5040 10852 5096 10854
rect 5120 10852 5176 10854
rect 4802 9968 4858 10024
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4434 9016 4490 9072
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 3330 6840 3386 6896
rect 1398 5480 1454 5536
rect 1122 4800 1178 4856
rect 3422 6160 3478 6216
rect 4880 9818 4936 9820
rect 4960 9818 5016 9820
rect 5040 9818 5096 9820
rect 5120 9818 5176 9820
rect 4880 9766 4926 9818
rect 4926 9766 4936 9818
rect 4960 9766 4990 9818
rect 4990 9766 5002 9818
rect 5002 9766 5016 9818
rect 5040 9766 5054 9818
rect 5054 9766 5066 9818
rect 5066 9766 5096 9818
rect 5120 9766 5130 9818
rect 5130 9766 5176 9818
rect 4880 9764 4936 9766
rect 4960 9764 5016 9766
rect 5040 9764 5096 9766
rect 5120 9764 5176 9766
rect 5170 9580 5226 9616
rect 5170 9560 5172 9580
rect 5172 9560 5224 9580
rect 5224 9560 5226 9580
rect 5170 9288 5226 9344
rect 4880 8730 4936 8732
rect 4960 8730 5016 8732
rect 5040 8730 5096 8732
rect 5120 8730 5176 8732
rect 4880 8678 4926 8730
rect 4926 8678 4936 8730
rect 4960 8678 4990 8730
rect 4990 8678 5002 8730
rect 5002 8678 5016 8730
rect 5040 8678 5054 8730
rect 5054 8678 5066 8730
rect 5066 8678 5096 8730
rect 5120 8678 5130 8730
rect 5130 8678 5176 8730
rect 4880 8676 4936 8678
rect 4960 8676 5016 8678
rect 5040 8676 5096 8678
rect 5120 8676 5176 8678
rect 4880 7642 4936 7644
rect 4960 7642 5016 7644
rect 5040 7642 5096 7644
rect 5120 7642 5176 7644
rect 4880 7590 4926 7642
rect 4926 7590 4936 7642
rect 4960 7590 4990 7642
rect 4990 7590 5002 7642
rect 5002 7590 5016 7642
rect 5040 7590 5054 7642
rect 5054 7590 5066 7642
rect 5066 7590 5096 7642
rect 5120 7590 5130 7642
rect 5130 7590 5176 7642
rect 4880 7588 4936 7590
rect 4960 7588 5016 7590
rect 5040 7588 5096 7590
rect 5120 7588 5176 7590
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4880 6554 4936 6556
rect 4960 6554 5016 6556
rect 5040 6554 5096 6556
rect 5120 6554 5176 6556
rect 4880 6502 4926 6554
rect 4926 6502 4936 6554
rect 4960 6502 4990 6554
rect 4990 6502 5002 6554
rect 5002 6502 5016 6554
rect 5040 6502 5054 6554
rect 5054 6502 5066 6554
rect 5066 6502 5096 6554
rect 5120 6502 5130 6554
rect 5130 6502 5176 6554
rect 4880 6500 4936 6502
rect 4960 6500 5016 6502
rect 5040 6500 5096 6502
rect 5120 6500 5176 6502
rect 5630 9580 5686 9616
rect 5630 9560 5632 9580
rect 5632 9560 5684 9580
rect 5684 9560 5686 9580
rect 5538 9424 5594 9480
rect 5998 9288 6054 9344
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4880 5466 4936 5468
rect 4960 5466 5016 5468
rect 5040 5466 5096 5468
rect 5120 5466 5176 5468
rect 4880 5414 4926 5466
rect 4926 5414 4936 5466
rect 4960 5414 4990 5466
rect 4990 5414 5002 5466
rect 5002 5414 5016 5466
rect 5040 5414 5054 5466
rect 5054 5414 5066 5466
rect 5066 5414 5096 5466
rect 5120 5414 5130 5466
rect 5130 5414 5176 5466
rect 4880 5412 4936 5414
rect 4960 5412 5016 5414
rect 5040 5412 5096 5414
rect 5120 5412 5176 5414
rect 4880 4378 4936 4380
rect 4960 4378 5016 4380
rect 5040 4378 5096 4380
rect 5120 4378 5176 4380
rect 4880 4326 4926 4378
rect 4926 4326 4936 4378
rect 4960 4326 4990 4378
rect 4990 4326 5002 4378
rect 5002 4326 5016 4378
rect 5040 4326 5054 4378
rect 5054 4326 5066 4378
rect 5066 4326 5096 4378
rect 5120 4326 5130 4378
rect 5130 4326 5176 4378
rect 4880 4324 4936 4326
rect 4960 4324 5016 4326
rect 5040 4324 5096 4326
rect 5120 4324 5176 4326
rect 1490 4120 1546 4176
rect 6642 9424 6698 9480
rect 8114 9648 8170 9688
rect 8114 9632 8116 9648
rect 8116 9632 8168 9648
rect 8168 9632 8170 9648
rect 8022 9424 8078 9480
rect 10506 5480 10562 5536
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 938 3476 940 3496
rect 940 3476 992 3496
rect 992 3476 994 3496
rect 938 3440 994 3476
rect 4880 3290 4936 3292
rect 4960 3290 5016 3292
rect 5040 3290 5096 3292
rect 5120 3290 5176 3292
rect 4880 3238 4926 3290
rect 4926 3238 4936 3290
rect 4960 3238 4990 3290
rect 4990 3238 5002 3290
rect 5002 3238 5016 3290
rect 5040 3238 5054 3290
rect 5054 3238 5066 3290
rect 5066 3238 5096 3290
rect 5120 3238 5130 3290
rect 5130 3238 5176 3290
rect 4880 3236 4936 3238
rect 4960 3236 5016 3238
rect 5040 3236 5096 3238
rect 5120 3236 5176 3238
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 4880 2202 4936 2204
rect 4960 2202 5016 2204
rect 5040 2202 5096 2204
rect 5120 2202 5176 2204
rect 4880 2150 4926 2202
rect 4926 2150 4936 2202
rect 4960 2150 4990 2202
rect 4990 2150 5002 2202
rect 5002 2150 5016 2202
rect 5040 2150 5054 2202
rect 5054 2150 5066 2202
rect 5066 2150 5096 2202
rect 5120 2150 5130 2202
rect 5130 2150 5176 2202
rect 4880 2148 4936 2150
rect 4960 2148 5016 2150
rect 5040 2148 5096 2150
rect 5120 2148 5176 2150
<< metal3 >>
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 4870 10912 5186 10913
rect 4870 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5186 10912
rect 4870 10847 5186 10848
rect 4210 10368 4526 10369
rect 0 10298 800 10328
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 0 10238 2790 10298
rect 0 10208 800 10238
rect 2730 10026 2790 10238
rect 4797 10026 4863 10029
rect 2730 10024 4863 10026
rect 2730 9968 4802 10024
rect 4858 9968 4863 10024
rect 2730 9966 4863 9968
rect 4797 9963 4863 9966
rect 4870 9824 5186 9825
rect 4870 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5186 9824
rect 4870 9759 5186 9760
rect 8109 9690 8175 9693
rect 8109 9688 8218 9690
rect 8109 9632 8114 9688
rect 8170 9632 8218 9688
rect 8109 9627 8218 9632
rect 5165 9618 5231 9621
rect 5625 9618 5691 9621
rect 5165 9616 5691 9618
rect 5165 9560 5170 9616
rect 5226 9560 5630 9616
rect 5686 9560 5691 9616
rect 5165 9558 5691 9560
rect 5165 9555 5231 9558
rect 5625 9555 5691 9558
rect 5533 9482 5599 9485
rect 6637 9482 6703 9485
rect 4662 9480 6703 9482
rect 4662 9424 5538 9480
rect 5594 9424 6642 9480
rect 6698 9424 6703 9480
rect 4662 9422 6703 9424
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 4429 9074 4495 9077
rect 4662 9074 4722 9422
rect 5533 9419 5599 9422
rect 6637 9419 6703 9422
rect 8017 9482 8083 9485
rect 8158 9482 8218 9627
rect 8017 9480 8218 9482
rect 8017 9424 8022 9480
rect 8078 9424 8218 9480
rect 8017 9422 8218 9424
rect 8017 9419 8083 9422
rect 5165 9346 5231 9349
rect 5993 9346 6059 9349
rect 5165 9344 6059 9346
rect 5165 9288 5170 9344
rect 5226 9288 5998 9344
rect 6054 9288 6059 9344
rect 5165 9286 6059 9288
rect 5165 9283 5231 9286
rect 5993 9283 6059 9286
rect 4429 9072 4722 9074
rect 4429 9016 4434 9072
rect 4490 9016 4722 9072
rect 4429 9014 4722 9016
rect 4429 9011 4495 9014
rect 4870 8736 5186 8737
rect 4870 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5186 8736
rect 4870 8671 5186 8672
rect 0 8258 800 8288
rect 1117 8258 1183 8261
rect 0 8256 1183 8258
rect 0 8200 1122 8256
rect 1178 8200 1183 8256
rect 0 8198 1183 8200
rect 0 8168 800 8198
rect 1117 8195 1183 8198
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 4870 7648 5186 7649
rect 0 7578 800 7608
rect 4870 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5186 7648
rect 4870 7583 5186 7584
rect 1393 7578 1459 7581
rect 0 7576 1459 7578
rect 0 7520 1398 7576
rect 1454 7520 1459 7576
rect 0 7518 1459 7520
rect 0 7488 800 7518
rect 1393 7515 1459 7518
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 0 6898 800 6928
rect 3325 6898 3391 6901
rect 0 6896 3391 6898
rect 0 6840 3330 6896
rect 3386 6840 3391 6896
rect 0 6838 3391 6840
rect 0 6808 800 6838
rect 3325 6835 3391 6838
rect 4870 6560 5186 6561
rect 4870 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5186 6560
rect 4870 6495 5186 6496
rect 0 6218 800 6248
rect 3417 6218 3483 6221
rect 0 6216 3483 6218
rect 0 6160 3422 6216
rect 3478 6160 3483 6216
rect 0 6158 3483 6160
rect 0 6128 800 6158
rect 3417 6155 3483 6158
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 0 5538 800 5568
rect 1393 5538 1459 5541
rect 0 5536 1459 5538
rect 0 5480 1398 5536
rect 1454 5480 1459 5536
rect 0 5478 1459 5480
rect 0 5448 800 5478
rect 1393 5475 1459 5478
rect 10501 5538 10567 5541
rect 10793 5538 11593 5568
rect 10501 5536 11593 5538
rect 10501 5480 10506 5536
rect 10562 5480 11593 5536
rect 10501 5478 11593 5480
rect 10501 5475 10567 5478
rect 4870 5472 5186 5473
rect 4870 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5186 5472
rect 10793 5448 11593 5478
rect 4870 5407 5186 5408
rect 4210 4928 4526 4929
rect 0 4858 800 4888
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 1117 4858 1183 4861
rect 0 4856 1183 4858
rect 0 4800 1122 4856
rect 1178 4800 1183 4856
rect 0 4798 1183 4800
rect 0 4768 800 4798
rect 1117 4795 1183 4798
rect 4870 4384 5186 4385
rect 4870 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5186 4384
rect 4870 4319 5186 4320
rect 0 4178 800 4208
rect 1485 4178 1551 4181
rect 0 4176 1551 4178
rect 0 4120 1490 4176
rect 1546 4120 1551 4176
rect 0 4118 1551 4120
rect 0 4088 800 4118
rect 1485 4115 1551 4118
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 798 3574 1042 3634
rect 798 3528 858 3574
rect 0 3438 858 3528
rect 982 3501 1042 3574
rect 933 3496 1042 3501
rect 933 3440 938 3496
rect 994 3440 1042 3496
rect 933 3438 1042 3440
rect 0 3408 800 3438
rect 933 3435 999 3438
rect 4870 3296 5186 3297
rect 4870 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5186 3296
rect 4870 3231 5186 3232
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 4870 2208 5186 2209
rect 4870 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5186 2208
rect 4870 2143 5186 2144
<< via3 >>
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 4876 10908 4940 10912
rect 4876 10852 4880 10908
rect 4880 10852 4936 10908
rect 4936 10852 4940 10908
rect 4876 10848 4940 10852
rect 4956 10908 5020 10912
rect 4956 10852 4960 10908
rect 4960 10852 5016 10908
rect 5016 10852 5020 10908
rect 4956 10848 5020 10852
rect 5036 10908 5100 10912
rect 5036 10852 5040 10908
rect 5040 10852 5096 10908
rect 5096 10852 5100 10908
rect 5036 10848 5100 10852
rect 5116 10908 5180 10912
rect 5116 10852 5120 10908
rect 5120 10852 5176 10908
rect 5176 10852 5180 10908
rect 5116 10848 5180 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 4876 9820 4940 9824
rect 4876 9764 4880 9820
rect 4880 9764 4936 9820
rect 4936 9764 4940 9820
rect 4876 9760 4940 9764
rect 4956 9820 5020 9824
rect 4956 9764 4960 9820
rect 4960 9764 5016 9820
rect 5016 9764 5020 9820
rect 4956 9760 5020 9764
rect 5036 9820 5100 9824
rect 5036 9764 5040 9820
rect 5040 9764 5096 9820
rect 5096 9764 5100 9820
rect 5036 9760 5100 9764
rect 5116 9820 5180 9824
rect 5116 9764 5120 9820
rect 5120 9764 5176 9820
rect 5176 9764 5180 9820
rect 5116 9760 5180 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 4876 8732 4940 8736
rect 4876 8676 4880 8732
rect 4880 8676 4936 8732
rect 4936 8676 4940 8732
rect 4876 8672 4940 8676
rect 4956 8732 5020 8736
rect 4956 8676 4960 8732
rect 4960 8676 5016 8732
rect 5016 8676 5020 8732
rect 4956 8672 5020 8676
rect 5036 8732 5100 8736
rect 5036 8676 5040 8732
rect 5040 8676 5096 8732
rect 5096 8676 5100 8732
rect 5036 8672 5100 8676
rect 5116 8732 5180 8736
rect 5116 8676 5120 8732
rect 5120 8676 5176 8732
rect 5176 8676 5180 8732
rect 5116 8672 5180 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 4876 7644 4940 7648
rect 4876 7588 4880 7644
rect 4880 7588 4936 7644
rect 4936 7588 4940 7644
rect 4876 7584 4940 7588
rect 4956 7644 5020 7648
rect 4956 7588 4960 7644
rect 4960 7588 5016 7644
rect 5016 7588 5020 7644
rect 4956 7584 5020 7588
rect 5036 7644 5100 7648
rect 5036 7588 5040 7644
rect 5040 7588 5096 7644
rect 5096 7588 5100 7644
rect 5036 7584 5100 7588
rect 5116 7644 5180 7648
rect 5116 7588 5120 7644
rect 5120 7588 5176 7644
rect 5176 7588 5180 7644
rect 5116 7584 5180 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 4876 6556 4940 6560
rect 4876 6500 4880 6556
rect 4880 6500 4936 6556
rect 4936 6500 4940 6556
rect 4876 6496 4940 6500
rect 4956 6556 5020 6560
rect 4956 6500 4960 6556
rect 4960 6500 5016 6556
rect 5016 6500 5020 6556
rect 4956 6496 5020 6500
rect 5036 6556 5100 6560
rect 5036 6500 5040 6556
rect 5040 6500 5096 6556
rect 5096 6500 5100 6556
rect 5036 6496 5100 6500
rect 5116 6556 5180 6560
rect 5116 6500 5120 6556
rect 5120 6500 5176 6556
rect 5176 6500 5180 6556
rect 5116 6496 5180 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 4876 5468 4940 5472
rect 4876 5412 4880 5468
rect 4880 5412 4936 5468
rect 4936 5412 4940 5468
rect 4876 5408 4940 5412
rect 4956 5468 5020 5472
rect 4956 5412 4960 5468
rect 4960 5412 5016 5468
rect 5016 5412 5020 5468
rect 4956 5408 5020 5412
rect 5036 5468 5100 5472
rect 5036 5412 5040 5468
rect 5040 5412 5096 5468
rect 5096 5412 5100 5468
rect 5036 5408 5100 5412
rect 5116 5468 5180 5472
rect 5116 5412 5120 5468
rect 5120 5412 5176 5468
rect 5176 5412 5180 5468
rect 5116 5408 5180 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 4876 4380 4940 4384
rect 4876 4324 4880 4380
rect 4880 4324 4936 4380
rect 4936 4324 4940 4380
rect 4876 4320 4940 4324
rect 4956 4380 5020 4384
rect 4956 4324 4960 4380
rect 4960 4324 5016 4380
rect 5016 4324 5020 4380
rect 4956 4320 5020 4324
rect 5036 4380 5100 4384
rect 5036 4324 5040 4380
rect 5040 4324 5096 4380
rect 5096 4324 5100 4380
rect 5036 4320 5100 4324
rect 5116 4380 5180 4384
rect 5116 4324 5120 4380
rect 5120 4324 5176 4380
rect 5176 4324 5180 4380
rect 5116 4320 5180 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 4876 3292 4940 3296
rect 4876 3236 4880 3292
rect 4880 3236 4936 3292
rect 4936 3236 4940 3292
rect 4876 3232 4940 3236
rect 4956 3292 5020 3296
rect 4956 3236 4960 3292
rect 4960 3236 5016 3292
rect 5016 3236 5020 3292
rect 4956 3232 5020 3236
rect 5036 3292 5100 3296
rect 5036 3236 5040 3292
rect 5040 3236 5096 3292
rect 5096 3236 5100 3292
rect 5036 3232 5100 3236
rect 5116 3292 5180 3296
rect 5116 3236 5120 3292
rect 5120 3236 5176 3292
rect 5176 3236 5180 3292
rect 5116 3232 5180 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 4876 2204 4940 2208
rect 4876 2148 4880 2204
rect 4880 2148 4936 2204
rect 4936 2148 4940 2204
rect 4876 2144 4940 2148
rect 4956 2204 5020 2208
rect 4956 2148 4960 2204
rect 4960 2148 5016 2204
rect 5016 2148 5020 2204
rect 4956 2144 5020 2148
rect 5036 2204 5100 2208
rect 5036 2148 5040 2204
rect 5040 2148 5096 2204
rect 5096 2148 5100 2204
rect 5036 2144 5100 2148
rect 5116 2204 5180 2208
rect 5116 2148 5120 2204
rect 5120 2148 5176 2204
rect 5176 2148 5180 2204
rect 5116 2144 5180 2148
<< metal4 >>
rect 4208 11456 4528 11472
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 4868 10912 5188 11472
rect 4868 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5188 10912
rect 4868 9824 5188 10848
rect 4868 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5188 9824
rect 4868 8736 5188 9760
rect 4868 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5188 8736
rect 4868 7648 5188 8672
rect 4868 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5188 7648
rect 4868 6560 5188 7584
rect 4868 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5188 6560
rect 4868 5472 5188 6496
rect 4868 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5188 5472
rect 4868 4384 5188 5408
rect 4868 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5188 4384
rect 4868 3296 5188 4320
rect 4868 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5188 3296
rect 4868 2208 5188 3232
rect 4868 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5188 2208
rect 4868 2128 5188 2144
use sky130_fd_sc_hd__inv_2  _050_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform 1 0 2024 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _051_
timestamp 1707688321
transform 1 0 1840 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and4bb_1  _052_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform -1 0 7268 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__and3b_1  _053_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform -1 0 6992 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _054_
timestamp 1707688321
transform -1 0 7728 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _055_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform -1 0 5152 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_1  _056_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform -1 0 7820 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _057_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform 1 0 1472 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _058_
timestamp 1707688321
transform -1 0 5612 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or4bb_1  _059_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform 1 0 3680 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _060_
timestamp 1707688321
transform -1 0 4048 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  _061_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform -1 0 6164 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__nor3b_1  _062_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform 1 0 3680 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__nor3b_1  _063_
timestamp 1707688321
transform 1 0 4784 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _064_
timestamp 1707688321
transform 1 0 6348 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__nor3b_1  _065_
timestamp 1707688321
transform -1 0 4784 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _066_
timestamp 1707688321
transform 1 0 5612 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _067_
timestamp 1707688321
transform 1 0 5612 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _068_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform -1 0 5796 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _069_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform -1 0 2116 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_2  _070_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform 1 0 5796 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _071_
timestamp 1707688321
transform -1 0 6256 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _072_
timestamp 1707688321
transform -1 0 4416 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__o21bai_1  _073_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform 1 0 4508 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a211oi_1  _074_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform -1 0 4324 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _075_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform -1 0 5520 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _076_
timestamp 1707688321
transform 1 0 6992 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o21bai_1  _077_
timestamp 1707688321
transform 1 0 5152 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _078_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform 1 0 6624 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__o311a_1  _079_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform 1 0 6348 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _080_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform -1 0 8004 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _081_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform -1 0 8648 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _082_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform -1 0 8280 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _083_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform 1 0 6808 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _084_
timestamp 1707688321
transform 1 0 5152 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _085_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform 1 0 6532 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__o211a_1  _086_
timestamp 1707688321
transform -1 0 7084 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _087_
timestamp 1707688321
transform 1 0 8924 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o2bb2a_1  _088_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform -1 0 9292 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _089_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform -1 0 8464 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _090_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform -1 0 8740 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _091_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform 1 0 7360 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__and4_1  _092_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform -1 0 8096 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _093_
timestamp 1707688321
transform -1 0 8740 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _094_
timestamp 1707688321
transform 1 0 5612 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_1  _095_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform 1 0 6716 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _096_
timestamp 1707688321
transform -1 0 6624 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o32a_1  _097_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform 1 0 4784 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _098_
timestamp 1707688321
transform -1 0 5704 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _099_
timestamp 1707688321
transform 1 0 5612 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _100_
timestamp 1707688321
transform -1 0 5980 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o2bb2a_1  _101_
timestamp 1707688321
transform 1 0 4784 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _102_
timestamp 1707688321
transform 1 0 3864 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _103_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform 1 0 4692 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _104_
timestamp 1707688321
transform -1 0 3680 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a41o_1  _105_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform 1 0 3772 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _106_
timestamp 1707688321
transform -1 0 5152 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o21ba_1  _107_
timestamp 1707688321
transform 1 0 2944 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _108_
timestamp 1707688321
transform -1 0 2300 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _109_
timestamp 1707688321
transform -1 0 2944 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a41o_1  _110_
timestamp 1707688321
transform 1 0 2668 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _111_
timestamp 1707688321
transform 1 0 2392 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _112_
timestamp 1707688321
transform -1 0 2392 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__dfrtp_1  _113_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform 1 0 2576 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _114_
timestamp 1707688321
transform 1 0 3772 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _115_
timestamp 1707688321
transform 1 0 4416 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _116_
timestamp 1707688321
transform -1 0 6992 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _117_
timestamp 1707688321
transform -1 0 8832 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _118_
timestamp 1707688321
transform -1 0 8924 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _119_
timestamp 1707688321
transform 1 0 6164 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _120_
timestamp 1707688321
transform -1 0 8556 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _121_
timestamp 1707688321
transform 1 0 6348 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _122_
timestamp 1707688321
transform 1 0 6624 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _123_
timestamp 1707688321
transform 1 0 4416 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _124_
timestamp 1707688321
transform 1 0 4140 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _125_
timestamp 1707688321
transform 1 0 2300 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _126_
timestamp 1707688321
transform 1 0 2852 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _127_
timestamp 1707688321
transform 1 0 1380 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _128_
timestamp 1707688321
transform -1 0 3220 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _129_
timestamp 1707688321
transform 1 0 1840 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _130_
timestamp 1707688321
transform 1 0 1380 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__conb_1  _130__27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform 1 0 1748 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _131_
timestamp 1707688321
transform 1 0 1380 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_osc_ck $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform 1 0 4784 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_osc_ck
timestamp 1707688321
transform -1 0 4416 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_osc_ck
timestamp 1707688321
transform 1 0 7728 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_2  fanout22 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform -1 0 3680 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout23
timestamp 1707688321
transform 1 0 7820 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout24 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform -1 0 4600 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout25
timestamp 1707688321
transform 1 0 5612 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout26 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform -1 0 6716 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_15 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform 1 0 2484 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_39
timestamp 1707688321
transform 1 0 4692 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_57
timestamp 1707688321
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_63 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform 1 0 6900 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_70
timestamp 1707688321
transform 1 0 7544 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_77
timestamp 1707688321
transform 1 0 8188 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_85
timestamp 1707688321
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_97
timestamp 1707688321
transform 1 0 10028 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1707688321
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1707688321
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_27
timestamp 1707688321
transform 1 0 3588 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_46
timestamp 1707688321
transform 1 0 5336 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_64
timestamp 1707688321
transform 1 0 6992 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_76
timestamp 1707688321
transform 1 0 8096 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_88 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform 1 0 9200 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_96
timestamp 1707688321
transform 1 0 9936 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_6
timestamp 1707688321
transform 1 0 1656 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_18
timestamp 1707688321
transform 1 0 2760 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_26
timestamp 1707688321
transform 1 0 3496 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_29
timestamp 1707688321
transform 1 0 3772 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_35
timestamp 1707688321
transform 1 0 4324 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_42 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform 1 0 4968 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_55
timestamp 1707688321
transform 1 0 6164 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_67
timestamp 1707688321
transform 1 0 7268 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_79
timestamp 1707688321
transform 1 0 8372 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 1707688321
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_85
timestamp 1707688321
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_97
timestamp 1707688321
transform 1 0 10028 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_13
timestamp 1707688321
transform 1 0 2300 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_25 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform 1 0 3404 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_31
timestamp 1707688321
transform 1 0 3956 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_38
timestamp 1707688321
transform 1 0 4600 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_48
timestamp 1707688321
transform 1 0 5520 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_53
timestamp 1707688321
transform 1 0 5980 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_57
timestamp 1707688321
transform 1 0 6348 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_61
timestamp 1707688321
transform 1 0 6716 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp 1707688321
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_81
timestamp 1707688321
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_93
timestamp 1707688321
transform 1 0 9660 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_23
timestamp 1707688321
transform 1 0 3220 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1707688321
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_50
timestamp 1707688321
transform 1 0 5704 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_64
timestamp 1707688321
transform 1 0 6992 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_77
timestamp 1707688321
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 1707688321
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_85
timestamp 1707688321
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_97
timestamp 1707688321
transform 1 0 10028 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_6
timestamp 1707688321
transform 1 0 1656 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_14
timestamp 1707688321
transform 1 0 2392 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_85
timestamp 1707688321
transform 1 0 8924 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_97
timestamp 1707688321
transform 1 0 10028 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1707688321
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_43
timestamp 1707688321
transform 1 0 5060 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_85
timestamp 1707688321
transform 1 0 8924 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_93
timestamp 1707688321
transform 1 0 9660 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_3
timestamp 1707688321
transform 1 0 1380 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_44
timestamp 1707688321
transform 1 0 5152 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_53
timestamp 1707688321
transform 1 0 5980 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_78
timestamp 1707688321
transform 1 0 8280 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_90
timestamp 1707688321
transform 1 0 9384 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_98
timestamp 1707688321
transform 1 0 10120 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1707688321
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_82
timestamp 1707688321
transform 1 0 8648 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_90
timestamp 1707688321
transform 1 0 9384 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_98
timestamp 1707688321
transform 1 0 10120 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_7
timestamp 1707688321
transform 1 0 1748 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_92
timestamp 1707688321
transform 1 0 9568 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_98
timestamp 1707688321
transform 1 0 10120 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_80
timestamp 1707688321
transform 1 0 8464 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_93
timestamp 1707688321
transform 1 0 9660 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_3
timestamp 1707688321
transform 1 0 1380 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_25
timestamp 1707688321
transform 1 0 3404 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_37
timestamp 1707688321
transform 1 0 4508 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_60
timestamp 1707688321
transform 1 0 6624 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_89
timestamp 1707688321
transform 1 0 9292 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_97
timestamp 1707688321
transform 1 0 10028 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_23
timestamp 1707688321
transform 1 0 3220 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_56
timestamp 1707688321
transform 1 0 6256 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_73
timestamp 1707688321
transform 1 0 7820 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_82
timestamp 1707688321
transform 1 0 8648 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_85
timestamp 1707688321
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_97
timestamp 1707688321
transform 1 0 10028 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_3
timestamp 1707688321
transform 1 0 1380 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_20
timestamp 1707688321
transform 1 0 2944 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_28
timestamp 1707688321
transform 1 0 3680 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_43
timestamp 1707688321
transform 1 0 5060 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_54
timestamp 1707688321
transform 1 0 6072 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_57
timestamp 1707688321
transform 1 0 6348 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_83
timestamp 1707688321
transform 1 0 8740 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_95
timestamp 1707688321
transform 1 0 9844 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_3
timestamp 1707688321
transform 1 0 1380 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_7
timestamp 1707688321
transform 1 0 1748 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_37
timestamp 1707688321
transform 1 0 4508 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_53
timestamp 1707688321
transform 1 0 5980 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_83
timestamp 1707688321
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_85
timestamp 1707688321
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_97
timestamp 1707688321
transform 1 0 10028 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_3
timestamp 1707688321
transform 1 0 1380 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_11
timestamp 1707688321
transform 1 0 2116 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_85
timestamp 1707688321
transform 1 0 8924 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_97
timestamp 1707688321
transform 1 0 10028 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_3
timestamp 1707688321
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_15
timestamp 1707688321
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_27
timestamp 1707688321
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_29
timestamp 1707688321
transform 1 0 3772 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_37
timestamp 1707688321
transform 1 0 4508 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_50
timestamp 1707688321
transform 1 0 5704 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_65
timestamp 1707688321
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_77
timestamp 1707688321
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_83
timestamp 1707688321
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_85
timestamp 1707688321
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_97
timestamp 1707688321
transform 1 0 10028 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform 1 0 4416 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1707688321
transform -1 0 2852 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1707688321
transform -1 0 7820 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1707688321
transform -1 0 4508 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1707688321
transform -1 0 2576 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1707688321
transform -1 0 9660 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1707688321
transform -1 0 6256 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 1707688321
transform -1 0 5980 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 1707688321
transform -1 0 5060 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 1707688321
transform -1 0 7084 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 1707688321
transform 1 0 7912 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp 1707688321
transform -1 0 4784 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 1707688321
transform -1 0 8924 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold14
timestamp 1707688321
transform -1 0 6624 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold15
timestamp 1707688321
transform 1 0 1932 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform -1 0 1656 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1707688321
transform -1 0 1656 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1707688321
transform -1 0 1656 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input4 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform -1 0 10212 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input5 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform 1 0 9108 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input6
timestamp 1707688321
transform 1 0 2668 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input7
timestamp 1707688321
transform 1 0 3772 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input8
timestamp 1707688321
transform 1 0 2116 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output9
timestamp 1707688321
transform -1 0 1748 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output10
timestamp 1707688321
transform 1 0 3220 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output11
timestamp 1707688321
transform 1 0 6532 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output12
timestamp 1707688321
transform 1 0 3956 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output13
timestamp 1707688321
transform 1 0 4876 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output14
timestamp 1707688321
transform 1 0 7176 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output15
timestamp 1707688321
transform 1 0 4600 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output16
timestamp 1707688321
transform 1 0 7820 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output17
timestamp 1707688321
transform 1 0 8464 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output18
timestamp 1707688321
transform 1 0 5244 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output19
timestamp 1707688321
transform -1 0 3588 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output20
timestamp 1707688321
transform -1 0 6256 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output21
timestamp 1707688321
transform -1 0 1748 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_17
timestamp 1707688321
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1707688321
transform -1 0 10488 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_18
timestamp 1707688321
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1707688321
transform -1 0 10488 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_19
timestamp 1707688321
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1707688321
transform -1 0 10488 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_20
timestamp 1707688321
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1707688321
transform -1 0 10488 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_21
timestamp 1707688321
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1707688321
transform -1 0 10488 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_22
timestamp 1707688321
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1707688321
transform -1 0 10488 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_23
timestamp 1707688321
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1707688321
transform -1 0 10488 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_24
timestamp 1707688321
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1707688321
transform -1 0 10488 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_25
timestamp 1707688321
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1707688321
transform -1 0 10488 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_26
timestamp 1707688321
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1707688321
transform -1 0 10488 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_27
timestamp 1707688321
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 1707688321
transform -1 0 10488 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_28
timestamp 1707688321
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 1707688321
transform -1 0 10488 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_29
timestamp 1707688321
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 1707688321
transform -1 0 10488 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_30
timestamp 1707688321
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 1707688321
transform -1 0 10488 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_31
timestamp 1707688321
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 1707688321
transform -1 0 10488 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_32
timestamp 1707688321
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 1707688321
transform -1 0 10488 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_33
timestamp 1707688321
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 1707688321
transform -1 0 10488 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_34 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_35
timestamp 1707688321
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_36
timestamp 1707688321
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_37
timestamp 1707688321
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_38
timestamp 1707688321
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_39
timestamp 1707688321
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_40
timestamp 1707688321
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_41
timestamp 1707688321
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_42
timestamp 1707688321
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_43
timestamp 1707688321
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_44
timestamp 1707688321
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_45
timestamp 1707688321
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_46
timestamp 1707688321
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_47
timestamp 1707688321
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_48
timestamp 1707688321
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_49
timestamp 1707688321
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_50
timestamp 1707688321
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_51
timestamp 1707688321
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_52
timestamp 1707688321
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_53
timestamp 1707688321
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_54
timestamp 1707688321
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_55
timestamp 1707688321
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_56
timestamp 1707688321
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_57
timestamp 1707688321
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_58
timestamp 1707688321
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_59
timestamp 1707688321
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_60
timestamp 1707688321
transform 1 0 6256 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_61
timestamp 1707688321
transform 1 0 8832 0 1 10880
box -38 -48 130 592
<< labels >>
flabel metal4 s 4868 2128 5188 11472 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 4208 2128 4528 11472 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 0 5448 800 5568 0 FreeSans 480 0 0 0 force_dis_rc_osc
port 2 nsew signal input
flabel metal3 s 0 7488 800 7608 0 FreeSans 480 0 0 0 force_ena_rc_osc
port 3 nsew signal input
flabel metal3 s 0 3408 800 3528 0 FreeSans 480 0 0 0 force_pdn
port 4 nsew signal input
flabel metal3 s 0 4088 800 4208 0 FreeSans 480 0 0 0 force_pdnb
port 5 nsew signal output
flabel metal3 s 10793 5448 11593 5568 0 FreeSans 480 0 0 0 force_short_oneshot
port 6 nsew signal input
flabel metal3 s 0 10208 800 10328 0 FreeSans 480 0 0 0 osc_ck
port 7 nsew signal input
flabel metal3 s 0 6128 800 6248 0 FreeSans 480 0 0 0 osc_ena
port 8 nsew signal output
flabel metal2 s 9034 0 9090 800 0 FreeSans 224 90 0 0 otrip[0]
port 9 nsew signal input
flabel metal2 s 2594 0 2650 800 0 FreeSans 224 90 0 0 otrip[1]
port 10 nsew signal input
flabel metal2 s 3238 0 3294 800 0 FreeSans 224 90 0 0 otrip[2]
port 11 nsew signal input
flabel metal2 s 6458 0 6514 800 0 FreeSans 224 90 0 0 otrip_decoded[0]
port 12 nsew signal output
flabel metal2 s 3882 0 3938 800 0 FreeSans 224 90 0 0 otrip_decoded[1]
port 13 nsew signal output
flabel metal2 s 5170 0 5226 800 0 FreeSans 224 90 0 0 otrip_decoded[2]
port 14 nsew signal output
flabel metal2 s 7102 0 7158 800 0 FreeSans 224 90 0 0 otrip_decoded[3]
port 15 nsew signal output
flabel metal2 s 4526 0 4582 800 0 FreeSans 224 90 0 0 otrip_decoded[4]
port 16 nsew signal output
flabel metal2 s 7746 0 7802 800 0 FreeSans 224 90 0 0 otrip_decoded[5]
port 17 nsew signal output
flabel metal2 s 8390 0 8446 800 0 FreeSans 224 90 0 0 otrip_decoded[6]
port 18 nsew signal output
flabel metal2 s 5814 0 5870 800 0 FreeSans 224 90 0 0 otrip_decoded[7]
port 19 nsew signal output
flabel metal3 s 0 6808 800 6928 0 FreeSans 480 0 0 0 por_timed_out
port 20 nsew signal output
flabel metal2 s 5814 12937 5870 13737 0 FreeSans 224 90 0 0 por_unbuf
port 21 nsew signal output
flabel metal3 s 0 4768 800 4888 0 FreeSans 480 0 0 0 pwup_filt
port 22 nsew signal input
flabel metal3 s 0 8168 800 8288 0 FreeSans 480 0 0 0 startup_timed_out
port 23 nsew signal output
rlabel metal1 5796 10880 5796 10880 0 VGND
rlabel metal1 5796 11424 5796 11424 0 VPWR
rlabel metal1 3588 4794 3588 4794 0 _000_
rlabel metal1 4370 5746 4370 5746 0 _001_
rlabel metal1 5106 4794 5106 4794 0 _002_
rlabel metal1 6532 5338 6532 5338 0 _003_
rlabel metal1 8470 5882 8470 5882 0 _004_
rlabel metal1 8004 4046 8004 4046 0 _005_
rlabel metal1 6532 9690 6532 9690 0 _006_
rlabel metal1 8372 8398 8372 8398 0 _007_
rlabel metal2 7406 10132 7406 10132 0 _008_
rlabel metal1 6854 7514 6854 7514 0 _009_
rlabel metal2 4738 7854 4738 7854 0 _010_
rlabel metal2 4830 10404 4830 10404 0 _011_
rlabel metal1 4186 10540 4186 10540 0 _012_
rlabel metal1 3174 6392 3174 6392 0 _013_
rlabel via1 1695 6970 1695 6970 0 _014_
rlabel via1 2904 9146 2904 9146 0 _015_
rlabel metal2 1794 9724 1794 9724 0 _016_
rlabel metal2 5658 7718 5658 7718 0 _017_
rlabel metal1 5198 8364 5198 8364 0 _018_
rlabel metal1 5704 10030 5704 10030 0 _019_
rlabel metal1 4002 9554 4002 9554 0 _020_
rlabel metal1 5290 9894 5290 9894 0 _021_
rlabel metal1 4600 9486 4600 9486 0 _022_
rlabel metal1 3358 7854 3358 7854 0 _023_
rlabel metal2 3818 7888 3818 7888 0 _024_
rlabel metal1 3174 7888 3174 7888 0 _025_
rlabel metal1 2300 9486 2300 9486 0 _026_
rlabel metal2 2714 9010 2714 9010 0 _027_
rlabel metal1 1886 5338 1886 5338 0 _028_
rlabel metal1 6486 6426 6486 6426 0 _029_
rlabel metal1 7038 5270 7038 5270 0 _030_
rlabel metal1 4370 8466 4370 8466 0 _031_
rlabel metal1 4324 8262 4324 8262 0 _032_
rlabel metal2 2714 8092 2714 8092 0 _033_
rlabel via2 5198 9571 5198 9571 0 _034_
rlabel metal1 4554 8602 4554 8602 0 _035_
rlabel metal1 6026 10642 6026 10642 0 _036_
rlabel metal1 3818 5678 3818 5678 0 _037_
rlabel metal1 5612 4590 5612 4590 0 _038_
rlabel metal1 6118 4726 6118 4726 0 _039_
rlabel metal1 6854 5134 6854 5134 0 _040_
rlabel metal1 7636 6086 7636 6086 0 _041_
rlabel metal1 8188 6290 8188 6290 0 _042_
rlabel metal2 8878 8908 8878 8908 0 _043_
rlabel metal1 8694 8398 8694 8398 0 _044_
rlabel metal1 8510 6698 8510 6698 0 _045_
rlabel metal2 7682 9860 7682 9860 0 _046_
rlabel metal1 8418 9894 8418 9894 0 _047_
rlabel metal1 7406 6970 7406 6970 0 _048_
rlabel metal1 5612 9690 5612 9690 0 _049_
rlabel metal1 5244 7718 5244 7718 0 clknet_0_osc_ck
rlabel metal1 2346 10710 2346 10710 0 clknet_1_0__leaf_osc_ck
rlabel metal1 6256 10098 6256 10098 0 clknet_1_1__leaf_osc_ck
rlabel metal1 8832 9554 8832 9554 0 cnt_por\[0\]
rlabel metal2 4462 9860 4462 9860 0 cnt_por\[10\]
rlabel metal1 8740 9418 8740 9418 0 cnt_por\[1\]
rlabel metal1 8188 9962 8188 9962 0 cnt_por\[2\]
rlabel metal1 8970 7990 8970 7990 0 cnt_por\[3\]
rlabel metal2 5474 10355 5474 10355 0 cnt_por\[4\]
rlabel metal1 6302 11050 6302 11050 0 cnt_por\[5\]
rlabel metal1 4186 10438 4186 10438 0 cnt_por\[6\]
rlabel metal2 4646 7582 4646 7582 0 cnt_por\[7\]
rlabel metal2 2438 7888 2438 7888 0 cnt_por\[8\]
rlabel metal1 1472 8466 1472 8466 0 cnt_por\[9\]
rlabel metal1 4600 4658 4600 4658 0 cnt_rsb
rlabel metal2 3174 5508 3174 5508 0 cnt_rsb_stg1
rlabel metal1 6118 6630 6118 6630 0 cnt_st\[0\]
rlabel metal1 5474 6970 5474 6970 0 cnt_st\[1\]
rlabel metal1 6900 6290 6900 6290 0 cnt_st\[2\]
rlabel metal1 6440 5202 6440 5202 0 cnt_st\[3\]
rlabel metal2 7314 6528 7314 6528 0 cnt_st\[4\]
rlabel metal1 7038 5134 7038 5134 0 cnt_st\[5\]
rlabel metal3 1050 5508 1050 5508 0 force_dis_rc_osc
rlabel metal3 1050 7548 1050 7548 0 force_ena_rc_osc
rlabel metal3 751 3468 751 3468 0 force_pdn
rlabel metal3 1096 4148 1096 4148 0 force_pdnb
rlabel metal1 10166 5644 10166 5644 0 force_short_oneshot
rlabel metal1 1748 5202 1748 5202 0 net1
rlabel metal2 2070 5984 2070 5984 0 net10
rlabel metal1 6348 2414 6348 2414 0 net11
rlabel metal1 3864 3162 3864 3162 0 net12
rlabel metal1 4876 2414 4876 2414 0 net13
rlabel metal1 7084 2414 7084 2414 0 net14
rlabel metal1 4692 3162 4692 3162 0 net15
rlabel metal1 7590 2414 7590 2414 0 net16
rlabel metal1 8510 2380 8510 2380 0 net17
rlabel metal1 5336 2414 5336 2414 0 net18
rlabel metal1 3634 6766 3634 6766 0 net19
rlabel metal2 1610 7004 1610 7004 0 net2
rlabel metal2 6118 10336 6118 10336 0 net20
rlabel metal2 7866 5610 7866 5610 0 net21
rlabel metal1 5060 6086 5060 6086 0 net22
rlabel metal1 2231 7378 2231 7378 0 net23
rlabel metal1 6079 7378 6079 7378 0 net24
rlabel metal2 7222 9622 7222 9622 0 net25
rlabel metal1 5198 4556 5198 4556 0 net26
rlabel metal1 1748 4250 1748 4250 0 net27
rlabel metal1 4784 4454 4784 4454 0 net28
rlabel metal1 1787 5882 1787 5882 0 net29
rlabel metal1 1840 3706 1840 3706 0 net3
rlabel metal1 7084 4114 7084 4114 0 net30
rlabel metal1 2461 9554 2461 9554 0 net31
rlabel metal1 1978 7514 1978 7514 0 net32
rlabel metal1 7406 7344 7406 7344 0 net33
rlabel metal1 5428 8398 5428 8398 0 net34
rlabel metal1 4784 5678 4784 5678 0 net35
rlabel metal1 4508 5882 4508 5882 0 net36
rlabel metal1 5704 10098 5704 10098 0 net37
rlabel metal1 8648 8466 8648 8466 0 net38
rlabel metal1 3634 7820 3634 7820 0 net39
rlabel metal1 6716 7378 6716 7378 0 net4
rlabel metal1 8050 9520 8050 9520 0 net40
rlabel metal1 5704 4182 5704 4182 0 net41
rlabel metal1 2760 8398 2760 8398 0 net42
rlabel metal1 8096 3094 8096 3094 0 net5
rlabel metal1 3450 2958 3450 2958 0 net6
rlabel metal2 4002 2720 4002 2720 0 net7
rlabel metal2 2346 4760 2346 4760 0 net8
rlabel metal1 1702 4080 1702 4080 0 net9
rlabel metal3 1717 10268 1717 10268 0 osc_ck
rlabel metal2 3450 6035 3450 6035 0 osc_ena
rlabel metal2 9062 1027 9062 1027 0 otrip[0]
rlabel metal2 2622 1588 2622 1588 0 otrip[1]
rlabel metal2 3266 1588 3266 1588 0 otrip[2]
rlabel metal2 6486 1520 6486 1520 0 otrip_decoded[0]
rlabel metal1 4048 3366 4048 3366 0 otrip_decoded[1]
rlabel metal2 5198 959 5198 959 0 otrip_decoded[2]
rlabel metal2 7130 1520 7130 1520 0 otrip_decoded[3]
rlabel metal2 4554 1231 4554 1231 0 otrip_decoded[4]
rlabel metal2 7774 1520 7774 1520 0 otrip_decoded[5]
rlabel metal2 8418 1520 8418 1520 0 otrip_decoded[6]
rlabel metal2 5842 1520 5842 1520 0 otrip_decoded[7]
rlabel metal2 3358 6749 3358 6749 0 por_timed_out
rlabel metal1 5934 11322 5934 11322 0 por_unbuf
rlabel metal3 912 4828 912 4828 0 pwup_filt
rlabel metal1 1334 7514 1334 7514 0 startup_timed_out
<< properties >>
string FIXED_BBOX 0 0 11593 13737
<< end >>
