../../por_dig.out.spice