magic
tech sky130A
magscale 1 2
timestamp 1712973328
<< pwell >>
rect -1182 40391 42901 40527
rect -1182 -559 -1046 40391
rect 42765 -559 42901 40391
rect -1182 -695 42901 -559
<< psubdiff >>
rect -1146 40457 -1086 40491
rect 42805 40457 42865 40491
rect -1146 40431 -1112 40457
rect -1146 -625 -1112 -599
rect 42831 40431 42865 40457
rect 42831 -625 42865 -599
rect -1146 -659 -1086 -625
rect 42805 -659 42865 -625
<< psubdiffcont >>
rect -1086 40457 42805 40491
rect -1146 -599 -1112 40431
rect 42831 -599 42865 40431
rect -1086 -659 42805 -625
<< locali >>
rect -1146 40457 -1086 40491
rect 42805 40457 42865 40491
rect -1146 40431 -1112 40457
rect -1146 -625 -1112 -599
rect 42831 40431 42865 40457
rect 42831 -625 42865 -599
rect -1146 -659 -1086 -625
rect 42805 -659 42865 -625
<< viali >>
rect -1086 40457 42805 40491
rect -1146 -556 -1112 40404
rect 42831 -567 42865 40393
rect -1086 -659 42805 -625
<< metal1 >>
rect 41177 40601 41325 40612
rect 41177 40531 41188 40601
rect -1186 40491 41188 40531
rect 41314 40531 41325 40601
rect 41314 40491 42905 40531
rect -1186 40457 -1086 40491
rect 42805 40457 42905 40491
rect -1186 40404 42905 40457
rect -1186 -556 -1146 40404
rect -1112 40393 42905 40404
rect -1112 40391 42831 40393
rect -1112 -556 -1046 40391
rect 42223 27573 42301 27619
rect 42255 27563 42301 27573
rect 42067 27404 42131 27468
rect 42255 27303 42301 27471
rect 42223 27257 42301 27303
rect 42134 27088 42198 27152
rect 42255 26987 42301 27257
rect 42223 26941 42301 26987
rect 42024 26763 42088 26827
rect 42255 26671 42301 26941
rect 42223 26625 42301 26671
rect 42084 26451 42158 26525
rect 42255 26355 42301 26625
rect 42223 26309 42301 26355
rect 42104 26133 42178 26207
rect 42255 26039 42301 26309
rect 42223 25993 42301 26039
rect 42096 25819 42170 25893
rect 42255 25723 42301 25993
rect 42223 25677 42301 25723
rect 42134 25505 42198 25569
rect 42255 25407 42301 25677
rect 42223 25388 42301 25407
rect 42765 25388 42831 40391
rect 42223 25361 42831 25388
rect 42255 25281 42831 25361
rect 42036 25189 42100 25253
rect 42255 25193 42301 25281
rect 42255 25091 42301 25119
rect 42223 25045 42301 25091
rect -1186 -559 -1046 -556
rect 42765 -559 42831 25281
rect -1186 -567 42831 -559
rect 42865 -567 42905 40393
rect -1186 -625 42905 -567
rect -1186 -659 -1086 -625
rect 42805 -659 42905 -625
rect -1186 -699 42905 -659
<< via1 >>
rect 41188 40491 41314 40601
rect 41188 40475 41314 40491
<< metal2 >>
rect 41177 40603 41325 40612
rect 41177 40473 41186 40603
rect 41316 40473 41325 40603
rect 41177 40464 41325 40473
rect 1111 40272 1507 40292
rect 1111 39982 1131 40272
rect 1471 39982 1507 40272
rect 1111 39265 1507 39982
rect 1577 39865 1962 39896
rect 1577 39606 1599 39865
rect 1934 39606 1962 39865
rect 1577 39251 1962 39606
rect 10 -707 396 1690
rect 493 -110 893 1899
rect 493 -519 893 -510
rect 10 -1039 28 -707
rect 383 -1039 396 -707
rect 10 -1056 396 -1039
<< via2 >>
rect 41186 40601 41316 40603
rect 41186 40475 41188 40601
rect 41188 40475 41314 40601
rect 41314 40475 41316 40601
rect 41186 40473 41316 40475
rect 1131 39982 1471 40272
rect 1599 39606 1934 39865
rect 493 -510 893 -110
rect 28 -1039 383 -707
<< metal3 >>
rect -1604 41276 43293 41282
rect -1604 40888 -1598 41276
rect -1210 40888 42899 41276
rect 43287 40888 43293 41276
rect -1604 40882 43293 40888
rect -1604 40816 43293 40822
rect -1604 40428 -1138 40816
rect -750 40603 42439 40816
rect -750 40473 41186 40603
rect 41316 40473 42439 40603
rect -750 40428 42439 40473
rect 42827 40428 43293 40816
rect -1604 40422 43293 40428
rect -1604 40356 43293 40362
rect -1604 39968 -678 40356
rect -290 40272 41979 40356
rect -290 39982 1131 40272
rect 1471 39982 41979 40272
rect -290 39968 41979 39982
rect 42367 39968 43293 40356
rect -1604 39962 43293 39968
rect -1604 39896 43293 39902
rect -1604 39508 -218 39896
rect 170 39865 41519 39896
rect 170 39606 1599 39865
rect 1934 39606 41519 39865
rect 170 39508 41519 39606
rect 41907 39508 43293 39896
rect -1604 39502 43293 39508
rect 947 39492 1357 39502
rect 488 -110 898 -105
rect 488 -207 493 -110
rect -1604 -213 493 -207
rect -1604 -601 -218 -213
rect 170 -510 493 -213
rect 893 -207 898 -110
rect 893 -213 43293 -207
rect 893 -510 41519 -213
rect 170 -601 41519 -510
rect 41907 -601 43293 -213
rect -1604 -607 43293 -601
rect -1604 -673 43293 -667
rect -1604 -1061 -678 -673
rect -290 -707 41979 -673
rect -290 -1039 28 -707
rect 383 -1039 41979 -707
rect -290 -1061 41979 -1039
rect 42367 -1061 43293 -673
rect -1604 -1067 43293 -1061
rect -1604 -1133 43293 -1127
rect -1604 -1521 -1138 -1133
rect -750 -1521 42439 -1133
rect 42827 -1521 43293 -1133
rect -1604 -1527 43293 -1521
rect -1604 -1593 43293 -1587
rect -1604 -1981 -1598 -1593
rect -1210 -1981 42899 -1593
rect 43287 -1981 43293 -1593
rect -1604 -1987 43293 -1981
<< via3 >>
rect -1598 40888 -1210 41276
rect 42899 40888 43287 41276
rect -1138 40428 -750 40816
rect 42439 40428 42827 40816
rect -678 39968 -290 40356
rect 41979 39968 42367 40356
rect -218 39508 170 39896
rect 41519 39508 41907 39896
rect -218 -601 170 -213
rect 41519 -601 41907 -213
rect -678 -1061 -290 -673
rect 41979 -1061 42367 -673
rect -1138 -1521 -750 -1133
rect 42439 -1521 42827 -1133
rect -1598 -1981 -1210 -1593
rect 42899 -1981 43287 -1593
<< metal4 >>
rect -1604 41276 -1204 41283
rect -1604 40888 -1598 41276
rect -1210 40888 -1204 41276
rect -1604 -1593 -1204 40888
rect -1604 -1981 -1598 -1593
rect -1210 -1981 -1204 -1593
rect -1604 -1987 -1204 -1981
rect -1144 40816 -744 41283
rect -1144 40428 -1138 40816
rect -750 40428 -744 40816
rect -1144 -1133 -744 40428
rect -1144 -1521 -1138 -1133
rect -750 -1521 -744 -1133
rect -1144 -1987 -744 -1521
rect -684 40356 -284 41283
rect -684 39968 -678 40356
rect -290 39968 -284 40356
rect -684 -673 -284 39968
rect -684 -1061 -678 -673
rect -290 -1061 -284 -673
rect -684 -1987 -284 -1061
rect -224 39896 176 41283
rect -224 39508 -218 39896
rect 170 39508 176 39896
rect -224 7639 176 39508
rect 41513 39896 41913 41283
rect 41513 39508 41519 39896
rect 41907 39508 41913 39896
rect -224 7237 180 7639
rect -224 -213 176 7237
rect -224 -601 -218 -213
rect 170 -601 176 -213
rect -224 -1987 176 -601
rect 41513 -213 41913 39508
rect 41513 -601 41519 -213
rect 41907 -601 41913 -213
rect 41513 -1987 41913 -601
rect 41973 40356 42373 41283
rect 41973 39968 41979 40356
rect 42367 39968 42373 40356
rect 41973 -673 42373 39968
rect 41973 -1061 41979 -673
rect 42367 -1061 42373 -673
rect 41973 -1987 42373 -1061
rect 42433 40816 42833 41283
rect 42433 40428 42439 40816
rect 42827 40428 42833 40816
rect 42433 -1133 42833 40428
rect 42433 -1521 42439 -1133
rect 42827 -1521 42833 -1133
rect 42433 -1987 42833 -1521
rect 42893 41276 43293 41283
rect 42893 40888 42899 41276
rect 43287 40888 43293 41276
rect 42893 -1593 43293 40888
rect 42893 -1981 42899 -1593
rect 43287 -1981 43293 -1593
rect 42893 -1987 43293 -1981
use sky130_fd_pr__nfet_g5v0d10v5_PXF6AN  sky130_fd_pr__nfet_g5v0d10v5_PXF6AN_0
timestamp 1712947988
transform 0 1 42123 -1 0 26332
box -1463 -358 1463 358
<< labels >>
flabel metal3 1723 -1527 1723 -1527 0 FreeSans 1600 0 0 0 dvss
port 6 nsew
flabel metal3 1723 -1987 1723 -1987 0 FreeSans 1600 0 0 0 dvdd
port 4 nsew
flabel metal3 1723 -607 1723 -607 0 FreeSans 1600 0 0 0 avss
port 2 nsew
flabel metal3 1723 -1067 1723 -1067 0 FreeSans 1600 0 0 0 avdd
port 1 nsew
<< end >>
