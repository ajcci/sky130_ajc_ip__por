** sch_path: /home/rtsang/chipalooza/sky130_ajc_ip__por/xschem/tb_por.sch
**.subckt tb_por
Vavss avss GND 0
Vena force_pdn GND pwl (0 0 500u 0 500.01u dvdd 600u dvdd 600.01u 0)
Vavdd avdd GND pwl (0 0 20u 0 400u avdd 700u avdd 900u 2 1000u 2 1200u avdd)
.save i(vavdd)
Vbg vbg_1v2 GND 1.2
Ibias vbp avss 200n
XM1 ibg_200n vbp avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM0 vbp vbp avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
Vdvss dvss GND 0
Vdvdd dvdd GND dvdd
.save i(vdvdd)
R1 itest GND 1e6 m=1
C1 porb_h GND 20p m=1
C2 porb GND 20p m=1
C3 por GND 20p m=1
xIpor porb_h avdd avss porb dvdd por dvss osc_ck vbg_1v2 osc_ck_256 otrip_2_ otrip_1_ otrip_0_ itest pwup_filt force_pdn vin
+ force_rc_osc force_short_oneshot startup_timed_out por_timed_out isrc_sel ibg_200n por
Vvotrip0 otrip_0_ GND DC 0
.save i(vvotrip0)
Vvotrip1 otrip_1_ GND DC 0
.save i(vvotrip1)
Vvotrip2 otrip_2_ GND DC 0
.save i(vvotrip2)
**** begin user architecture code


.param avdd=3.3
.param dvdd=1.8

.lib libs.tech/ngspice/sky130.lib.spice tt
.include libs.ref/sky130_fd_sc_hvl/spice/sky130_fd_sc_hvl.spice
.include libs.ref/sky130_fd_sc_hd/spice/sky130_fd_sc_hd.spice

*dig pull up/down to set test bits
R000 force_pdn dvss 1e9
R001 force_rc_osc dvss 1e9
R002 force_short_oneshot dvdd 1e9
R003 isrc_sel dvss 1e9

.temp 25
.save all
.save @m.xipor.xiana.xirsmux.xmena.msky130_fd_pr__nfet_g5v0d10v5[id]

.control
tran 10u 1400u
plot pwup_filt itest avdd force_pdn vbg_1v2 vin xipor.xiana.dcomp xipor.xiana.dcomp_filt
plot i(Vavdd) i(Vdvdd)
plot porb avdd pwup_filt
plot @m.xipor.xiana.xirsmux.xmena.msky130_fd_pr__nfet_g5v0d10v5[id]

.endc


**** end user architecture code
**.ends

* expanding   symbol:  xschem/por.sym # of pins=21
** sym_path: /home/rtsang/chipalooza/sky130_ajc_ip__por/xschem/por.sym
** sch_path: /home/rtsang/chipalooza/sky130_ajc_ip__por/xschem/por.sch
.subckt por porb_h avdd avss porb dvdd por dvss osc_ck vbg_1v2 osc_ck_256 otrip_2_ otrip_1_ otrip_0_ itest pwup_filt force_pdn vin
+ force_rc_osc force_short_oneshot startup_timed_out por_timed_out isrc_sel ibg_200n
*.ipin avdd
*.ipin avss
*.ipin dvdd
*.ipin dvss
*.ipin vbg_1v2
*.ipin otrip_2_,otrip_1_,otrip_0_
*.ipin force_pdn
*.ipin force_rc_osc
*.ipin force_short_oneshot
*.ipin isrc_sel
*.ipin ibg_200n
*.opin vin
*.opin porb_h
*.opin porb
*.opin por
*.opin osc_ck
*.opin osc_ck_256
*.opin pwup_filt
*.opin itest
*.opin startup_timed_out
*.opin por_timed_out
xIana otrip_decoded_7_ otrip_decoded_6_ otrip_decoded_5_ otrip_decoded_4_ otrip_decoded_3_ otrip_decoded_2_ otrip_decoded_1_
+ otrip_decoded_0_ vin vbg_1v2 avdd itest force_pdnb avss ibg_200n dvdd dvss isrc_sel pwup_filt osc_ck osc_ena porb_h por_unbuf por porb por_ana
**** begin user architecture code



*XSPICE CO-SIM netlist
.include por_dig.out.spice
xipor_dig dvss dvdd force_pdn force_pdnb force_rc_osc force_short_oneshot osc_ck osc_ck_256 osc_ena
+otrip_0_ otrip_1_ otrip_2_
+otrip_decoded_0_ otrip_decoded_1_ otrip_decoded_2_ otrip_decoded_3_ otrip_decoded_4_ otrip_decoded_5_ otrip_decoded_6_ otrip_decoded_7_
+por_timed_out por_unbuf pwup_filt startup_timed_out por_dig


**** end user architecture code
.ends


* expanding   symbol:  xschem/por_ana.sym # of pins=18
** sym_path: /home/rtsang/chipalooza/sky130_ajc_ip__por/xschem/por_ana.sym
** sch_path: /home/rtsang/chipalooza/sky130_ajc_ip__por/xschem/por_ana.sch
.subckt por_ana otrip_decoded_7_ otrip_decoded_6_ otrip_decoded_5_ otrip_decoded_4_ otrip_decoded_3_ otrip_decoded_2_
+ otrip_decoded_1_ otrip_decoded_0_ vin vbg_1v2 avdd itest force_pdnb avss ibg_200n dvdd dvss isrc_sel pwup_filt osc_ck osc_ena porb_h por_unbuf por
+ porb
*.ipin vbg_1v2
*.ipin avdd
*.ipin avss
*.ipin dvdd
*.ipin dvss
*.ipin force_pdnb
*.ipin isrc_sel
*.ipin ibg_200n
*.opin pwup_filt
*.opin itest
*.ipin osc_ena
*.opin osc_ck
*.ipin
*+ otrip_decoded_7_,otrip_decoded_6_,otrip_decoded_5_,otrip_decoded_4_,otrip_decoded_3_,otrip_decoded_2_,otrip_decoded_1_,otrip_decoded_0_
*.opin vin
*.ipin por_unbuf
*.opin porb_h
*.opin por
*.opin porb
XR1 dcomp_filt dcomp avss sky130_fd_pr__res_xhigh_po W=2 L=1000 mult=1 m=1
xIlvls0 dcomp_filt dvdd avss avss avdd avdd pwup_filt sky130_fd_sc_hvl__lsbufhv2lv_1
XC1 dcomp_filt avss sky130_fd_pr__cap_mim_m3_1 W=30 L=30 MF=3 m=3
XC2 dcomp_filt avss sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=3 m=3
xIlvls0_7_ otrip_decoded_7_ dvdd avss avss avdd avdd otrip_decoded_avdd_7_ sky130_fd_sc_hvl__lsbuflv2hv_1
xIlvls0_6_ otrip_decoded_6_ dvdd avss avss avdd avdd otrip_decoded_avdd_6_ sky130_fd_sc_hvl__lsbuflv2hv_1
xIlvls0_5_ otrip_decoded_5_ dvdd avss avss avdd avdd otrip_decoded_avdd_5_ sky130_fd_sc_hvl__lsbuflv2hv_1
xIlvls0_4_ otrip_decoded_4_ dvdd avss avss avdd avdd otrip_decoded_avdd_4_ sky130_fd_sc_hvl__lsbuflv2hv_1
xIlvls0_3_ otrip_decoded_3_ dvdd avss avss avdd avdd otrip_decoded_avdd_3_ sky130_fd_sc_hvl__lsbuflv2hv_1
xIlvls0_2_ otrip_decoded_2_ dvdd avss avss avdd avdd otrip_decoded_avdd_2_ sky130_fd_sc_hvl__lsbuflv2hv_1
xIlvls0_1_ otrip_decoded_1_ dvdd avss avss avdd avdd otrip_decoded_avdd_1_ sky130_fd_sc_hvl__lsbuflv2hv_1
xIlvls0_0_ otrip_decoded_0_ dvdd avss avss avdd avdd otrip_decoded_avdd_0_ sky130_fd_sc_hvl__lsbuflv2hv_1
xIlvls1 force_pdnb dvdd avss avss avdd avdd force_pdnb_avdd sky130_fd_sc_hvl__lsbuflv2hv_1
xIlvls2 isrc_sel dvdd avss avss avdd avdd isrc_sel_avdd sky130_fd_sc_hvl__lsbuflv2hv_1
xIrsmux avdd vin otrip_decoded_avdd_7_ otrip_decoded_avdd_6_ otrip_decoded_avdd_5_ otrip_decoded_avdd_4_ otrip_decoded_avdd_3_
+ otrip_decoded_avdd_2_ otrip_decoded_avdd_1_ otrip_decoded_avdd_0_ dvdd dvss force_pdnb_avdd avss rstring_mux
xIcomp avdd ibias dcomp force_pdnb_avdd vbg_1v2 vin avss comparator
xIbiasgen avdd itest ibias ibg_200n vbg_1v2 isrc_sel_avdd force_pdnb_avdd avss ibias_gen
xIosc dvdd osc_ck osc_ena dvss rc_osc
xIlvls3 por_unbuf dvdd avss avss avdd avdd net1 sky130_fd_sc_hvl__lsbuflv2hv_1
xIinv1 net1 avss avss avdd avdd net2 sky130_fd_sc_hvl__inv_1
xIinv2 net2 avss avss avdd avdd net3 sky130_fd_sc_hvl__inv_4
xIinv3 net3 avss avss avdd avdd porb_h sky130_fd_sc_hvl__inv_16
xIinv4 por_unbuf dvss dvss dvdd dvdd net4 sky130_fd_sc_hd__inv_4
xIinv5 net4 dvss dvss dvdd dvdd por sky130_fd_sc_hd__inv_16
xIinv7 net6 dvss dvss dvdd dvdd net5 sky130_fd_sc_hd__inv_4
xIinv88 net5 dvss dvss dvdd dvdd porb sky130_fd_sc_hd__inv_16
xIinv6 por_unbuf dvss dvss dvdd dvdd net6 sky130_fd_sc_hd__inv_1
.ends


* expanding   symbol:  rstring_mux.sym # of pins=7
** sym_path: /home/rtsang/chipalooza/sky130_ajc_ip__por/xschem/rstring_mux.sym
** sch_path: /home/rtsang/chipalooza/sky130_ajc_ip__por/xschem/rstring_mux.sch
.subckt rstring_mux avdd vout otrip_decoded_avdd_7_ otrip_decoded_avdd_6_ otrip_decoded_avdd_5_ otrip_decoded_avdd_4_
+ otrip_decoded_avdd_3_ otrip_decoded_avdd_2_ otrip_decoded_avdd_1_ otrip_decoded_avdd_0_ dvdd dvss ena avss
*.ipin avdd
*.ipin avss
*.opin vout
*.ipin ena
*.ipin
*+ otrip_decoded_avdd_7_,otrip_decoded_avdd_6_,otrip_decoded_avdd_5_,otrip_decoded_avdd_4_,otrip_decoded_avdd_3_,otrip_decoded_avdd_2_,otrip_decoded_avdd_1_,otrip_decoded_avdd_0_
*.ipin dvss
*.ipin dvdd
XR1 net2 net3 avss sky130_fd_pr__res_xhigh_po W=2 L=50 mult=1 m=1
XR2 net3 net4 avss sky130_fd_pr__res_xhigh_po W=2 L=50 mult=1 m=1
XR0 net1 net2 avss sky130_fd_pr__res_xhigh_po W=2 L=50 mult=1 m=1
XR3 net4 net5 avss sky130_fd_pr__res_xhigh_po W=2 L=50 mult=1 m=1
XR4 net5 net6 avss sky130_fd_pr__res_xhigh_po W=2 L=50 mult=1 m=1
XR5 net6 net7 avss sky130_fd_pr__res_xhigh_po W=2 L=50 mult=1 m=1
XR6 net7 net8 avss sky130_fd_pr__res_xhigh_po W=2 L=50 mult=1 m=1
XR7 net8 net9 avss sky130_fd_pr__res_xhigh_po W=2 L=50 mult=1 m=1
XR8 net9 net10 avss sky130_fd_pr__res_xhigh_po W=2 L=50 mult=1 m=1
XR9 net10 net11 avss sky130_fd_pr__res_xhigh_po W=2 L=50 mult=1 m=1
XR10 net11 net12 avss sky130_fd_pr__res_xhigh_po W=2 L=50 mult=1 m=1
XR11 net12 net13 avss sky130_fd_pr__res_xhigh_po W=2 L=50 mult=1 m=1
XR12 net13 net14 avss sky130_fd_pr__res_xhigh_po W=2 L=50 mult=1 m=1
XR13 net14 net15 avss sky130_fd_pr__res_xhigh_po W=2 L=50 mult=1 m=1
XR14 net15 net16 avss sky130_fd_pr__res_xhigh_po W=2 L=50 mult=1 m=1
XR15 net16 net17 avss sky130_fd_pr__res_xhigh_po W=2 L=50 mult=1 m=1
XR16 net17 net18 avss sky130_fd_pr__res_xhigh_po W=2 L=50 mult=1 m=1
XR17 net18 net19 avss sky130_fd_pr__res_xhigh_po W=2 L=50 mult=1 m=1
XR18 net19 net20 avss sky130_fd_pr__res_xhigh_po W=2 L=50 mult=1 m=1
XR19 net20 net21 avss sky130_fd_pr__res_xhigh_po W=2 L=50 mult=1 m=1
XR20 net21 net22 avss sky130_fd_pr__res_xhigh_po W=2 L=50 mult=1 m=1
XR21 net22 net23 avss sky130_fd_pr__res_xhigh_po W=2 L=50 mult=1 m=1
XR22 net23 net24 avss sky130_fd_pr__res_xhigh_po W=2 L=50 mult=1 m=1
XR23 net24 net25 avss sky130_fd_pr__res_xhigh_po W=2 L=50 mult=1 m=1
XR24 net25 net26 avss sky130_fd_pr__res_xhigh_po W=2 L=50 mult=1 m=1
XR25 net26 net27 avss sky130_fd_pr__res_xhigh_po W=2 L=50 mult=1 m=1
XR26 net27 net28 avss sky130_fd_pr__res_xhigh_po W=2 L=50 mult=1 m=1
XR27 net28 vtrip7 avss sky130_fd_pr__res_xhigh_po W=2 L=50 mult=1 m=1
XR28 vtrip7 vtrip6 avss sky130_fd_pr__res_xhigh_po W=2 L=50 mult=1 m=1
XR29 vtrip6 vtrip5 avss sky130_fd_pr__res_xhigh_po W=2 L=50 mult=1 m=1
XR30 vtrip5 vtrip4 avss sky130_fd_pr__res_xhigh_po W=2 L=50 mult=1 m=1
XR31 vtrip4 vtrip3 avss sky130_fd_pr__res_xhigh_po W=2 L=50 mult=1 m=1
XR32 vtrip3 vtrip2 avss sky130_fd_pr__res_xhigh_po W=2 L=50 mult=1 m=1
XR33 vtrip2 vtrip1 avss sky130_fd_pr__res_xhigh_po W=2 L=50 mult=1 m=1
XR34 vtrip1 vtrip0 avss sky130_fd_pr__res_xhigh_po W=2 L=50 mult=1 m=1
XR35 vtrip0 net29 avss sky130_fd_pr__res_xhigh_po W=2 L=50 mult=1 m=1
XR36 net29 net30 avss sky130_fd_pr__res_xhigh_po W=2 L=50 mult=1 m=1
XR37 net30 net31 avss sky130_fd_pr__res_xhigh_po W=2 L=50 mult=1 m=1
XR38 net31 net32 avss sky130_fd_pr__res_xhigh_po W=2 L=50 mult=1 m=1
XR39 net32 net33 avss sky130_fd_pr__res_xhigh_po W=2 L=50 mult=1 m=1
XR40 net33 net34 avss sky130_fd_pr__res_xhigh_po W=2 L=50 mult=1 m=1
XR41 net34 net35 avss sky130_fd_pr__res_xhigh_po W=2 L=50 mult=1 m=1
XR42 net35 net36 avss sky130_fd_pr__res_xhigh_po W=2 L=50 mult=1 m=1
XR43 net36 net37 avss sky130_fd_pr__res_xhigh_po W=2 L=50 mult=1 m=1
XR44 net37 net38 avss sky130_fd_pr__res_xhigh_po W=2 L=50 mult=1 m=1
XR45 net38 net39 avss sky130_fd_pr__res_xhigh_po W=2 L=50 mult=1 m=1
XR46 net39 net40 avss sky130_fd_pr__res_xhigh_po W=2 L=50 mult=1 m=1
XR47 net40 net41 avss sky130_fd_pr__res_xhigh_po W=2 L=50 mult=1 m=1
XR48 net41 net42 avss sky130_fd_pr__res_xhigh_po W=2 L=50 mult=1 m=1
XR49 net42 net43 avss sky130_fd_pr__res_xhigh_po W=2 L=50 mult=1 m=1
XR50 net43 net44 avss sky130_fd_pr__res_xhigh_po W=2 L=50 mult=1 m=1
XR51 net44 net45 avss sky130_fd_pr__res_xhigh_po W=2 L=50 mult=1 m=1
XR52 net45 net46 avss sky130_fd_pr__res_xhigh_po W=2 L=50 mult=1 m=1
XR53 net46 net47 avss sky130_fd_pr__res_xhigh_po W=2 L=50 mult=1 m=1
XR54 net47 net48 avss sky130_fd_pr__res_xhigh_po W=2 L=50 mult=1 m=1
XR55 net48 net49 avss sky130_fd_pr__res_xhigh_po W=2 L=50 mult=1 m=1
XR56 net49 net50 avss sky130_fd_pr__res_xhigh_po W=2 L=50 mult=1 m=1
XR57 net50 net51 avss sky130_fd_pr__res_xhigh_po W=2 L=50 mult=1 m=1
XR58 net51 net52 avss sky130_fd_pr__res_xhigh_po W=2 L=50 mult=1 m=1
XR59 net52 net53 avss sky130_fd_pr__res_xhigh_po W=2 L=50 mult=1 m=1
XR60 net53 net54 avss sky130_fd_pr__res_xhigh_po W=2 L=50 mult=1 m=1
XR61 net54 net55 avss sky130_fd_pr__res_xhigh_po W=2 L=50 mult=1 m=1
XR62 net55 net56 avss sky130_fd_pr__res_xhigh_po W=2 L=50 mult=1 m=1
XR63 net56 net57 avss sky130_fd_pr__res_xhigh_po W=2 L=50 mult=1 m=1
XR64 net57 net58 avss sky130_fd_pr__res_xhigh_po W=2 L=50 mult=1 m=1
XR65 net58 net59 avss sky130_fd_pr__res_xhigh_po W=2 L=50 mult=1 m=1
XR66 net59 net60 avss sky130_fd_pr__res_xhigh_po W=2 L=50 mult=1 m=1
XR67 net60 net61 avss sky130_fd_pr__res_xhigh_po W=2 L=50 mult=1 m=1
XR68 net61 net62 avss sky130_fd_pr__res_xhigh_po W=2 L=50 mult=1 m=1
XR69 net62 avdd avss sky130_fd_pr__res_xhigh_po W=2 L=50 mult=1 m=1
XMtp_7_ vtrip7 otrip_decoded_b_avdd_7_ vout avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XMtp_6_ vtrip6 otrip_decoded_b_avdd_6_ vout avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XMtp_5_ vtrip5 otrip_decoded_b_avdd_5_ vout avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XMtp_4_ vtrip4 otrip_decoded_b_avdd_4_ vout avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XMtp_3_ vtrip3 otrip_decoded_b_avdd_3_ vout avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XMtp_2_ vtrip2 otrip_decoded_b_avdd_2_ vout avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XMtp_1_ vtrip1 otrip_decoded_b_avdd_1_ vout avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XMtp_0_ vtrip0 otrip_decoded_b_avdd_0_ vout avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XMtn_7_ vout otrip_decoded_avdd_7_ vtrip7 avss sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XMtn_6_ vout otrip_decoded_avdd_6_ vtrip6 avss sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XMtn_5_ vout otrip_decoded_avdd_5_ vtrip5 avss sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XMtn_4_ vout otrip_decoded_avdd_4_ vtrip4 avss sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XMtn_3_ vout otrip_decoded_avdd_3_ vtrip3 avss sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XMtn_2_ vout otrip_decoded_avdd_2_ vtrip2 avss sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XMtn_1_ vout otrip_decoded_avdd_1_ vtrip1 avss sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XMtn_0_ vout otrip_decoded_avdd_0_ vtrip0 avss sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XMena net1 ena avss avss sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=16 m=16
xIinv_7_ otrip_decoded_avdd_7_ avss avss avdd avdd otrip_decoded_b_avdd_7_ sky130_fd_sc_hvl__inv_1
xIinv_6_ otrip_decoded_avdd_6_ avss avss avdd avdd otrip_decoded_b_avdd_6_ sky130_fd_sc_hvl__inv_1
xIinv_5_ otrip_decoded_avdd_5_ avss avss avdd avdd otrip_decoded_b_avdd_5_ sky130_fd_sc_hvl__inv_1
xIinv_4_ otrip_decoded_avdd_4_ avss avss avdd avdd otrip_decoded_b_avdd_4_ sky130_fd_sc_hvl__inv_1
xIinv_3_ otrip_decoded_avdd_3_ avss avss avdd avdd otrip_decoded_b_avdd_3_ sky130_fd_sc_hvl__inv_1
xIinv_2_ otrip_decoded_avdd_2_ avss avss avdd avdd otrip_decoded_b_avdd_2_ sky130_fd_sc_hvl__inv_1
xIinv_1_ otrip_decoded_avdd_1_ avss avss avdd avdd otrip_decoded_b_avdd_1_ sky130_fd_sc_hvl__inv_1
xIinv_0_ otrip_decoded_avdd_0_ avss avss avdd avdd otrip_decoded_b_avdd_0_ sky130_fd_sc_hvl__inv_1
.ends


* expanding   symbol:  comparator.sym # of pins=7
** sym_path: /home/rtsang/chipalooza/sky130_ajc_ip__por/xschem/comparator.sym
** sch_path: /home/rtsang/chipalooza/sky130_ajc_ip__por/xschem/comparator.sch
.subckt comparator avdd ibias out ena vinn vinp avss
*.ipin ena
*.ipin avdd
*.ipin avss
*.ipin ibias
*.ipin vinn
*.ipin vinp
*.opin out
XMb vn vn avss avss sky130_fd_pr__nfet_g5v0d10v5 L=8 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XMta vt vn avss avss sky130_fd_pr__nfet_g5v0d10v5 L=8 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XMl0 vn ena_b avss avss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMinv0 ena_b ena avss avss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMinv1 ena_b ena avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMi0 vnn vinn vt vt sky130_fd_pr__nfet_g5v0d10v5 L=8 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=4 m=4
XMi1 vpp vinp vt vt sky130_fd_pr__nfet_g5v0d10v5 L=8 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=4 m=4
XMld1 vpp vpp avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=8 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XMh1 vnn vpp avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XMh0 vpp vnn avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XMld0 vnn vnn avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=8 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XMpp1 n0 vpp avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=8 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XMnn1 n0 vm avss avss sky130_fd_pr__nfet_g5v0d10v5 L=8 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XMpp0 vm vnn avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=8 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XMnn0 vm vm avss avss sky130_fd_pr__nfet_g5v0d10v5 L=8 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XMinv3 n1 n0 avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XMinv2 n1 n0 avss avss sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XMinv5 out n1 avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=8 m=8
XMinv4 out n1 avss avss sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=8 m=8
XMl1 vm ena_b avss avss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMl3 vnn ena avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMl4 vpp ena avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMt1 ibias ena vn avss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMt0 vn ena_b ibias avdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMl2 n0 ena_b avss avss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  ibias_gen.sym # of pins=8
** sym_path: /home/rtsang/chipalooza/sky130_ajc_ip__por/xschem/ibias_gen.sym
** sch_path: /home/rtsang/chipalooza/sky130_ajc_ip__por/xschem/ibias_gen.sch
.subckt ibias_gen avdd itest ibias ibg_200n vbg_1v2 isrc_sel ena avss
*.ipin vbg_1v2
*.ipin ena
*.opin ibias
*.ipin ibg_200n
*.ipin isrc_sel
*.ipin avdd
*.ipin avss
*.opin itest
XR1 avss net3 avss sky130_fd_pr__res_xhigh_po W=2 L=1000 mult=1 m=1
XQ1 avss avss net2 sky130_fd_pr__pnp_05v5_W0p68L0p68 m=1 mult=1
XM17 net1 vbg_1v2 vn0 avss sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=10 m=10
XMt9 net1 ena_b net4 avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMn0 vn0 vn0 net2 avss sky130_fd_pr__nfet_g5v0d10v5 L=4 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XMp0 vn0 vp0 avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=4 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XMn1 vp0 vn0 net3 avss sky130_fd_pr__nfet_g5v0d10v5 L=4 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XMp1 vp0 vp0 avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=4 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XMp ibias vp avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=4 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XMt0 vp0 isrc_sel vp avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMt1 vp isrc_sel_b vp0 avss sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMl6 vp ena avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=2 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMl3 vp0 ena avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=2 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMl1 vn0 ena_b avss avss sky130_fd_pr__nfet_g5v0d10v5 L=2 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMnn1 vp1 vn1 avss avss sky130_fd_pr__nfet_g5v0d10v5 L=8 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=8 m=8
XMnn0 vn1 vn1 avss avss sky130_fd_pr__nfet_g5v0d10v5 L=8 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XMl9 vn1 isrc_sel_b avss avss sky130_fd_pr__nfet_g5v0d10v5 L=2 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMt6 net5 isrc_sel vn1 avss sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMt7 vn1 isrc_sel_b net6 avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMpp1 vp1 vp1 avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=4 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XMt2 vp isrc_sel_b vp1 avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMt3 vp1 isrc_sel vp avss sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMt4 ibg_200n ena net5 avss sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMt5 net6 ena_b ibg_200n avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMl7 vp1 isrc_sel avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=2 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMl8 vp1 ena avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=2 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMl10 vn1 ena_b avss avss sky130_fd_pr__nfet_g5v0d10v5 L=2 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMl2 vp0 isrc_sel_b avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=2 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMl0 vn0 isrc_sel avss avss sky130_fd_pr__nfet_g5v0d10v5 L=2 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMt8 net4 isrc_sel avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMn2 ena_b ena avss avss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMp2 ena_b ena avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMn3 isrc_sel_b isrc_sel avss avss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMp3 isrc_sel_b isrc_sel avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMtst itest vp avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=4 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
.ends


* expanding   symbol:  rc_osc.sym # of pins=4
** sym_path: /home/rtsang/chipalooza/sky130_ajc_ip__por/xschem/rc_osc.sym
** sch_path: /home/rtsang/chipalooza/sky130_ajc_ip__por/xschem/rc_osc.sch
.subckt rc_osc dvdd out ena dvss
*.ipin dvdd
*.ipin dvss
*.opin out
*.ipin ena
XM1 m in dvss dvss sky130_fd_pr__nfet_01v8 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XM3 m in dvdd dvdd sky130_fd_pr__pfet_01v8 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=4 m=4
XM2 m n dvss dvss sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM4 m n dvdd dvdd sky130_fd_pr__pfet_01v8 L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XM5 n m dvss dvss sky130_fd_pr__nfet_01v8 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM6 n m dvdd dvdd sky130_fd_pr__pfet_01v8 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XM7 out n dvss dvss sky130_fd_pr__nfet_01v8 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM8 out n dvdd dvdd sky130_fd_pr__pfet_01v8 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XC1 in dvss sky130_fd_pr__cap_mim_m3_1 W=25 L=25 MF=1 m=1
XR1 in net1 dvss sky130_fd_pr__res_xhigh_po W=2 L=305 mult=1 m=1
XM12 in ena dvdd dvdd sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XC2 in dvss sky130_fd_pr__cap_mim_m3_2 W=25 L=25 MF=1 m=1
XM9 out ena net1 dvss sky130_fd_pr__nfet_01v8 L=0.18 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM10 out ena_b net1 dvdd sky130_fd_pr__pfet_01v8 L=0.18 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM11 ena_b ena dvss dvss sky130_fd_pr__nfet_01v8 L=0.6 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM13 ena_b ena dvdd dvdd sky130_fd_pr__pfet_01v8 L=0.6 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends

.GLOBAL GND
.end
