* NGSPICE file created from por_ana.ext - technology: sky130A

.subckt sky130_fd_sc_hd__inv_16 A VGND VNB VPB VPWR Y
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X16 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X17 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X18 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X19 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X20 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X21 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X22 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X23 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X24 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X25 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X26 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X27 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X28 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X29 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X30 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X31 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
C0 Y A 1.4347f
C1 VGND Y 1.06261f
C2 VPB VPWR 0.159316f
C3 A VPB 0.525745f
C4 A VPWR 0.280261f
C5 VGND VPWR 0.160762f
C6 Y VPWR 1.46621f
C7 VGND A 0.265874f
C8 VGND VNB 0.864536f
C9 VPWR VNB 0.737072f
C10 A VNB 1.54575f
C11 VPB VNB 1.49072f
.ends

.subckt sky130_fd_sc_hvl__lsbufhv2lv_1 A LVPWR VGND VNB VPB VPWR X
X0 a_30_1337# A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.1197 ps=1.41 w=0.42 l=0.5
X1 VGND a_30_1337# a_30_207# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.178875 pd=1.26 as=0.1197 ps=1.41 w=0.42 l=0.5
X2 VGND a_30_207# a_389_141# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.105 ps=1.03 w=0.75 l=0.5
X3 VGND a_30_207# a_389_141# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.19875 ps=2.03 w=0.75 l=0.5
X4 a_389_1337# a_30_1337# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.105 ps=1.03 w=0.75 l=0.5
X5 VGND a_30_207# a_389_141# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.19875 ps=2.03 w=0.75 l=0.5
X6 VGND A a_30_1337# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.178875 pd=1.26 as=0.1197 ps=1.41 w=0.42 l=0.5
X7 VGND a_30_1337# a_389_1337# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.19875 ps=2.03 w=0.75 l=0.5
X8 a_389_141# a_30_207# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.178875 ps=1.26 w=0.75 l=0.5
X9 VGND a_30_1337# a_389_1337# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X10 LVPWR a_389_141# X LVPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1568 pd=1.4 as=0.2968 ps=2.77 w=1.12 l=0.15
X11 VGND a_389_141# X VNB sky130_fd_pr__nfet_01v8 ad=0.1961 pd=2.01 as=0.1961 ps=2.01 w=0.74 l=0.15
X12 a_389_1337# a_30_1337# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.178875 ps=1.26 w=0.75 l=0.5
X13 LVPWR a_389_1337# a_389_141# LVPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2968 pd=2.77 as=0.2968 ps=2.77 w=1.12 l=0.15
X14 a_30_207# a_30_1337# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.1197 ps=1.41 w=0.42 l=0.5
X15 a_389_1337# a_389_141# LVPWR LVPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2968 pd=2.77 as=0.1568 ps=1.4 w=1.12 l=0.15
C0 LVPWR X 0.171836f
C1 a_389_141# a_30_1337# 0.166612f
C2 a_30_207# a_30_1337# 0.170258f
C3 VPWR a_389_1337# 0.113209f
C4 VGND X 0.22925f
C5 VPWR VPB 2.11464f
C6 LVPWR VPWR 1.07584f
C7 a_389_141# X 0.116307f
C8 VGND VPWR 0.179222f
C9 LVPWR a_389_1337# 0.443515f
C10 A a_30_1337# 0.187128f
C11 VGND a_389_1337# 0.349538f
C12 VPWR a_389_141# 0.164733f
C13 LVPWR VGND 0.248568f
C14 VPWR a_30_1337# 0.215762f
C15 a_389_141# a_389_1337# 0.136815f
C16 a_30_1337# a_389_1337# 0.249533f
C17 LVPWR a_389_141# 0.469283f
C18 a_30_1337# VPB 0.29963f
C19 VGND a_389_141# 0.378288f
C20 a_30_207# VGND 0.254325f
C21 VGND a_30_1337# 0.296817f
C22 A VPB 0.193945f
C23 a_30_207# a_389_141# 0.249269f
C24 VPWR VNB 0.294478f
C25 VGND VNB 2.76278f
C26 A VNB 0.284924f
C27 LVPWR VNB 0.712212f
C28 VPB VNB 1.87844f
C29 a_30_207# VNB 0.665049f
C30 a_389_141# VNB 0.635783f
C31 a_389_1337# VNB 0.510776f
C32 a_30_1337# VNB 1.03613f
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_K8JYEQ a_n3678_n531# a_296_n557# a_950_n531#
+ a_n2374_n557# a_3976_n531# a_2908_n531# a_n1306_n557# a_n3442_n557# a_n2076_n531#
+ a_n3144_n531# a_2610_n557# a_1542_n557# a_n950_n557# a_n1008_n531# a_n4212_n531#
+ a_3442_n531# a_2374_n531# a_1306_n531# a_n652_n531# a_1898_n557# a_n3798_n557# a_2966_n557#
+ a_772_n531# a_118_n557# a_3798_n531# a_n1720_n531# a_n1128_n557# a_n2196_n557# a_n3264_n557#
+ a_1364_n557# a_3500_n557# a_2432_n557# a_n772_n557# a_2196_n531# a_n474_n531# a_n4034_n531#
+ a_3264_n531# a_1128_n531# a_830_n557# a_3856_n557# a_2788_n557# a_n1840_n557# a_594_n531#
+ a_n1542_n531# a_n2610_n531# a_n3086_n557# a_2254_n557# a_1186_n557# a_n594_n557#
+ a_n2018_n557# a_n4154_n557# a_1840_n531# a_3322_n557# a_3086_n531# a_n296_n531#
+ a_n1898_n531# a_n2966_n531# a_4154_n531# a_2018_n531# a_60_n531# a_652_n557# a_3678_n557#
+ a_n1662_n557# a_n2730_n557# a_n1364_n531# a_n60_n557# a_416_n531# a_n2432_n531#
+ a_1662_n531# a_n3500_n531# a_3144_n557# a_2076_n557# a_1008_n557# a_2730_n531# a_n416_n557#
+ a_n2788_n531# a_n3856_n531# a_474_n557# a_n118_n531# a_n1484_n557# a_n2552_n557#
+ a_n3620_n557# a_238_n531# a_n1186_n531# a_n2254_n531# a_1720_n557# a_n3322_n531#
+ a_n4346_n691# a_2552_n531# a_1484_n531# a_n830_n531# a_4034_n557# a_n3976_n557#
+ a_3620_n531# a_n238_n557# a_n2908_n557#
X0 a_n3856_n531# a_n3976_n557# a_n4034_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X1 a_2196_n531# a_2076_n557# a_2018_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X2 a_n2610_n531# a_n2730_n557# a_n2788_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X3 a_n2254_n531# a_n2374_n557# a_n2432_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X4 a_n652_n531# a_n772_n557# a_n830_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X5 a_2018_n531# a_1898_n557# a_1840_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X6 a_n1008_n531# a_n1128_n557# a_n1186_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X7 a_594_n531# a_474_n557# a_416_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X8 a_3264_n531# a_3144_n557# a_3086_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X9 a_n3322_n531# a_n3442_n557# a_n3500_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X10 a_60_n531# a_n60_n557# a_n118_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X11 a_3086_n531# a_2966_n557# a_2908_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X12 a_1484_n531# a_1364_n557# a_1306_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X13 a_n1542_n531# a_n1662_n557# a_n1720_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X14 a_2552_n531# a_2432_n557# a_2374_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X15 a_n3678_n531# a_n3798_n557# a_n3856_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X16 a_950_n531# a_830_n557# a_772_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X17 a_3620_n531# a_3500_n557# a_3442_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X18 a_n2076_n531# a_n2196_n557# a_n2254_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X19 a_n830_n531# a_n950_n557# a_n1008_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X20 a_n474_n531# a_n594_n557# a_n652_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X21 a_1840_n531# a_1720_n557# a_1662_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X22 a_n3500_n531# a_n3620_n557# a_n3678_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X23 a_416_n531# a_296_n557# a_238_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X24 a_n3144_n531# a_n3264_n557# a_n3322_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X25 a_2908_n531# a_2788_n557# a_2730_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X26 a_n1898_n531# a_n2018_n557# a_n2076_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X27 a_4154_n531# a_4034_n557# a_3976_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=0.6
X28 a_n296_n531# a_n416_n557# a_n474_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X29 a_1306_n531# a_1186_n557# a_1128_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X30 a_3976_n531# a_3856_n557# a_3798_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X31 a_n1720_n531# a_n1840_n557# a_n1898_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X32 a_n1364_n531# a_n1484_n557# a_n1542_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X33 a_238_n531# a_118_n557# a_60_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X34 a_2374_n531# a_2254_n557# a_2196_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X35 a_n2788_n531# a_n2908_n557# a_n2966_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X36 a_n2432_n531# a_n2552_n557# a_n2610_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X37 a_1128_n531# a_1008_n557# a_950_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X38 a_n1186_n531# a_n1306_n557# a_n1364_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X39 a_772_n531# a_652_n557# a_594_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X40 a_3442_n531# a_3322_n557# a_3264_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X41 a_1662_n531# a_1542_n557# a_1484_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X42 a_n2966_n531# a_n3086_n557# a_n3144_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X43 a_2730_n531# a_2610_n557# a_2552_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X44 a_n4034_n531# a_n4154_n557# a_n4212_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=0.6
X45 a_n118_n531# a_n238_n557# a_n296_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X46 a_3798_n531# a_3678_n557# a_3620_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
C0 a_n2788_n531# a_n2610_n531# 0.396241f
C1 a_1306_n531# a_1128_n531# 0.396241f
C2 a_1484_n531# a_1662_n531# 0.396241f
C3 a_n1898_n531# a_n2076_n531# 0.396241f
C4 a_3264_n531# a_3442_n531# 0.396241f
C5 a_3442_n531# a_3620_n531# 0.396241f
C6 a_n3678_n531# a_n3856_n531# 0.396241f
C7 a_2196_n531# a_2374_n531# 0.396241f
C8 a_n1186_n531# a_n1008_n531# 0.396241f
C9 a_3620_n531# a_3798_n531# 0.396241f
C10 a_238_n531# a_416_n531# 0.396241f
C11 a_1662_n531# a_1840_n531# 0.396241f
C12 a_416_n531# a_594_n531# 0.396241f
C13 a_2018_n531# a_2196_n531# 0.396241f
C14 a_2374_n531# a_2552_n531# 0.396241f
C15 a_n1008_n531# a_n830_n531# 0.396241f
C16 a_3798_n531# a_3976_n531# 0.396241f
C17 a_n4212_n531# a_n4034_n531# 0.396241f
C18 a_1840_n531# a_2018_n531# 0.396241f
C19 a_3086_n531# a_3264_n531# 0.396241f
C20 a_2552_n531# a_2730_n531# 0.396241f
C21 a_n830_n531# a_n652_n531# 0.396241f
C22 a_3976_n531# a_4154_n531# 0.396241f
C23 a_60_n531# a_238_n531# 0.396241f
C24 a_n3500_n531# a_n3322_n531# 0.396241f
C25 a_n4034_n531# a_n3856_n531# 0.396241f
C26 a_2730_n531# a_2908_n531# 0.396241f
C27 a_n474_n531# a_n652_n531# 0.396241f
C28 a_n2610_n531# a_n2432_n531# 0.396241f
C29 a_n1898_n531# a_n1720_n531# 0.396241f
C30 a_594_n531# a_772_n531# 0.396241f
C31 a_n3144_n531# a_n2966_n531# 0.396241f
C32 a_n2432_n531# a_n2254_n531# 0.396241f
C33 a_n1720_n531# a_n1542_n531# 0.396241f
C34 a_n474_n531# a_n296_n531# 0.396241f
C35 a_n3678_n531# a_n3500_n531# 0.396241f
C36 a_n2966_n531# a_n2788_n531# 0.396241f
C37 a_n2254_n531# a_n2076_n531# 0.396241f
C38 a_n1542_n531# a_n1364_n531# 0.396241f
C39 a_n296_n531# a_n118_n531# 0.396241f
C40 a_772_n531# a_950_n531# 0.396241f
C41 a_n118_n531# a_60_n531# 0.396241f
C42 a_1306_n531# a_1484_n531# 0.396241f
C43 a_950_n531# a_1128_n531# 0.396241f
C44 a_n1186_n531# a_n1364_n531# 0.396241f
C45 a_n3144_n531# a_n3322_n531# 0.396241f
C46 a_2908_n531# a_3086_n531# 0.396241f
C47 a_4154_n531# a_n4346_n691# 0.533824f
C48 a_3976_n531# a_n4346_n691# 0.125488f
C49 a_3798_n531# a_n4346_n691# 0.125488f
C50 a_3620_n531# a_n4346_n691# 0.125488f
C51 a_3442_n531# a_n4346_n691# 0.125488f
C52 a_3264_n531# a_n4346_n691# 0.125488f
C53 a_3086_n531# a_n4346_n691# 0.125488f
C54 a_2908_n531# a_n4346_n691# 0.125488f
C55 a_2730_n531# a_n4346_n691# 0.125488f
C56 a_2552_n531# a_n4346_n691# 0.125488f
C57 a_2374_n531# a_n4346_n691# 0.125488f
C58 a_2196_n531# a_n4346_n691# 0.125488f
C59 a_2018_n531# a_n4346_n691# 0.125488f
C60 a_1840_n531# a_n4346_n691# 0.125488f
C61 a_1662_n531# a_n4346_n691# 0.125488f
C62 a_1484_n531# a_n4346_n691# 0.125488f
C63 a_1306_n531# a_n4346_n691# 0.125488f
C64 a_1128_n531# a_n4346_n691# 0.125488f
C65 a_950_n531# a_n4346_n691# 0.125488f
C66 a_772_n531# a_n4346_n691# 0.125488f
C67 a_594_n531# a_n4346_n691# 0.125488f
C68 a_416_n531# a_n4346_n691# 0.125488f
C69 a_238_n531# a_n4346_n691# 0.125488f
C70 a_60_n531# a_n4346_n691# 0.125488f
C71 a_n118_n531# a_n4346_n691# 0.125488f
C72 a_n296_n531# a_n4346_n691# 0.125488f
C73 a_n474_n531# a_n4346_n691# 0.125488f
C74 a_n652_n531# a_n4346_n691# 0.125488f
C75 a_n830_n531# a_n4346_n691# 0.125488f
C76 a_n1008_n531# a_n4346_n691# 0.125488f
C77 a_n1186_n531# a_n4346_n691# 0.125488f
C78 a_n1364_n531# a_n4346_n691# 0.125488f
C79 a_n1542_n531# a_n4346_n691# 0.125488f
C80 a_n1720_n531# a_n4346_n691# 0.125488f
C81 a_n1898_n531# a_n4346_n691# 0.125488f
C82 a_n2076_n531# a_n4346_n691# 0.125488f
C83 a_n2254_n531# a_n4346_n691# 0.125488f
C84 a_n2432_n531# a_n4346_n691# 0.125488f
C85 a_n2610_n531# a_n4346_n691# 0.125488f
C86 a_n2788_n531# a_n4346_n691# 0.125488f
C87 a_n2966_n531# a_n4346_n691# 0.125488f
C88 a_n3144_n531# a_n4346_n691# 0.125488f
C89 a_n3322_n531# a_n4346_n691# 0.125488f
C90 a_n3500_n531# a_n4346_n691# 0.125488f
C91 a_n3678_n531# a_n4346_n691# 0.125488f
C92 a_n3856_n531# a_n4346_n691# 0.125488f
C93 a_n4034_n531# a_n4346_n691# 0.125488f
C94 a_n4212_n531# a_n4346_n691# 0.533824f
C95 a_4034_n557# a_n4346_n691# 0.307672f
C96 a_3856_n557# a_n4346_n691# 0.27141f
C97 a_3678_n557# a_n4346_n691# 0.27141f
C98 a_3500_n557# a_n4346_n691# 0.27141f
C99 a_3322_n557# a_n4346_n691# 0.27141f
C100 a_3144_n557# a_n4346_n691# 0.27141f
C101 a_2966_n557# a_n4346_n691# 0.27141f
C102 a_2788_n557# a_n4346_n691# 0.27141f
C103 a_2610_n557# a_n4346_n691# 0.27141f
C104 a_2432_n557# a_n4346_n691# 0.27141f
C105 a_2254_n557# a_n4346_n691# 0.27141f
C106 a_2076_n557# a_n4346_n691# 0.27141f
C107 a_1898_n557# a_n4346_n691# 0.27141f
C108 a_1720_n557# a_n4346_n691# 0.27141f
C109 a_1542_n557# a_n4346_n691# 0.27141f
C110 a_1364_n557# a_n4346_n691# 0.27141f
C111 a_1186_n557# a_n4346_n691# 0.27141f
C112 a_1008_n557# a_n4346_n691# 0.27141f
C113 a_830_n557# a_n4346_n691# 0.27141f
C114 a_652_n557# a_n4346_n691# 0.27141f
C115 a_474_n557# a_n4346_n691# 0.27141f
C116 a_296_n557# a_n4346_n691# 0.27141f
C117 a_118_n557# a_n4346_n691# 0.27141f
C118 a_n60_n557# a_n4346_n691# 0.27141f
C119 a_n238_n557# a_n4346_n691# 0.27141f
C120 a_n416_n557# a_n4346_n691# 0.27141f
C121 a_n594_n557# a_n4346_n691# 0.27141f
C122 a_n772_n557# a_n4346_n691# 0.27141f
C123 a_n950_n557# a_n4346_n691# 0.27141f
C124 a_n1128_n557# a_n4346_n691# 0.27141f
C125 a_n1306_n557# a_n4346_n691# 0.27141f
C126 a_n1484_n557# a_n4346_n691# 0.27141f
C127 a_n1662_n557# a_n4346_n691# 0.27141f
C128 a_n1840_n557# a_n4346_n691# 0.27141f
C129 a_n2018_n557# a_n4346_n691# 0.27141f
C130 a_n2196_n557# a_n4346_n691# 0.27141f
C131 a_n2374_n557# a_n4346_n691# 0.27141f
C132 a_n2552_n557# a_n4346_n691# 0.27141f
C133 a_n2730_n557# a_n4346_n691# 0.27141f
C134 a_n2908_n557# a_n4346_n691# 0.27141f
C135 a_n3086_n557# a_n4346_n691# 0.27141f
C136 a_n3264_n557# a_n4346_n691# 0.27141f
C137 a_n3442_n557# a_n4346_n691# 0.27141f
C138 a_n3620_n557# a_n4346_n691# 0.27141f
C139 a_n3798_n557# a_n4346_n691# 0.27141f
C140 a_n3976_n557# a_n4346_n691# 0.27141f
C141 a_n4154_n557# a_n4346_n691# 0.307672f
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_4Z8MHY a_652_n562# a_n1186_n536# a_238_n536#
+ a_n1662_n562# a_3678_n562# a_n2254_n536# a_n2730_n562# a_n3322_n536# a_n60_n562#
+ a_1484_n536# a_2552_n536# a_n830_n536# a_3620_n536# w_n4412_n762# a_2076_n562# a_3144_n562#
+ a_1008_n562# a_n3678_n536# a_n416_n562# a_950_n536# a_474_n562# a_3976_n536# a_2908_n536#
+ a_n1484_n562# a_n2076_n536# a_n2552_n562# a_n3144_n536# a_n1008_n536# a_n3620_n562#
+ a_n4212_n536# a_1720_n562# a_2374_n536# a_n652_n536# a_1306_n536# a_3442_n536# a_n3976_n562#
+ a_4034_n562# a_n238_n562# a_772_n536# a_n2908_n562# a_296_n562# a_3798_n536# a_n1720_n536#
+ a_n2374_n562# a_n3442_n562# a_n1306_n562# a_n4034_n536# a_1542_n562# a_2196_n536#
+ a_n474_n536# a_2610_n562# a_n950_n562# a_1128_n536# a_3264_n536# a_n3798_n562# a_594_n536#
+ a_1898_n562# a_2966_n562# a_n1542_n536# a_n2610_n536# a_118_n562# a_n2196_n562#
+ 0 a_1840_n536# a_n3264_n562# a_n1128_n562# a_1364_n562# a_n1898_n536# a_n296_n536#
+ a_2432_n562# a_n2966_n536# a_n772_n562# a_3086_n536# a_3500_n562# a_2018_n536# a_4154_n536#
+ a_60_n536# a_830_n562# a_2788_n562# a_n1364_n536# a_416_n536# a_n1840_n562# a_3856_n562#
+ a_n2432_n536# a_n3500_n536# a_1662_n536# a_n3086_n562# a_2730_n536# a_n4154_n562#
+ a_n2018_n562# a_1186_n562# a_2254_n562# a_n2788_n536# a_n594_n562# a_3322_n562#
+ a_n3856_n536# a_n118_n536#
X0 a_2552_n536# a_2432_n562# a_2374_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X1 a_950_n536# a_830_n562# a_772_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X2 a_3620_n536# a_3500_n562# a_3442_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X3 a_n3678_n536# a_n3798_n562# a_n3856_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X4 a_n830_n536# a_n950_n562# a_n1008_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X5 a_n2076_n536# a_n2196_n562# a_n2254_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X6 a_n474_n536# a_n594_n562# a_n652_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X7 a_1840_n536# a_1720_n562# a_1662_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X8 a_416_n536# a_296_n562# a_238_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X9 a_n3500_n536# a_n3620_n562# a_n3678_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X10 a_n3144_n536# a_n3264_n562# a_n3322_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X11 a_2908_n536# a_2788_n562# a_2730_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X12 a_4154_n536# a_4034_n562# a_3976_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=0.6
X13 a_n1898_n536# a_n2018_n562# a_n2076_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X14 a_n296_n536# a_n416_n562# a_n474_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X15 a_1306_n536# a_1186_n562# a_1128_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X16 a_n1720_n536# a_n1840_n562# a_n1898_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X17 a_n1364_n536# a_n1484_n562# a_n1542_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X18 a_238_n536# a_118_n562# a_60_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X19 a_3976_n536# a_3856_n562# a_3798_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X20 a_n2788_n536# a_n2908_n562# a_n2966_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X21 a_2374_n536# a_2254_n562# a_2196_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X22 a_n2432_n536# a_n2552_n562# a_n2610_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X23 a_1128_n536# a_1008_n562# a_950_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X24 a_n1186_n536# a_n1306_n562# a_n1364_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X25 a_772_n536# a_652_n562# a_594_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X26 a_3442_n536# a_3322_n562# a_3264_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X27 a_1662_n536# a_1542_n562# a_1484_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X28 a_n2966_n536# a_n3086_n562# a_n3144_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X29 a_2730_n536# a_2610_n562# a_2552_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X30 a_n4034_n536# a_n4154_n562# a_n4212_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=0.6
X31 a_n118_n536# a_n238_n562# a_n296_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X32 a_3798_n536# a_3678_n562# a_3620_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X33 a_n3856_n536# a_n3976_n562# a_n4034_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X34 a_n2610_n536# a_n2730_n562# a_n2788_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X35 a_2196_n536# a_2076_n562# a_2018_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X36 a_n2254_n536# a_n2374_n562# a_n2432_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X37 a_n652_n536# a_n772_n562# a_n830_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X38 a_2018_n536# a_1898_n562# a_1840_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X39 a_n1008_n536# a_n1128_n562# a_n1186_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X40 a_594_n536# a_474_n562# a_416_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X41 a_3264_n536# a_3144_n562# a_3086_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X42 a_n3322_n536# a_n3442_n562# a_n3500_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X43 a_60_n536# a_n60_n562# a_n118_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X44 a_3086_n536# a_2966_n562# a_2908_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X45 a_1484_n536# a_1364_n562# a_1306_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X46 a_n1542_n536# a_n1662_n562# a_n1720_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
C0 a_n1186_n536# a_n1364_n536# 0.396241f
C1 a_n4212_n536# a_n4034_n536# 0.396241f
C2 a_n60_n562# w_n4412_n762# 0.154143f
C3 w_n4412_n762# a_n4154_n562# 0.178797f
C4 a_1720_n562# w_n4412_n762# 0.154143f
C5 w_n4412_n762# a_n2374_n562# 0.154143f
C6 a_n474_n536# a_n296_n536# 0.396241f
C7 a_n3678_n536# a_n3500_n536# 0.396241f
C8 a_n2018_n562# w_n4412_n762# 0.154143f
C9 a_4034_n562# w_n4412_n762# 0.178797f
C10 w_n4412_n762# a_n3798_n562# 0.154143f
C11 w_n4412_n762# a_n1484_n562# 0.154143f
C12 a_238_n536# a_60_n536# 0.396241f
C13 a_n2254_n536# a_n2432_n536# 0.396241f
C14 a_n3500_n536# a_n3322_n536# 0.396241f
C15 a_n1542_n536# a_n1364_n536# 0.396241f
C16 a_n2966_n536# a_n3144_n536# 0.396241f
C17 a_n2908_n562# w_n4412_n762# 0.154143f
C18 a_2908_n536# a_2730_n536# 0.396241f
C19 a_238_n536# a_416_n536# 0.396241f
C20 w_n4412_n762# a_n3442_n562# 0.154143f
C21 a_1364_n562# w_n4412_n762# 0.154143f
C22 a_n2432_n536# a_n2610_n536# 0.396241f
C23 a_3500_n562# w_n4412_n762# 0.154143f
C24 w_n4412_n762# a_1186_n562# 0.154143f
C25 a_n1306_n562# w_n4412_n762# 0.154143f
C26 a_n950_n562# w_n4412_n762# 0.154143f
C27 a_n2788_n536# a_n2610_n536# 0.396241f
C28 a_n4212_n536# w_n4412_n762# 0.306477f
C29 a_3620_n536# a_3798_n536# 0.396241f
C30 a_4154_n536# w_n4412_n762# 0.306477f
C31 a_n1662_n562# w_n4412_n762# 0.154143f
C32 a_n3086_n562# w_n4412_n762# 0.154143f
C33 a_2966_n562# w_n4412_n762# 0.154143f
C34 a_1662_n536# a_1840_n536# 0.396241f
C35 a_1128_n536# a_950_n536# 0.396241f
C36 a_2196_n536# a_2018_n536# 0.396241f
C37 a_772_n536# a_950_n536# 0.396241f
C38 a_1840_n536# a_2018_n536# 0.396241f
C39 a_n416_n562# w_n4412_n762# 0.154143f
C40 w_n4412_n762# a_1542_n562# 0.154143f
C41 a_3442_n536# a_3264_n536# 0.396241f
C42 a_3976_n536# a_4154_n536# 0.396241f
C43 a_1662_n536# a_1484_n536# 0.396241f
C44 a_1306_n536# a_1484_n536# 0.396241f
C45 a_2552_n536# a_2374_n536# 0.396241f
C46 a_2076_n562# w_n4412_n762# 0.154143f
C47 a_n830_n536# a_n652_n536# 0.396241f
C48 a_2610_n562# w_n4412_n762# 0.154143f
C49 a_n1008_n536# a_n1186_n536# 0.396241f
C50 a_3322_n562# w_n4412_n762# 0.154143f
C51 a_n474_n536# a_n652_n536# 0.396241f
C52 a_416_n536# a_594_n536# 0.396241f
C53 a_60_n536# a_n118_n536# 0.396241f
C54 w_n4412_n762# a_n3976_n562# 0.154143f
C55 a_n2196_n562# w_n4412_n762# 0.154143f
C56 a_n3264_n562# w_n4412_n762# 0.154143f
C57 a_474_n562# w_n4412_n762# 0.154143f
C58 a_3086_n536# a_3264_n536# 0.396241f
C59 a_118_n562# w_n4412_n762# 0.154143f
C60 w_n4412_n762# a_n3620_n562# 0.154143f
C61 a_n1720_n536# a_n1898_n536# 0.396241f
C62 a_n1008_n536# a_n830_n536# 0.396241f
C63 w_n4412_n762# a_652_n562# 0.154143f
C64 a_n594_n562# w_n4412_n762# 0.154143f
C65 a_3856_n562# w_n4412_n762# 0.154143f
C66 a_n3678_n536# a_n3856_n536# 0.396241f
C67 w_n4412_n762# a_296_n562# 0.154143f
C68 a_n3322_n536# a_n3144_n536# 0.396241f
C69 a_2432_n562# w_n4412_n762# 0.154143f
C70 a_n1128_n562# w_n4412_n762# 0.154143f
C71 a_n1840_n562# w_n4412_n762# 0.154143f
C72 a_n2730_n562# w_n4412_n762# 0.154143f
C73 w_n4412_n762# a_3678_n562# 0.154143f
C74 a_n772_n562# w_n4412_n762# 0.154143f
C75 a_n2966_n536# a_n2788_n536# 0.396241f
C76 w_n4412_n762# a_1898_n562# 0.154143f
C77 a_n1542_n536# a_n1720_n536# 0.396241f
C78 w_n4412_n762# a_2788_n562# 0.154143f
C79 a_830_n562# w_n4412_n762# 0.154143f
C80 a_2552_n536# a_2730_n536# 0.396241f
C81 a_3086_n536# a_2908_n536# 0.396241f
C82 a_n2076_n536# a_n2254_n536# 0.396241f
C83 a_1306_n536# a_1128_n536# 0.396241f
C84 a_3976_n536# a_3798_n536# 0.396241f
C85 w_n4412_n762# a_2254_n562# 0.154143f
C86 a_1008_n562# w_n4412_n762# 0.154143f
C87 a_2196_n536# a_2374_n536# 0.396241f
C88 a_3144_n562# w_n4412_n762# 0.154143f
C89 a_n2552_n562# w_n4412_n762# 0.154143f
C90 w_n4412_n762# a_n238_n562# 0.154143f
C91 a_n296_n536# a_n118_n536# 0.396241f
C92 a_n3856_n536# a_n4034_n536# 0.396241f
C93 a_772_n536# a_594_n536# 0.396241f
C94 a_n2076_n536# a_n1898_n536# 0.396241f
C95 a_3442_n536# a_3620_n536# 0.396241f
C96 a_4154_n536# 0 0.229314f
C97 a_3976_n536# 0 0.102508f
C98 a_3798_n536# 0 0.102508f
C99 a_3620_n536# 0 0.102508f
C100 a_3442_n536# 0 0.102508f
C101 a_3264_n536# 0 0.102508f
C102 a_3086_n536# 0 0.102508f
C103 a_2908_n536# 0 0.102508f
C104 a_2730_n536# 0 0.102508f
C105 a_2552_n536# 0 0.102508f
C106 a_2374_n536# 0 0.102508f
C107 a_2196_n536# 0 0.102508f
C108 a_2018_n536# 0 0.102508f
C109 a_1840_n536# 0 0.102508f
C110 a_1662_n536# 0 0.102508f
C111 a_1484_n536# 0 0.102508f
C112 a_1306_n536# 0 0.102508f
C113 a_1128_n536# 0 0.102508f
C114 a_950_n536# 0 0.102508f
C115 a_772_n536# 0 0.102508f
C116 a_594_n536# 0 0.102508f
C117 a_416_n536# 0 0.102508f
C118 a_238_n536# 0 0.102508f
C119 a_60_n536# 0 0.102508f
C120 a_n118_n536# 0 0.102508f
C121 a_n296_n536# 0 0.102508f
C122 a_n474_n536# 0 0.102508f
C123 a_n652_n536# 0 0.102508f
C124 a_n830_n536# 0 0.102508f
C125 a_n1008_n536# 0 0.102508f
C126 a_n1186_n536# 0 0.102508f
C127 a_n1364_n536# 0 0.102508f
C128 a_n1542_n536# 0 0.102508f
C129 a_n1720_n536# 0 0.102508f
C130 a_n1898_n536# 0 0.102508f
C131 a_n2076_n536# 0 0.102508f
C132 a_n2254_n536# 0 0.102508f
C133 a_n2432_n536# 0 0.102508f
C134 a_n2610_n536# 0 0.102508f
C135 a_n2788_n536# 0 0.102508f
C136 a_n2966_n536# 0 0.102508f
C137 a_n3144_n536# 0 0.102508f
C138 a_n3322_n536# 0 0.102508f
C139 a_n3500_n536# 0 0.102508f
C140 a_n3678_n536# 0 0.102508f
C141 a_n3856_n536# 0 0.102508f
C142 a_n4034_n536# 0 0.102508f
C143 a_n4212_n536# 0 0.229314f
C144 a_4034_n562# 0 0.135281f
C145 a_3856_n562# 0 0.1219f
C146 a_3678_n562# 0 0.1219f
C147 a_3500_n562# 0 0.1219f
C148 a_3322_n562# 0 0.1219f
C149 a_3144_n562# 0 0.1219f
C150 a_2966_n562# 0 0.1219f
C151 a_2788_n562# 0 0.1219f
C152 a_2610_n562# 0 0.1219f
C153 a_2432_n562# 0 0.1219f
C154 a_2254_n562# 0 0.1219f
C155 a_2076_n562# 0 0.1219f
C156 a_1898_n562# 0 0.1219f
C157 a_1720_n562# 0 0.1219f
C158 a_1542_n562# 0 0.1219f
C159 a_1364_n562# 0 0.1219f
C160 a_1186_n562# 0 0.1219f
C161 a_1008_n562# 0 0.1219f
C162 a_830_n562# 0 0.1219f
C163 a_652_n562# 0 0.1219f
C164 a_474_n562# 0 0.1219f
C165 a_296_n562# 0 0.1219f
C166 a_118_n562# 0 0.1219f
C167 a_n60_n562# 0 0.1219f
C168 a_n238_n562# 0 0.1219f
C169 a_n416_n562# 0 0.1219f
C170 a_n594_n562# 0 0.1219f
C171 a_n772_n562# 0 0.1219f
C172 a_n950_n562# 0 0.1219f
C173 a_n1128_n562# 0 0.1219f
C174 a_n1306_n562# 0 0.1219f
C175 a_n1484_n562# 0 0.1219f
C176 a_n1662_n562# 0 0.1219f
C177 a_n1840_n562# 0 0.1219f
C178 a_n2018_n562# 0 0.1219f
C179 a_n2196_n562# 0 0.1219f
C180 a_n2374_n562# 0 0.1219f
C181 a_n2552_n562# 0 0.1219f
C182 a_n2730_n562# 0 0.1219f
C183 a_n2908_n562# 0 0.1219f
C184 a_n3086_n562# 0 0.1219f
C185 a_n3264_n562# 0 0.1219f
C186 a_n3442_n562# 0 0.1219f
C187 a_n3620_n562# 0 0.1219f
C188 a_n3798_n562# 0 0.1219f
C189 a_n3976_n562# 0 0.1219f
C190 a_n4154_n562# 0 0.135281f
C191 w_n4412_n762# 0 46.4171f
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_WY4TLZ a_n919_n536# a_207_n562# a_n1217_n562#
+ w_n1653_n762# a_n385_n536# a_1039_n536# a_n861_n562# a_n1453_n536# a_505_n536# a_1275_n562#
+ a_29_n562# a_n1039_n562# a_n683_n562# a_n207_n536# a_741_n562# a_327_n536# a_n1275_n536#
+ a_1097_n562# a_n505_n562# a_n29_n536# a_n1097_n536# a_563_n562# a_149_n536# a_1395_n536#
+ 0 a_n741_n536# a_919_n562# a_861_n536# a_n327_n562# a_385_n562# a_n1395_n562# a_1217_n536#
+ a_n563_n536# a_683_n536# a_n149_n562#
X0 a_n207_n536# a_n327_n562# a_n385_n536# w_n1653_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X1 a_1217_n536# a_1097_n562# a_1039_n536# w_n1653_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X2 a_n1275_n536# a_n1395_n562# a_n1453_n536# w_n1653_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=0.6
X3 a_n741_n536# a_n861_n562# a_n919_n536# w_n1653_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X4 a_n1097_n536# a_n1217_n562# a_n1275_n536# w_n1653_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X5 a_683_n536# a_563_n562# a_505_n536# w_n1653_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X6 a_1039_n536# a_919_n562# a_861_n536# w_n1653_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X7 a_n29_n536# a_n149_n562# a_n207_n536# w_n1653_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X8 a_n563_n536# a_n683_n562# a_n741_n536# w_n1653_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X9 a_n919_n536# a_n1039_n562# a_n1097_n536# w_n1653_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X10 a_505_n536# a_385_n562# a_327_n536# w_n1653_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X11 a_n385_n536# a_n505_n562# a_n563_n536# w_n1653_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X12 a_1395_n536# a_1275_n562# a_1217_n536# w_n1653_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=0.6
X13 a_327_n536# a_207_n562# a_149_n536# w_n1653_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X14 a_149_n536# a_29_n562# a_n29_n536# w_n1653_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X15 a_861_n536# a_741_n562# a_683_n536# w_n1653_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
C0 a_327_n536# a_149_n536# 0.396241f
C1 a_n1217_n562# w_n1653_n762# 0.154143f
C2 a_1275_n562# w_n1653_n762# 0.178797f
C3 a_n563_n536# a_n741_n536# 0.396241f
C4 a_683_n536# a_861_n536# 0.396241f
C5 a_919_n562# w_n1653_n762# 0.154143f
C6 a_n919_n536# a_n741_n536# 0.396241f
C7 a_n29_n536# a_n207_n536# 0.396241f
C8 a_n683_n562# w_n1653_n762# 0.154143f
C9 a_n149_n562# w_n1653_n762# 0.154143f
C10 a_1039_n536# a_1217_n536# 0.396241f
C11 a_29_n562# w_n1653_n762# 0.154143f
C12 a_n1395_n562# w_n1653_n762# 0.178797f
C13 a_n563_n536# a_n385_n536# 0.396241f
C14 a_741_n562# w_n1653_n762# 0.154143f
C15 a_327_n536# a_505_n536# 0.396241f
C16 a_1395_n536# w_n1653_n762# 0.306477f
C17 a_n29_n536# a_149_n536# 0.396241f
C18 a_1097_n562# w_n1653_n762# 0.154143f
C19 a_n1453_n536# w_n1653_n762# 0.306477f
C20 a_n861_n562# w_n1653_n762# 0.154143f
C21 a_n1097_n536# a_n1275_n536# 0.396241f
C22 a_n505_n562# w_n1653_n762# 0.154143f
C23 a_n1039_n562# w_n1653_n762# 0.154143f
C24 a_1395_n536# a_1217_n536# 0.396241f
C25 a_n919_n536# a_n1097_n536# 0.396241f
C26 a_1039_n536# a_861_n536# 0.396241f
C27 a_n327_n562# w_n1653_n762# 0.154143f
C28 a_563_n562# w_n1653_n762# 0.154143f
C29 a_385_n562# w_n1653_n762# 0.154143f
C30 a_683_n536# a_505_n536# 0.396241f
C31 a_n1453_n536# a_n1275_n536# 0.396241f
C32 a_207_n562# w_n1653_n762# 0.154143f
C33 a_n385_n536# a_n207_n536# 0.396241f
C34 a_1395_n536# 0 0.229314f
C35 a_1217_n536# 0 0.102508f
C36 a_1039_n536# 0 0.102508f
C37 a_861_n536# 0 0.102508f
C38 a_683_n536# 0 0.102508f
C39 a_505_n536# 0 0.102508f
C40 a_327_n536# 0 0.102508f
C41 a_149_n536# 0 0.102508f
C42 a_n29_n536# 0 0.102508f
C43 a_n207_n536# 0 0.102508f
C44 a_n385_n536# 0 0.102508f
C45 a_n563_n536# 0 0.102508f
C46 a_n741_n536# 0 0.102508f
C47 a_n919_n536# 0 0.102508f
C48 a_n1097_n536# 0 0.102508f
C49 a_n1275_n536# 0 0.102508f
C50 a_n1453_n536# 0 0.229314f
C51 a_1275_n562# 0 0.135281f
C52 a_1097_n562# 0 0.1219f
C53 a_919_n562# 0 0.1219f
C54 a_741_n562# 0 0.1219f
C55 a_563_n562# 0 0.1219f
C56 a_385_n562# 0 0.1219f
C57 a_207_n562# 0 0.1219f
C58 a_29_n562# 0 0.1219f
C59 a_n149_n562# 0 0.1219f
C60 a_n327_n562# 0 0.1219f
C61 a_n505_n562# 0 0.1219f
C62 a_n683_n562# 0 0.1219f
C63 a_n861_n562# 0 0.1219f
C64 a_n1039_n562# 0 0.1219f
C65 a_n1217_n562# 0 0.1219f
C66 a_n1395_n562# 0 0.135281f
C67 w_n1653_n762# 0 17.7208f
.ends

.subckt sky130_fd_sc_hvl__inv_1 A VGND VNB VPB VPWR Y
X0 Y A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X1 Y A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
C0 Y VPWR 0.136398f
C1 VPWR VPB 0.245656f
C2 A Y 0.101326f
C3 A VPWR 0.114724f
C4 VGND VNB 0.303489f
C5 Y VNB 0.158366f
C6 A VNB 0.320027f
C7 VPB VNB 0.793675f
.ends

.subckt sky130_fd_pr__res_xhigh_po_1p41_9VZRJ2 a_n7134_n3916# a_n8646_3484# a_7230_3484#
+ a_n5244_3484# a_8364_n3916# a_12144_3484# a_n7512_n3916# a_6096_n3916# a_n9024_3484#
+ a_n5244_n3916# a_n12048_n3916# a_8742_n3916# a_6474_n3916# a_n330_n3916# a_n708_n3916#
+ a_n12426_n3916# a_48_n3916# a_n5622_n3916# a_n7890_3484# a_7986_3484# a_n12804_3484#
+ a_4584_3484# a_n2598_3484# a_n3354_n3916# a_n10158_n3916# a_n13182_3484# a_1182_3484#
+ a_6852_n3916# a_n12804_n3916# a_11388_n3916# a_4584_n3916# a_n1086_n3916# a_8364_3484#
+ a_n10536_n3916# a_n3732_n3916# a_n6378_3484# a_11766_n3916# a_4962_n3916# a_n1464_n3916#
+ a_n10914_n3916# a_2694_n3916# a_n1842_n3916# a_n9780_n3916# a_n1842_3484# a_1938_3484#
+ a_48_3484# a_n10536_3484# a_n5622_3484# a_5718_3484# a_9498_3484# a_n2220_3484#
+ a_n7890_n3916# a_2316_3484# a_6096_3484# a_12522_3484# a_9120_n3916# a_n9402_3484#
+ a_n6000_3484# a_n6000_n3916# a_7230_n3916# a_7608_n3916# a_426_n3916# a_4962_3484#
+ a_1560_3484# a_n2976_3484# a_804_n3916# a_n4110_n3916# a_8742_3484# a_n6756_3484#
+ a_5340_3484# a_12144_n3916# a_n3354_3484# a_5340_n3916# a_5718_n3916# a_n13312_n4046#
+ a_n12048_3484# a_10254_3484# a_3072_n3916# a_9120_3484# a_12522_n3916# a_n2220_n3916#
+ a_n7134_3484# a_426_3484# a_10254_n3916# a_3450_n3916# a_3828_n3916# a_12900_n3916#
+ a_n708_3484# a_1182_n3916# a_n8268_n3916# a_10632_n3916# a_n10914_3484# a_2694_3484#
+ a_n11292_3484# a_9498_n3916# a_n8646_n3916# a_n9780_3484# a_1560_n3916# a_1938_n3916#
+ a_9876_3484# a_6474_3484# a_12900_3484# a_n4488_3484# a_3072_3484# a_9876_n3916#
+ a_n1086_3484# a_n6378_n3916# a_11388_3484# a_n8268_3484# a_n13182_n3916# a_n6756_n3916#
+ a_n330_3484# a_7986_n3916# a_n4488_n3916# a_n11292_n3916# a_n4866_n3916# a_n2598_n3916#
+ a_n3732_3484# a_3828_3484# a_n11670_n3916# a_n12426_3484# a_10632_3484# a_n2976_n3916#
+ a_n7512_3484# a_7608_3484# a_804_3484# a_n4110_3484# a_4206_3484# a_4206_n3916#
+ a_11010_3484# a_11010_n3916# a_n11670_3484# a_2316_n3916# a_n9024_n3916# a_6852_3484#
+ a_3450_3484# a_n4866_3484# a_n9402_n3916# a_n1464_3484# a_n10158_3484# a_11766_3484#
X0 a_n9024_3484# a_n9024_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X1 a_9876_3484# a_9876_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X2 a_n11670_3484# a_n11670_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X3 a_n330_3484# a_n330_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X4 a_3072_3484# a_3072_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X5 a_5718_3484# a_5718_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X6 a_6474_3484# a_6474_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X7 a_8742_3484# a_8742_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X8 a_n11292_3484# a_n11292_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X9 a_n10536_3484# a_n10536_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X10 a_n7890_3484# a_n7890_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X11 a_2316_3484# a_2316_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X12 a_5340_3484# a_5340_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X13 a_n12804_3484# a_n12804_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X14 a_n6756_3484# a_n6756_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X15 a_n4488_3484# a_n4488_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X16 a_n1086_3484# a_n1086_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X17 a_12144_3484# a_12144_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X18 a_n5622_3484# a_n5622_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X19 a_n3354_3484# a_n3354_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X20 a_11010_3484# a_11010_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X21 a_6096_3484# a_6096_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X22 a_9498_3484# a_9498_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X23 a_7608_3484# a_7608_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X24 a_8364_3484# a_8364_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X25 a_n13182_3484# a_n13182_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X26 a_n10158_3484# a_n10158_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X27 a_n9780_3484# a_n9780_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X28 a_4206_3484# a_4206_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X29 a_7230_3484# a_7230_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X30 a_n12426_3484# a_n12426_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X31 a_n8646_3484# a_n8646_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X32 a_n6378_3484# a_n6378_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X33 a_n7512_3484# a_n7512_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X34 a_n5244_3484# a_n5244_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X35 a_n2220_3484# a_n2220_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X36 a_1938_3484# a_1938_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X37 a_2694_3484# a_2694_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X38 a_4962_3484# a_4962_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X39 a_1560_3484# a_1560_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X40 a_11766_3484# a_11766_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X41 a_n2976_3484# a_n2976_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X42 a_48_3484# a_48_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X43 a_10632_3484# a_10632_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X44 a_12900_3484# a_12900_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X45 a_n1842_3484# a_n1842_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X46 a_804_3484# a_804_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X47 a_9120_3484# a_9120_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X48 a_n12048_3484# a_n12048_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X49 a_n8268_3484# a_n8268_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X50 a_n7134_3484# a_n7134_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X51 a_n4110_3484# a_n4110_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X52 a_7986_3484# a_7986_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X53 a_n9402_3484# a_n9402_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X54 a_4584_3484# a_4584_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X55 a_n6000_3484# a_n6000_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X56 a_n708_3484# a_n708_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X57 a_1182_3484# a_1182_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X58 a_3828_3484# a_3828_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X59 a_6852_3484# a_6852_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X60 a_11388_3484# a_11388_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X61 a_n2598_3484# a_n2598_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X62 a_3450_3484# a_3450_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X63 a_10254_3484# a_10254_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X64 a_n10914_3484# a_n10914_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X65 a_n4866_3484# a_n4866_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X66 a_12522_3484# a_12522_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X67 a_n3732_3484# a_n3732_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X68 a_n1464_3484# a_n1464_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X69 a_426_3484# a_426_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
C0 a_12144_n3916# a_12522_n3916# 0.296258f
C1 a_n7134_3484# a_n6756_3484# 0.296258f
C2 a_10632_3484# a_11010_3484# 0.296258f
C3 a_n12426_n3916# a_n12048_n3916# 0.296258f
C4 a_1560_n3916# a_1182_n3916# 0.296258f
C5 a_n11670_n3916# a_n12048_n3916# 0.296258f
C6 a_4206_3484# a_4584_3484# 0.296258f
C7 a_n708_n3916# a_n330_n3916# 0.296258f
C8 a_7986_3484# a_8364_3484# 0.296258f
C9 a_n708_3484# a_n1086_3484# 0.296258f
C10 a_3450_3484# a_3828_3484# 0.296258f
C11 a_n9402_3484# a_n9780_3484# 0.296258f
C12 a_n1842_3484# a_n1464_3484# 0.296258f
C13 a_n1842_3484# a_n2220_3484# 0.296258f
C14 a_n12804_3484# a_n13182_3484# 0.296258f
C15 a_6474_n3916# a_6852_n3916# 0.296258f
C16 a_n8646_3484# a_n9024_3484# 0.296258f
C17 a_n5622_3484# a_n5244_3484# 0.296258f
C18 a_n6000_3484# a_n6378_3484# 0.296258f
C19 a_10632_n3916# a_11010_n3916# 0.296258f
C20 a_7608_3484# a_7986_3484# 0.296258f
C21 a_3072_3484# a_3450_3484# 0.296258f
C22 a_n6000_n3916# a_n6378_n3916# 0.296258f
C23 a_n5244_3484# a_n4866_3484# 0.296258f
C24 a_9120_n3916# a_9498_n3916# 0.296258f
C25 a_n8268_n3916# a_n8646_n3916# 0.296258f
C26 a_n4110_3484# a_n4488_3484# 0.296258f
C27 a_6096_n3916# a_6474_n3916# 0.296258f
C28 a_n4866_n3916# a_n4488_n3916# 0.296258f
C29 a_n10536_3484# a_n10914_3484# 0.296258f
C30 a_11010_3484# a_11388_3484# 0.296258f
C31 a_n7890_3484# a_n7512_3484# 0.296258f
C32 a_n1464_n3916# a_n1086_n3916# 0.296258f
C33 a_6096_n3916# a_5718_n3916# 0.296258f
C34 a_3450_n3916# a_3828_n3916# 0.296258f
C35 a_n11292_n3916# a_n10914_n3916# 0.296258f
C36 a_9498_3484# a_9876_3484# 0.296258f
C37 a_n12804_n3916# a_n13182_n3916# 0.296258f
C38 a_48_n3916# a_426_n3916# 0.296258f
C39 a_7230_3484# a_7608_3484# 0.296258f
C40 a_5340_n3916# a_5718_n3916# 0.296258f
C41 a_1938_n3916# a_2316_n3916# 0.296258f
C42 a_n2598_3484# a_n2976_3484# 0.296258f
C43 a_n9780_3484# a_n10158_3484# 0.296258f
C44 a_n9402_n3916# a_n9024_n3916# 0.296258f
C45 a_n4110_n3916# a_n3732_n3916# 0.296258f
C46 a_11010_n3916# a_11388_n3916# 0.296258f
C47 a_804_3484# a_1182_3484# 0.296258f
C48 a_n2220_3484# a_n2598_3484# 0.296258f
C49 a_6852_3484# a_7230_3484# 0.296258f
C50 a_n1464_3484# a_n1086_3484# 0.296258f
C51 a_n10536_n3916# a_n10914_n3916# 0.296258f
C52 a_4962_n3916# a_5340_n3916# 0.296258f
C53 a_8364_n3916# a_8742_n3916# 0.296258f
C54 a_1560_n3916# a_1938_n3916# 0.296258f
C55 a_1560_3484# a_1182_3484# 0.296258f
C56 a_11388_3484# a_11766_3484# 0.296258f
C57 a_n11670_3484# a_n12048_3484# 0.296258f
C58 a_n1842_n3916# a_n2220_n3916# 0.296258f
C59 a_n1842_n3916# a_n1464_n3916# 0.296258f
C60 a_n6756_3484# a_n6378_3484# 0.296258f
C61 a_48_n3916# a_n330_n3916# 0.296258f
C62 a_n11292_3484# a_n11670_3484# 0.296258f
C63 a_6474_3484# a_6852_3484# 0.296258f
C64 a_n10536_n3916# a_n10158_n3916# 0.296258f
C65 a_n8268_3484# a_n7890_3484# 0.296258f
C66 a_n3732_3484# a_n3354_3484# 0.296258f
C67 a_4584_n3916# a_4962_n3916# 0.296258f
C68 a_9498_n3916# a_9876_n3916# 0.296258f
C69 a_n5244_n3916# a_n5622_n3916# 0.296258f
C70 a_6474_3484# a_6096_3484# 0.296258f
C71 a_3828_3484# a_4206_3484# 0.296258f
C72 a_n10536_3484# a_n10158_3484# 0.296258f
C73 a_n708_3484# a_n330_3484# 0.296258f
C74 a_12900_3484# a_12522_3484# 0.296258f
C75 a_48_3484# a_n330_3484# 0.296258f
C76 a_11388_n3916# a_11766_n3916# 0.296258f
C77 a_5718_3484# a_6096_3484# 0.296258f
C78 a_n3732_n3916# a_n3354_n3916# 0.296258f
C79 a_2694_n3916# a_2316_n3916# 0.296258f
C80 a_n1086_n3916# a_n708_n3916# 0.296258f
C81 a_9876_3484# a_10254_3484# 0.296258f
C82 a_n9402_3484# a_n9024_3484# 0.296258f
C83 a_8742_3484# a_9120_3484# 0.296258f
C84 a_2316_3484# a_2694_3484# 0.296258f
C85 a_n12048_3484# a_n12426_3484# 0.296258f
C86 a_n2976_n3916# a_n2598_n3916# 0.296258f
C87 a_n6000_n3916# a_n5622_n3916# 0.296258f
C88 a_426_n3916# a_804_n3916# 0.296258f
C89 a_n7890_n3916# a_n7512_n3916# 0.296258f
C90 a_4206_n3916# a_4584_n3916# 0.296258f
C91 a_804_n3916# a_1182_n3916# 0.296258f
C92 a_7986_n3916# a_8364_n3916# 0.296258f
C93 a_11766_3484# a_12144_3484# 0.296258f
C94 a_n6000_3484# a_n5622_3484# 0.296258f
C95 a_n10158_n3916# a_n9780_n3916# 0.296258f
C96 a_n6378_n3916# a_n6756_n3916# 0.296258f
C97 a_n12804_3484# a_n12426_3484# 0.296258f
C98 a_n2976_n3916# a_n3354_n3916# 0.296258f
C99 a_48_3484# a_426_3484# 0.296258f
C100 a_426_3484# a_804_3484# 0.296258f
C101 a_5340_3484# a_5718_3484# 0.296258f
C102 a_12900_n3916# a_12522_n3916# 0.296258f
C103 a_n7890_n3916# a_n8268_n3916# 0.296258f
C104 a_1938_3484# a_2316_3484# 0.296258f
C105 a_9876_n3916# a_10254_n3916# 0.296258f
C106 a_n7134_3484# a_n7512_3484# 0.296258f
C107 a_n3354_3484# a_n2976_3484# 0.296258f
C108 a_3828_n3916# a_4206_n3916# 0.296258f
C109 a_7608_n3916# a_7986_n3916# 0.296258f
C110 a_3072_n3916# a_3450_n3916# 0.296258f
C111 a_11766_n3916# a_12144_n3916# 0.296258f
C112 a_10254_3484# a_10632_3484# 0.296258f
C113 a_4962_3484# a_5340_3484# 0.296258f
C114 a_n8646_n3916# a_n9024_n3916# 0.296258f
C115 a_n5244_n3916# a_n4866_n3916# 0.296258f
C116 a_1560_3484# a_1938_3484# 0.296258f
C117 a_8742_n3916# a_9120_n3916# 0.296258f
C118 a_n9402_n3916# a_n9780_n3916# 0.296258f
C119 a_12144_3484# a_12522_3484# 0.296258f
C120 a_n4488_3484# a_n4866_3484# 0.296258f
C121 a_7230_n3916# a_7608_n3916# 0.296258f
C122 a_2694_n3916# a_3072_n3916# 0.296258f
C123 a_n8268_3484# a_n8646_3484# 0.296258f
C124 a_n2220_n3916# a_n2598_n3916# 0.296258f
C125 a_3072_3484# a_2694_3484# 0.296258f
C126 a_4584_3484# a_4962_3484# 0.296258f
C127 a_n7134_n3916# a_n6756_n3916# 0.296258f
C128 a_9120_3484# a_9498_3484# 0.296258f
C129 a_n11670_n3916# a_n11292_n3916# 0.296258f
C130 a_8364_3484# a_8742_3484# 0.296258f
C131 a_10254_n3916# a_10632_n3916# 0.296258f
C132 a_n7134_n3916# a_n7512_n3916# 0.296258f
C133 a_n4110_n3916# a_n4488_n3916# 0.296258f
C134 a_n12426_n3916# a_n12804_n3916# 0.296258f
C135 a_n11292_3484# a_n10914_3484# 0.296258f
C136 a_n3732_3484# a_n4110_3484# 0.296258f
C137 a_6852_n3916# a_7230_n3916# 0.296258f
C138 a_12900_n3916# a_n13312_n4046# 0.62945f
C139 a_12900_3484# a_n13312_n4046# 0.62945f
C140 a_12522_n3916# a_n13312_n4046# 0.419137f
C141 a_12522_3484# a_n13312_n4046# 0.419137f
C142 a_12144_n3916# a_n13312_n4046# 0.419137f
C143 a_12144_3484# a_n13312_n4046# 0.419137f
C144 a_11766_n3916# a_n13312_n4046# 0.419137f
C145 a_11766_3484# a_n13312_n4046# 0.419137f
C146 a_11388_n3916# a_n13312_n4046# 0.419137f
C147 a_11388_3484# a_n13312_n4046# 0.419137f
C148 a_11010_n3916# a_n13312_n4046# 0.419137f
C149 a_11010_3484# a_n13312_n4046# 0.419137f
C150 a_10632_n3916# a_n13312_n4046# 0.419137f
C151 a_10632_3484# a_n13312_n4046# 0.419137f
C152 a_10254_n3916# a_n13312_n4046# 0.419137f
C153 a_10254_3484# a_n13312_n4046# 0.419137f
C154 a_9876_n3916# a_n13312_n4046# 0.419137f
C155 a_9876_3484# a_n13312_n4046# 0.419137f
C156 a_9498_n3916# a_n13312_n4046# 0.419137f
C157 a_9498_3484# a_n13312_n4046# 0.419137f
C158 a_9120_n3916# a_n13312_n4046# 0.419137f
C159 a_9120_3484# a_n13312_n4046# 0.419137f
C160 a_8742_n3916# a_n13312_n4046# 0.419137f
C161 a_8742_3484# a_n13312_n4046# 0.419137f
C162 a_8364_n3916# a_n13312_n4046# 0.419137f
C163 a_8364_3484# a_n13312_n4046# 0.419137f
C164 a_7986_n3916# a_n13312_n4046# 0.419137f
C165 a_7986_3484# a_n13312_n4046# 0.419137f
C166 a_7608_n3916# a_n13312_n4046# 0.419137f
C167 a_7608_3484# a_n13312_n4046# 0.419137f
C168 a_7230_n3916# a_n13312_n4046# 0.419137f
C169 a_7230_3484# a_n13312_n4046# 0.419137f
C170 a_6852_n3916# a_n13312_n4046# 0.419137f
C171 a_6852_3484# a_n13312_n4046# 0.419137f
C172 a_6474_n3916# a_n13312_n4046# 0.419137f
C173 a_6474_3484# a_n13312_n4046# 0.419137f
C174 a_6096_n3916# a_n13312_n4046# 0.419137f
C175 a_6096_3484# a_n13312_n4046# 0.419137f
C176 a_5718_n3916# a_n13312_n4046# 0.419137f
C177 a_5718_3484# a_n13312_n4046# 0.419137f
C178 a_5340_n3916# a_n13312_n4046# 0.419137f
C179 a_5340_3484# a_n13312_n4046# 0.419137f
C180 a_4962_n3916# a_n13312_n4046# 0.419137f
C181 a_4962_3484# a_n13312_n4046# 0.419137f
C182 a_4584_n3916# a_n13312_n4046# 0.419137f
C183 a_4584_3484# a_n13312_n4046# 0.419137f
C184 a_4206_n3916# a_n13312_n4046# 0.419137f
C185 a_4206_3484# a_n13312_n4046# 0.419137f
C186 a_3828_n3916# a_n13312_n4046# 0.419137f
C187 a_3828_3484# a_n13312_n4046# 0.419137f
C188 a_3450_n3916# a_n13312_n4046# 0.419137f
C189 a_3450_3484# a_n13312_n4046# 0.419137f
C190 a_3072_n3916# a_n13312_n4046# 0.419137f
C191 a_3072_3484# a_n13312_n4046# 0.419137f
C192 a_2694_n3916# a_n13312_n4046# 0.419137f
C193 a_2694_3484# a_n13312_n4046# 0.419137f
C194 a_2316_n3916# a_n13312_n4046# 0.419137f
C195 a_2316_3484# a_n13312_n4046# 0.419137f
C196 a_1938_n3916# a_n13312_n4046# 0.419137f
C197 a_1938_3484# a_n13312_n4046# 0.419137f
C198 a_1560_n3916# a_n13312_n4046# 0.419137f
C199 a_1560_3484# a_n13312_n4046# 0.419137f
C200 a_1182_n3916# a_n13312_n4046# 0.419137f
C201 a_1182_3484# a_n13312_n4046# 0.419137f
C202 a_804_n3916# a_n13312_n4046# 0.419137f
C203 a_804_3484# a_n13312_n4046# 0.419137f
C204 a_426_n3916# a_n13312_n4046# 0.419137f
C205 a_426_3484# a_n13312_n4046# 0.419137f
C206 a_48_n3916# a_n13312_n4046# 0.419137f
C207 a_48_3484# a_n13312_n4046# 0.419137f
C208 a_n330_n3916# a_n13312_n4046# 0.419137f
C209 a_n330_3484# a_n13312_n4046# 0.419137f
C210 a_n708_n3916# a_n13312_n4046# 0.419137f
C211 a_n708_3484# a_n13312_n4046# 0.419137f
C212 a_n1086_n3916# a_n13312_n4046# 0.419137f
C213 a_n1086_3484# a_n13312_n4046# 0.419137f
C214 a_n1464_n3916# a_n13312_n4046# 0.419137f
C215 a_n1464_3484# a_n13312_n4046# 0.419137f
C216 a_n1842_n3916# a_n13312_n4046# 0.419137f
C217 a_n1842_3484# a_n13312_n4046# 0.419137f
C218 a_n2220_n3916# a_n13312_n4046# 0.419137f
C219 a_n2220_3484# a_n13312_n4046# 0.419137f
C220 a_n2598_n3916# a_n13312_n4046# 0.419137f
C221 a_n2598_3484# a_n13312_n4046# 0.419137f
C222 a_n2976_n3916# a_n13312_n4046# 0.419137f
C223 a_n2976_3484# a_n13312_n4046# 0.419137f
C224 a_n3354_n3916# a_n13312_n4046# 0.419137f
C225 a_n3354_3484# a_n13312_n4046# 0.419137f
C226 a_n3732_n3916# a_n13312_n4046# 0.419137f
C227 a_n3732_3484# a_n13312_n4046# 0.419137f
C228 a_n4110_n3916# a_n13312_n4046# 0.419137f
C229 a_n4110_3484# a_n13312_n4046# 0.419137f
C230 a_n4488_n3916# a_n13312_n4046# 0.419137f
C231 a_n4488_3484# a_n13312_n4046# 0.419137f
C232 a_n4866_n3916# a_n13312_n4046# 0.419137f
C233 a_n4866_3484# a_n13312_n4046# 0.419137f
C234 a_n5244_n3916# a_n13312_n4046# 0.419137f
C235 a_n5244_3484# a_n13312_n4046# 0.419137f
C236 a_n5622_n3916# a_n13312_n4046# 0.419137f
C237 a_n5622_3484# a_n13312_n4046# 0.419137f
C238 a_n6000_n3916# a_n13312_n4046# 0.419137f
C239 a_n6000_3484# a_n13312_n4046# 0.419137f
C240 a_n6378_n3916# a_n13312_n4046# 0.419137f
C241 a_n6378_3484# a_n13312_n4046# 0.419137f
C242 a_n6756_n3916# a_n13312_n4046# 0.419137f
C243 a_n6756_3484# a_n13312_n4046# 0.419137f
C244 a_n7134_n3916# a_n13312_n4046# 0.419137f
C245 a_n7134_3484# a_n13312_n4046# 0.419137f
C246 a_n7512_n3916# a_n13312_n4046# 0.419137f
C247 a_n7512_3484# a_n13312_n4046# 0.419137f
C248 a_n7890_n3916# a_n13312_n4046# 0.419137f
C249 a_n7890_3484# a_n13312_n4046# 0.419137f
C250 a_n8268_n3916# a_n13312_n4046# 0.419137f
C251 a_n8268_3484# a_n13312_n4046# 0.419137f
C252 a_n8646_n3916# a_n13312_n4046# 0.419137f
C253 a_n8646_3484# a_n13312_n4046# 0.419137f
C254 a_n9024_n3916# a_n13312_n4046# 0.419137f
C255 a_n9024_3484# a_n13312_n4046# 0.419137f
C256 a_n9402_n3916# a_n13312_n4046# 0.419137f
C257 a_n9402_3484# a_n13312_n4046# 0.419137f
C258 a_n9780_n3916# a_n13312_n4046# 0.419137f
C259 a_n9780_3484# a_n13312_n4046# 0.419137f
C260 a_n10158_n3916# a_n13312_n4046# 0.419137f
C261 a_n10158_3484# a_n13312_n4046# 0.419137f
C262 a_n10536_n3916# a_n13312_n4046# 0.419137f
C263 a_n10536_3484# a_n13312_n4046# 0.419137f
C264 a_n10914_n3916# a_n13312_n4046# 0.419137f
C265 a_n10914_3484# a_n13312_n4046# 0.419137f
C266 a_n11292_n3916# a_n13312_n4046# 0.419137f
C267 a_n11292_3484# a_n13312_n4046# 0.419137f
C268 a_n11670_n3916# a_n13312_n4046# 0.419137f
C269 a_n11670_3484# a_n13312_n4046# 0.419137f
C270 a_n12048_n3916# a_n13312_n4046# 0.419137f
C271 a_n12048_3484# a_n13312_n4046# 0.419137f
C272 a_n12426_n3916# a_n13312_n4046# 0.419137f
C273 a_n12426_3484# a_n13312_n4046# 0.419137f
C274 a_n12804_n3916# a_n13312_n4046# 0.419137f
C275 a_n12804_3484# a_n13312_n4046# 0.419137f
C276 a_n13182_n3916# a_n13312_n4046# 0.62945f
C277 a_n13182_3484# a_n13312_n4046# 0.62945f
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_CD9S2Z a_100_n100# a_n292_n322# a_n158_n100#
+ a_n100_n188#
X0 a_100_n100# a_n100_n188# a_n158_n100# a_n292_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
C0 a_100_n100# a_n292_n322# 0.137447f
C1 a_n158_n100# a_n292_n322# 0.137447f
C2 a_n100_n188# a_n292_n322# 0.688242f
.ends

.subckt rstring_mux vout_brout ena otrip_decoded_avdd[7] otrip_decoded_avdd[6] otrip_decoded_avdd[3]
+ otrip_decoded_avdd[1] m1_10352_4059# m1_24716_4059# m1_10730_n3340# m1_6572_4059#
+ m1_12998_n3340# m1_25850_n3340# m1_12242_n3340# m1_12620_4059# m1_3548_4059# m1_8840_4059#
+ m1_23204_4059# m1_6194_n3340# vtrip_decoded_avdd[3] m1_5060_4059# m1_13376_4059#
+ m1_22826_n3340# m1_20558_n3340# vtrip_decoded_avdd[1] vtrip_decoded_b_avdd[0] m1_902_n3340#
+ m1_17156_4059# m1_2036_4059# m1_19046_n3340# vtrip7 ena_b m1_24338_n3340# vtrip5
+ m1_2414_n3340# vtop m1_11864_4059# m1_21692_4059# m1_7706_n3340# m1_8084_4059# otrip_decoded_avdd[2]
+ otrip_decoded_avdd[4] otrip_decoded_avdd[0] m1_21314_n3340# m1_9218_n3340# vout_vunder
+ m1_7328_4059# m1_11486_n3340# m1_19802_n3340# m1_1658_n3340# vtrip0 vtrip_decoded_avdd[5]
+ m1_17534_n3340# vtrip_decoded_avdd[7] vtrip2 vtrip4 m1_4304_4059# vtrip6 m1_9596_4059#
+ m1_4682_n3340# m1_3170_n3340# vtrip_decoded_avdd[2] vtrip_decoded_avdd[4] m1_25472_4059#
+ vtrip_decoded_avdd[6] vtrip3 m1_5816_4059# m1_22070_n3340# avdd vtrip_decoded_b_avdd[7]
+ vtrip_decoded_avdd[0] otrip_decoded_avdd[5] vtrip1 avss
Xsky130_fd_pr__nfet_g5v0d10v5_K8JYEQ_0 vout_brout vtrip_decoded_avdd[0] vout_vunder
+ otrip_decoded_avdd[3] vtrip7 vtrip5 otrip_decoded_avdd[5] otrip_decoded_avdd[1]
+ vout_brout vout_brout avss avss otrip_decoded_avdd[6] vout_brout vout_brout vtrip6
+ vtrip4 vtrip2 vout_brout vtrip_decoded_avdd[3] avss vtrip_decoded_avdd[5] vtrip1
+ vtrip_decoded_avdd[0] vout_vunder vout_brout avss avss avss vtrip_decoded_avdd[2]
+ vtrip_decoded_avdd[6] vtrip_decoded_avdd[4] otrip_decoded_avdd[6] vout_vunder vout_brout
+ vtrip0 vout_vunder vout_vunder vtrip_decoded_avdd[1] vtrip_decoded_avdd[7] vtrip_decoded_avdd[5]
+ otrip_decoded_avdd[4] vout_vunder vout_brout vout_brout otrip_decoded_avdd[2] vtrip_decoded_avdd[4]
+ vtrip_decoded_avdd[2] avss otrip_decoded_avdd[4] otrip_decoded_avdd[0] vtrip3 vtrip_decoded_avdd[6]
+ vout_vunder vtrip7 vtrip4 vtrip2 vout_vunder vout_vunder vout_vunder vtrip_decoded_avdd[1]
+ avss avss avss vtrip5 avss vout_vunder vtrip3 vout_vunder vtrip1 avss avss avss
+ vout_vunder otrip_decoded_avdd[7] vout_brout vout_brout avss vout_brout otrip_decoded_avdd[5]
+ otrip_decoded_avdd[3] otrip_decoded_avdd[1] vtrip0 vout_brout vout_brout vtrip_decoded_avdd[3]
+ vout_brout avss vout_vunder vout_vunder vtrip6 vtrip_decoded_avdd[7] otrip_decoded_avdd[0]
+ vout_vunder otrip_decoded_avdd[7] otrip_decoded_avdd[2] sky130_fd_pr__nfet_g5v0d10v5_K8JYEQ
Xsky130_fd_pr__pfet_g5v0d10v5_4Z8MHY_0 vtrip_decoded_b_avdd[1] vout_brout vtrip0 avdd
+ avdd vout_brout avdd vout_brout avdd vout_vunder vout_vunder vtrip6 vout_vunder
+ avdd avdd avdd avdd vout_brout otrip_decoded_b_avdd[7] vout_vunder avdd vtrip7 vtrip5
+ otrip_decoded_b_avdd[5] vout_brout otrip_decoded_b_avdd[3] vout_brout vout_brout
+ otrip_decoded_b_avdd[1] vout_brout vtrip_decoded_b_avdd[3] vtrip4 vout_brout vtrip2
+ vtrip6 otrip_decoded_b_avdd[0] vtrip_decoded_b_avdd[7] otrip_decoded_b_avdd[7] vtrip1
+ otrip_decoded_b_avdd[2] vtrip_decoded_b_avdd[0] vout_vunder vout_brout otrip_decoded_b_avdd[3]
+ otrip_decoded_b_avdd[1] otrip_decoded_b_avdd[5] vtrip0 avdd vout_vunder vout_brout
+ avdd otrip_decoded_b_avdd[6] vout_vunder vout_vunder avdd vout_vunder vtrip_decoded_b_avdd[3]
+ vtrip_decoded_b_avdd[5] vout_brout vout_brout vtrip_decoded_b_avdd[0] avdd avss
+ vtrip3 avdd avdd vtrip_decoded_b_avdd[2] vtrip4 vtrip7 vtrip_decoded_b_avdd[4] vtrip2
+ otrip_decoded_b_avdd[6] vout_vunder vtrip_decoded_b_avdd[6] vout_vunder vout_vunder
+ vout_vunder vtrip_decoded_b_avdd[1] vtrip_decoded_b_avdd[5] vtrip5 vout_vunder otrip_decoded_b_avdd[4]
+ vtrip_decoded_b_avdd[7] vtrip3 vtrip1 vout_vunder otrip_decoded_b_avdd[2] vout_vunder
+ otrip_decoded_b_avdd[0] otrip_decoded_b_avdd[4] vtrip_decoded_b_avdd[2] vtrip_decoded_b_avdd[4]
+ vout_brout avdd vtrip_decoded_b_avdd[6] vout_brout vout_brout sky130_fd_pr__pfet_g5v0d10v5_4Z8MHY
Xsky130_fd_pr__pfet_g5v0d10v5_WY4TLZ_0 vtop ena_b ena_b avdd avdd avdd ena_b avdd
+ vtop ena_b ena_b ena_b ena_b vtop ena_b avdd vtop ena_b ena_b avdd avdd ena_b vtop
+ avdd avss avdd ena_b vtop ena_b ena_b ena_b vtop vtop avdd ena_b sky130_fd_pr__pfet_g5v0d10v5_WY4TLZ
Xsky130_fd_sc_hvl__inv_1_0[0] otrip_decoded_avdd[0] avss avss avdd avdd otrip_decoded_b_avdd[0]
+ sky130_fd_sc_hvl__inv_1
Xsky130_fd_sc_hvl__inv_1_0[1] otrip_decoded_avdd[1] avss avss avdd avdd otrip_decoded_b_avdd[1]
+ sky130_fd_sc_hvl__inv_1
Xsky130_fd_sc_hvl__inv_1_0[2] otrip_decoded_avdd[2] avss avss avdd avdd otrip_decoded_b_avdd[2]
+ sky130_fd_sc_hvl__inv_1
Xsky130_fd_sc_hvl__inv_1_0[3] otrip_decoded_avdd[3] avss avss avdd avdd otrip_decoded_b_avdd[3]
+ sky130_fd_sc_hvl__inv_1
Xsky130_fd_sc_hvl__inv_1_0[4] otrip_decoded_avdd[4] avss avss avdd avdd otrip_decoded_b_avdd[4]
+ sky130_fd_sc_hvl__inv_1
Xsky130_fd_sc_hvl__inv_1_0[5] otrip_decoded_avdd[5] avss avss avdd avdd otrip_decoded_b_avdd[5]
+ sky130_fd_sc_hvl__inv_1
Xsky130_fd_sc_hvl__inv_1_0[6] otrip_decoded_avdd[6] avss avss avdd avdd otrip_decoded_b_avdd[6]
+ sky130_fd_sc_hvl__inv_1
Xsky130_fd_sc_hvl__inv_1_0[7] otrip_decoded_avdd[7] avss avss avdd avdd otrip_decoded_b_avdd[7]
+ sky130_fd_sc_hvl__inv_1
Xsky130_fd_sc_hvl__inv_1_0[8] vtrip_decoded_avdd[0] avss avss avdd avdd vtrip_decoded_b_avdd[0]
+ sky130_fd_sc_hvl__inv_1
Xsky130_fd_sc_hvl__inv_1_0[9] vtrip_decoded_avdd[1] avss avss avdd avdd vtrip_decoded_b_avdd[1]
+ sky130_fd_sc_hvl__inv_1
Xsky130_fd_sc_hvl__inv_1_0[10] vtrip_decoded_avdd[2] avss avss avdd avdd vtrip_decoded_b_avdd[2]
+ sky130_fd_sc_hvl__inv_1
Xsky130_fd_sc_hvl__inv_1_0[11] vtrip_decoded_avdd[3] avss avss avdd avdd vtrip_decoded_b_avdd[3]
+ sky130_fd_sc_hvl__inv_1
Xsky130_fd_sc_hvl__inv_1_0[12] vtrip_decoded_avdd[4] avss avss avdd avdd vtrip_decoded_b_avdd[4]
+ sky130_fd_sc_hvl__inv_1
Xsky130_fd_sc_hvl__inv_1_0[13] vtrip_decoded_avdd[5] avss avss avdd avdd vtrip_decoded_b_avdd[5]
+ sky130_fd_sc_hvl__inv_1
Xsky130_fd_sc_hvl__inv_1_0[14] vtrip_decoded_avdd[6] avss avss avdd avdd vtrip_decoded_b_avdd[6]
+ sky130_fd_sc_hvl__inv_1
Xsky130_fd_sc_hvl__inv_1_0[15] vtrip_decoded_avdd[7] avss avss avdd avdd vtrip_decoded_b_avdd[7]
+ sky130_fd_sc_hvl__inv_1
Xsky130_fd_sc_hvl__inv_1_1 ena avss avss avdd avdd ena_b sky130_fd_sc_hvl__inv_1
Xsky130_fd_pr__res_xhigh_po_1p41_9VZRJ2_0 m1_6950_n3340# m1_5060_4059# m1_20936_4059#
+ m1_8840_4059# m1_22070_n3340# m1_26228_4059# m1_6194_n3340# m1_19802_n3340# m1_5060_4059#
+ m1_8462_n3340# m1_1658_n3340# m1_22826_n3340# m1_20558_n3340# vtrip0 m1_12998_n3340#
+ m1_1658_n3340# vtrip0 m1_8462_n3340# m1_5816_4059# m1_21692_4059# m1_1280_4059#
+ m1_18668_4059# m1_11108_4059# m1_10730_n3340# m1_3926_n3340# vtop vtrip3 m1_20558_n3340#
+ m1_902_n3340# m1_25094_n3340# m1_18290_n3340# m1_12998_n3340# m1_22448_4059# m1_3170_n3340#
+ m1_9974_n3340# m1_7328_4059# m1_25850_n3340# m1_19046_n3340# m1_12242_n3340# m1_3170_n3340#
+ m1_16778_n3340# m1_12242_n3340# m1_3926_n3340# m1_11864_4059# vtrip5 vtrip1 m1_3548_4059#
+ m1_8084_4059# m1_19424_4059# m1_23204_4059# m1_11864_4059# m1_6194_n3340# vtrip7
+ m1_20180_4059# m1_26228_4059# m1_22826_n3340# m1_4304_4059# m1_8084_4059# m1_7706_n3340#
+ m1_21314_n3340# m1_21314_n3340# vtrip2 m1_18668_4059# vtrip5 m1_11108_4059# vtrip2
+ m1_9974_n3340# m1_22448_4059# m1_7328_4059# m1_19424_4059# m1_25850_n3340# m1_10352_4059#
+ m1_19046_n3340# m1_19802_n3340# avss m1_2036_4059# m1_23960_4059# m1_16778_n3340#
+ m1_23204_4059# m1_26606_n3340# m1_11486_n3340# m1_6572_4059# vtrip1 m1_24338_n3340#
+ m1_17534_n3340# m1_17534_n3340# m1_26606_n3340# m1_13376_4059# vtrip4 m1_5438_n3340#
+ m1_24338_n3340# m1_2792_4059# vtrip7 m1_2792_4059# m1_23582_n3340# m1_5438_n3340#
+ m1_4304_4059# vtrip4 vtrip6 m1_23960_4059# m1_20180_4059# avss m1_9596_4059# m1_17156_4059#
+ m1_23582_n3340# m1_12620_4059# m1_7706_n3340# m1_25472_4059# m1_5816_4059# m1_902_n3340#
+ m1_6950_n3340# m1_13376_4059# m1_22070_n3340# m1_9218_n3340# m1_2414_n3340# m1_9218_n3340#
+ m1_11486_n3340# m1_10352_4059# m1_17912_4059# m1_2414_n3340# m1_1280_4059# m1_24716_4059#
+ m1_10730_n3340# m1_6572_4059# m1_21692_4059# vtrip3 m1_9596_4059# m1_17912_4059#
+ m1_18290_n3340# m1_24716_4059# m1_25094_n3340# m1_2036_4059# vtrip6 m1_4682_n3340#
+ m1_20936_4059# m1_17156_4059# m1_8840_4059# m1_4682_n3340# m1_12620_4059# m1_3548_4059#
+ m1_25472_4059# sky130_fd_pr__res_xhigh_po_1p41_9VZRJ2
Xsky130_fd_pr__nfet_g5v0d10v5_CD9S2Z_0 avss avss vtop ena_b sky130_fd_pr__nfet_g5v0d10v5_CD9S2Z
C0 vtop ena_b 1.269212f
C1 otrip_decoded_avdd[1] avdd 0.274776f
C2 vout_vunder vtrip_decoded_avdd[6] 0.728099f
C3 vtrip2 vtrip4 0.698261f
C4 vtrip7 otrip_decoded_avdd[7] 0.325806f
C5 otrip_decoded_avdd[5] vout_brout 0.724289f
C6 otrip_decoded_avdd[6] avdd 0.271582f
C7 vtrip1 vout_vunder 0.500536f
C8 vtrip_decoded_avdd[1] vtrip_decoded_b_avdd[0] 0.142261f
C9 vtrip_decoded_avdd[1] vout_vunder 0.722951f
C10 vtrip3 vtrip5 0.11433f
C11 vtrip_decoded_avdd[3] vtrip_decoded_b_avdd[2] 0.142261f
C12 vtop avdd 2.545652f
C13 otrip_decoded_b_avdd[6] vout_brout 0.187792f
C14 vout_brout vtrip4 0.679853f
C15 vtrip_decoded_b_avdd[3] vout_vunder 0.187792f
C16 vtrip5 avdd 0.386901f
C17 vtrip_decoded_b_avdd[6] vtrip_decoded_avdd[6] 0.459706f
C18 otrip_decoded_avdd[5] otrip_decoded_b_avdd[4] 0.142261f
C19 vtrip_decoded_avdd[2] avdd 0.271582f
C20 vtrip0 vtrip5 0.1051f
C21 vtrip1 vtrip4 0.210041f
C22 otrip_decoded_b_avdd[2] otrip_decoded_avdd[2] 0.459706f
C23 vout_brout otrip_decoded_avdd[7] 0.722855f
C24 otrip_decoded_b_avdd[1] avdd 0.245102f
C25 vtrip_decoded_b_avdd[5] vtrip_decoded_avdd[5] 0.459706f
C26 vout_brout otrip_decoded_b_avdd[7] 0.187792f
C27 vout_brout otrip_decoded_b_avdd[2] 0.187792f
C28 vtrip_decoded_avdd[4] avdd 0.271582f
C29 vtrip_decoded_avdd[3] vtrip3 0.297998f
C30 vtrip6 vtrip3 1.14511f
C31 vtrip_decoded_b_avdd[2] avdd 0.244353f
C32 vtrip_decoded_avdd[7] avdd 0.278971f
C33 vtrip_decoded_avdd[5] avdd 0.271726f
C34 vtrip_decoded_avdd[3] avdd 0.271582f
C35 vtrip6 avdd 0.907111f
C36 otrip_decoded_avdd[6] otrip_decoded_b_avdd[6] 0.459706f
C37 otrip_decoded_b_avdd[0] avdd 0.249227f
C38 vtrip5 vout_vunder 0.91347f
C39 otrip_decoded_avdd[5] vtrip5 0.386893f
C40 vtrip_decoded_avdd[2] vout_vunder 0.722952f
C41 vtrip_decoded_avdd[1] vtrip_decoded_b_avdd[1] 0.459706f
C42 ena_b avdd 2.443612f
C43 vtrip_decoded_b_avdd[5] avdd 0.244436f
C44 vtrip2 otrip_decoded_avdd[2] 0.325432f
C45 vtrip7 vout_brout 0.493971f
C46 vtrip_decoded_avdd[4] vout_vunder 0.722914f
C47 vout_brout otrip_decoded_avdd[4] 0.726903f
C48 vtrip4 vtrip5 2.03217f
C49 vtrip3 otrip_decoded_avdd[3] 0.327608f
C50 vout_brout vtrip2 0.510824f
C51 vtrip3 avdd 1.044079f
C52 vout_vunder vtrip_decoded_b_avdd[2] 0.187792f
C53 vtrip1 vtrip2 2.346093f
C54 vtrip_decoded_avdd[7] vout_vunder 0.728002f
C55 otrip_decoded_avdd[3] avdd 0.271582f
C56 vout_vunder vtrip_decoded_avdd[5] 0.725363f
C57 vtrip_decoded_avdd[3] vout_vunder 0.722951f
C58 otrip_decoded_b_avdd[3] otrip_decoded_avdd[4] 0.142261f
C59 vtrip6 vout_vunder 0.505947f
C60 vtrip0 avdd 0.384663f
C61 vout_brout otrip_decoded_b_avdd[5] 0.187792f
C62 vout_brout otrip_decoded_avdd[2] 0.728099f
C63 vtrip_decoded_avdd[4] vtrip4 0.343878f
C64 vtrip7 m1_17156_4059# 0.120895f
C65 otrip_decoded_avdd[4] otrip_decoded_b_avdd[4] 0.459706f
C66 vtrip_decoded_avdd[7] vtrip_decoded_b_avdd[7] 0.459706f
C67 vtrip_decoded_avdd[0] avdd 0.271582f
C68 vtrip_decoded_avdd[0] vtrip0 0.332173f
C69 vout_vunder vtrip_decoded_b_avdd[5] 0.187792f
C70 vout_brout vtrip1 0.509964f
C71 vtrip_decoded_avdd[2] vtrip_decoded_b_avdd[1] 0.142261f
C72 vtrip6 vtrip4 0.563736f
C73 vout_brout otrip_decoded_avdd[0] 0.398767f
C74 vtrip_decoded_b_avdd[6] vtrip_decoded_avdd[7] 0.142261f
C75 vtrip_decoded_b_avdd[0] avdd 0.244353f
C76 vtrip3 vout_vunder 0.449946f
C77 otrip_decoded_b_avdd[3] vout_brout 0.187793f
C78 vout_vunder avdd 1.776475f
C79 m1_12620_4059# vtrip0 0.139758f
C80 vtrip_decoded_avdd[1] vtrip1 0.328174f
C81 otrip_decoded_avdd[5] avdd 0.271582f
C82 vtrip0 vout_vunder 0.445016f
C83 vout_brout otrip_decoded_b_avdd[4] 0.187792f
C84 vtrip_decoded_avdd[0] vtrip_decoded_b_avdd[0] 0.459706f
C85 otrip_decoded_avdd[6] otrip_decoded_b_avdd[5] 0.142261f
C86 vtrip_decoded_b_avdd[7] avdd 0.254243f
C87 vout_brout otrip_decoded_avdd[1] 0.728098f
C88 vtrip7 m1_19424_4059# 0.117324f
C89 vtrip_decoded_avdd[0] vout_vunder 0.398307f
C90 vtrip3 vtrip4 0.485368f
C91 vtrip1 otrip_decoded_avdd[1] 0.324162f
C92 otrip_decoded_b_avdd[6] avdd 0.244353f
C93 vtrip_decoded_avdd[2] vtrip2 0.326798f
C94 otrip_decoded_avdd[6] vout_brout 0.722951f
C95 vtrip4 avdd 0.369463f
C96 vtrip0 vtrip4 0.655887f
C97 vout_vunder vtrip_decoded_b_avdd[0] 0.115806f
C98 vtrip_decoded_b_avdd[6] avdd 0.244986f
C99 vtrip7 m1_17912_4059# 0.117887f
C100 otrip_decoded_avdd[7] avdd 0.271582f
C101 vtrip7 vtrip_decoded_avdd[7] 0.331307f
C102 vtrip_decoded_avdd[4] vtrip_decoded_b_avdd[4] 0.459706f
C103 otrip_decoded_b_avdd[2] otrip_decoded_avdd[3] 0.142261f
C104 otrip_decoded_b_avdd[1] otrip_decoded_avdd[2] 0.142261f
C105 vout_brout vtrip5 0.723097f
C106 avdd otrip_decoded_b_avdd[7] 0.244353f
C107 otrip_decoded_b_avdd[2] avdd 0.244453f
C108 vtrip6 vtrip7 2.124565f
C109 vtrip1 vtrip5 0.105864f
C110 vout_vunder vtrip_decoded_b_avdd[7] 0.187792f
C111 vout_brout otrip_decoded_b_avdd[1] 0.187792f
C112 vtrip_decoded_avdd[5] vtrip_decoded_b_avdd[4] 0.142261f
C113 vtrip_decoded_b_avdd[1] avdd 0.244353f
C114 vtrip_decoded_avdd[0] otrip_decoded_b_avdd[7] 0.142261f
C115 m1_13376_4059# vtrip0 0.412491f
C116 vtrip4 vout_vunder 0.642078f
C117 vtrip_decoded_b_avdd[6] vout_vunder 0.187792f
C118 vtrip6 vtrip_decoded_avdd[6] 0.334965f
C119 vtrip7 m1_20180_4059# 0.117324f
C120 vtrip6 vout_brout 0.499729f
C121 vtrip7 avdd 0.537919f
C122 otrip_decoded_b_avdd[0] vout_brout 0.115916f
C123 otrip_decoded_avdd[4] avdd 0.271582f
C124 vtrip_decoded_b_avdd[3] vtrip_decoded_avdd[4] 0.142261f
C125 vtrip2 vtrip3 2.049601f
C126 otrip_decoded_b_avdd[0] otrip_decoded_avdd[0] 0.459787f
C127 otrip_decoded_b_avdd[1] otrip_decoded_avdd[1] 0.459706f
C128 vtrip2 avdd 0.812936f
C129 otrip_decoded_b_avdd[6] otrip_decoded_avdd[7] 0.142261f
C130 vtrip7 m1_18668_4059# 0.117324f
C131 vtrip_decoded_b_avdd[5] vtrip_decoded_avdd[6] 0.142261f
C132 vtrip0 vtrip2 0.552137f
C133 vtrip_decoded_b_avdd[4] avdd 0.244353f
C134 vout_vunder vtrip_decoded_b_avdd[1] 0.187792f
C135 otrip_decoded_b_avdd[5] avdd 0.244353f
C136 vtrip_decoded_b_avdd[3] vtrip_decoded_avdd[3] 0.459706f
C137 otrip_decoded_avdd[2] avdd 0.271961f
C138 vout_brout vtrip3 0.512881f
C139 vtrip_decoded_avdd[6] avdd 0.272528f
C140 vout_brout otrip_decoded_avdd[3] 0.728099f
C141 vout_brout avdd 1.733791f
C142 otrip_decoded_avdd[7] otrip_decoded_b_avdd[7] 0.459706f
C143 otrip_decoded_b_avdd[0] otrip_decoded_avdd[1] 0.142261f
C144 vout_brout vtrip0 0.621824f
C145 vtrip7 vout_vunder 0.498953f
C146 vtrip1 avdd 0.511967f
C147 otrip_decoded_avdd[6] vtrip6 0.3362f
C148 vtrip0 vtrip1 2.290143f
C149 otrip_decoded_avdd[0] avdd 0.378054f
C150 vtrip0 otrip_decoded_avdd[0] 0.355328f
C151 vtrip2 vout_vunder 0.498413f
C152 otrip_decoded_b_avdd[3] otrip_decoded_avdd[3] 0.459706f
C153 vtrip_decoded_avdd[0] vout_brout 0.252789f
C154 otrip_decoded_b_avdd[3] avdd 0.244353f
C155 vtrip_decoded_avdd[1] avdd 0.271582f
C156 vout_vunder vtrip_decoded_b_avdd[4] 0.187792f
C157 vtrip_decoded_b_avdd[3] avdd 0.244353f
C158 vtrip5 vtrip_decoded_avdd[5] 0.381025f
C159 otrip_decoded_b_avdd[4] avdd 0.244353f
C160 vtrip_decoded_avdd[2] vtrip_decoded_b_avdd[2] 0.459706f
C161 vtrip6 vtrip5 0.346416f
C162 otrip_decoded_avdd[5] otrip_decoded_b_avdd[5] 0.459706f
C163 vtrip4 otrip_decoded_avdd[4] 0.379796f
C164 m1_26606_n3340# avss 1.233559f
C165 m1_26228_4059# avss 1.030713f
C166 m1_25850_n3340# avss 0.969126f
C167 m1_25472_4059# avss 1.028466f
C168 m1_25094_n3340# avss 0.969045f
C169 m1_24716_4059# avss 1.028161f
C170 m1_24338_n3340# avss 0.969044f
C171 m1_23960_4059# avss 1.028161f
C172 m1_23582_n3340# avss 0.969045f
C173 m1_23204_4059# avss 1.028161f
C174 m1_22826_n3340# avss 0.969044f
C175 m1_22448_4059# avss 1.028161f
C176 m1_22070_n3340# avss 0.969045f
C177 m1_21692_4059# avss 1.028161f
C178 m1_21314_n3340# avss 0.969044f
C179 m1_20936_4059# avss 0.987074f
C180 m1_20558_n3340# avss 0.969045f
C181 m1_20180_4059# avss 0.968689f
C182 m1_19802_n3340# avss 0.969045f
C183 m1_19424_4059# avss 0.968302f
C184 m1_19046_n3340# avss 0.969045f
C185 m1_18668_4059# avss 0.968346f
C186 m1_18290_n3340# avss 0.969044f
C187 m1_17912_4059# avss 0.968235f
C188 m1_17534_n3340# avss 0.969044f
C189 m1_17156_4059# avss 0.968264f
C190 m1_16778_n3340# avss 0.969045f
C191 vtrip7 avss 3.325846f
C192 vtrip6 avss 3.589394f
C193 vtrip5 avss 2.461755f
C194 vtrip4 avss 3.147402f
C195 vtrip3 avss 2.563879f
C196 vtrip2 avss 3.412884f
C197 vtrip1 avss 2.744727f
C198 vtrip0 avss 3.894833f
C199 m1_13376_4059# avss 0.968235f
C200 m1_12998_n3340# avss 0.969044f
C201 m1_12620_4059# avss 0.984676f
C202 m1_12242_n3340# avss 0.969045f
C203 m1_11864_4059# avss 0.967778f
C204 m1_11486_n3340# avss 0.969044f
C205 m1_11108_4059# avss 0.967778f
C206 m1_10730_n3340# avss 0.969045f
C207 m1_10352_4059# avss 0.967778f
C208 m1_9974_n3340# avss 0.969045f
C209 m1_9596_4059# avss 0.967778f
C210 m1_9218_n3340# avss 0.969045f
C211 m1_8840_4059# avss 0.967778f
C212 m1_8462_n3340# avss 0.969045f
C213 m1_8084_4059# avss 0.967778f
C214 m1_7706_n3340# avss 0.969044f
C215 m1_7328_4059# avss 0.967778f
C216 m1_6950_n3340# avss 0.969045f
C217 m1_6572_4059# avss 0.967778f
C218 m1_6194_n3340# avss 0.969045f
C219 m1_5816_4059# avss 0.967778f
C220 m1_5438_n3340# avss 0.969045f
C221 m1_5060_4059# avss 0.967778f
C222 m1_4682_n3340# avss 0.969044f
C223 m1_4304_4059# avss 0.967778f
C224 m1_3926_n3340# avss 0.969045f
C225 m1_3548_4059# avss 0.967778f
C226 m1_3170_n3340# avss 0.969044f
C227 m1_2792_4059# avss 0.967778f
C228 m1_2414_n3340# avss 0.969045f
C229 m1_2036_4059# avss 0.967806f
C230 m1_1658_n3340# avss 0.969127f
C231 m1_1280_4059# avss 0.967978f
C232 m1_902_n3340# avss 1.234363f
C233 vtop avss 5.492615f
C234 ena avss 0.399955f
C235 ena_b avss 3.064275f
C236 avdd avss 0.100503p
C237 vtrip_decoded_b_avdd[7] avss 0.625077f
C238 vtrip_decoded_b_avdd[6] avss 0.512921f
C239 vtrip_decoded_b_avdd[5] avss 0.512472f
C240 vtrip_decoded_b_avdd[4] avss 0.512168f
C241 vtrip_decoded_b_avdd[3] avss 0.512168f
C242 vtrip_decoded_b_avdd[2] avss 0.512168f
C243 vtrip_decoded_b_avdd[1] avss 0.512176f
C244 vtrip_decoded_b_avdd[0] avss 0.512168f
C245 otrip_decoded_b_avdd[7] avss 0.512168f
C246 otrip_decoded_b_avdd[6] avss 0.512168f
C247 otrip_decoded_b_avdd[5] avss 0.512168f
C248 otrip_decoded_b_avdd[4] avss 0.512168f
C249 otrip_decoded_b_avdd[3] avss 0.512168f
C250 otrip_decoded_b_avdd[2] avss 0.512725f
C251 otrip_decoded_b_avdd[1] avss 0.515018f
C252 otrip_decoded_b_avdd[0] avss 0.547834f
C253 vout_vunder avss 5.81703f
C254 vout_brout avss 5.622336f
C255 vtrip_decoded_avdd[7] avss 1.32506f
C256 vtrip_decoded_avdd[6] avss 1.21963f
C257 vtrip_decoded_avdd[5] avss 1.219459f
C258 vtrip_decoded_avdd[4] avss 1.218783f
C259 vtrip_decoded_avdd[3] avss 1.21877f
C260 vtrip_decoded_avdd[2] avss 1.218783f
C261 vtrip_decoded_avdd[1] avss 1.222296f
C262 vtrip_decoded_avdd[0] avss 1.218775f
C263 otrip_decoded_avdd[7] avss 1.218775f
C264 otrip_decoded_avdd[6] avss 1.21914f
C265 otrip_decoded_avdd[5] avss 1.218782f
C266 otrip_decoded_avdd[4] avss 1.218766f
C267 otrip_decoded_avdd[3] avss 1.218763f
C268 otrip_decoded_avdd[2] avss 1.219219f
C269 otrip_decoded_avdd[1] avss 1.220117f
C270 otrip_decoded_avdd[0] avss 1.484734f
.ends

.subckt sky130_fd_sc_hvl__inv_4 A VGND VNB VPB VPWR Y
X0 VPWR A Y VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.21 ps=1.78 w=1.5 l=0.5
X1 Y A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X2 VGND A Y VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X3 Y A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.4275 ps=3.57 w=1.5 l=0.5
X4 VGND A Y VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.105 ps=1.03 w=0.75 l=0.5
X5 Y A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X6 Y A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.21375 ps=2.07 w=0.75 l=0.5
X7 VPWR A Y VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
C0 Y A 0.703999f
C1 VGND A 0.225758f
C2 Y VPWR 0.628131f
C3 A VPWR 0.342778f
C4 A VPB 0.348469f
C5 VPWR VPB 0.665325f
C6 Y VGND 0.376222f
C7 VGND VNB 0.728214f
C8 Y VNB 0.118981f
C9 VPWR VNB 0.118266f
C10 A VNB 1.08046f
C11 VPB VNB 1.7136f
.ends

.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
C0 Y A 0.359887f
C1 Y VPWR 0.361779f
C2 A VPB 0.141975f
C3 Y VGND 0.262586f
C4 VGND VNB 0.326816f
C5 VPWR VNB 0.296394f
C6 A VNB 0.451855f
C7 VPB VNB 0.516168f
.ends

.subckt sky130_fd_pr__nfet_01v8_SCV3UK a_50_n131# a_n50_n157# a_n526_n243# a_n108_n131#
+ a_n266_n131# a_n424_n131# a_208_n131# a_108_n157# a_n208_n157# a_366_n131# a_266_n157#
+ a_n366_n157#
X0 a_n108_n131# a_n208_n157# a_n266_n131# a_n526_n243# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X1 a_208_n131# a_108_n157# a_50_n131# a_n526_n243# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X2 a_n266_n131# a_n366_n157# a_n424_n131# a_n526_n243# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X3 a_366_n131# a_266_n157# a_208_n131# a_n526_n243# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X4 a_50_n131# a_n50_n157# a_n108_n131# a_n526_n243# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
C0 a_366_n131# a_n526_n243# 0.144549f
C1 a_n424_n131# a_n526_n243# 0.144549f
C2 a_266_n157# a_n526_n243# 0.283278f
C3 a_108_n157# a_n526_n243# 0.245808f
C4 a_n50_n157# a_n526_n243# 0.245716f
C5 a_n208_n157# a_n526_n243# 0.245808f
C6 a_n366_n157# a_n526_n243# 0.283278f
.ends

.subckt sky130_fd_pr__pfet_01v8_BZXTE7 a_208_n64# a_n108_n64# a_998_n64# a_n898_n64#
+ a_108_n161# a_50_n64# a_n208_n161# a_266_n161# a_n424_n64# a_524_n64# a_898_n161#
+ a_n366_n161# a_424_n161# a_n998_n161# a_n266_n64# a_366_n64# a_n524_n161# a_582_n161#
+ a_n50_n161# a_840_n64# a_n740_n64# a_n682_n161# 0 a_740_n161# a_682_n64# a_n582_n64#
+ a_n840_n161# w_n1194_n284# a_n1056_n64#
X0 a_n898_n64# a_n998_n161# a_n1056_n64# w_n1194_n284# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X1 a_n582_n64# a_n682_n161# a_n740_n64# w_n1194_n284# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X2 a_50_n64# a_n50_n161# a_n108_n64# w_n1194_n284# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X3 a_n740_n64# a_n840_n161# a_n898_n64# w_n1194_n284# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X4 a_n266_n64# a_n366_n161# a_n424_n64# w_n1194_n284# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X5 a_n424_n64# a_n524_n161# a_n582_n64# w_n1194_n284# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X6 a_n108_n64# a_n208_n161# a_n266_n64# w_n1194_n284# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X7 a_998_n64# a_898_n161# a_840_n64# w_n1194_n284# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X8 a_682_n64# a_582_n161# a_524_n64# w_n1194_n284# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X9 a_840_n64# a_740_n161# a_682_n64# w_n1194_n284# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X10 a_366_n64# a_266_n161# a_208_n64# w_n1194_n284# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X11 a_524_n64# a_424_n161# a_366_n64# w_n1194_n284# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X12 a_208_n64# a_108_n161# a_50_n64# w_n1194_n284# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
C0 w_n1194_n284# a_n998_n161# 0.162265f
C1 a_424_n161# w_n1194_n284# 0.139032f
C2 w_n1194_n284# a_108_n161# 0.139f
C3 w_n1194_n284# a_266_n161# 0.139012f
C4 w_n1194_n284# a_n50_n161# 0.138996f
C5 a_n366_n161# w_n1194_n284# 0.139012f
C6 w_n1194_n284# a_n524_n161# 0.139032f
C7 a_898_n161# w_n1194_n284# 0.162265f
C8 w_n1194_n284# a_740_n161# 0.139244f
C9 a_n682_n161# w_n1194_n284# 0.139085f
C10 w_n1194_n284# a_582_n161# 0.139085f
C11 w_n1194_n284# a_n840_n161# 0.139244f
C12 w_n1194_n284# a_n208_n161# 0.139f
C13 a_898_n161# 0 0.126262f
C14 a_740_n161# 0 0.110061f
C15 a_582_n161# 0 0.110061f
C16 a_424_n161# 0 0.110061f
C17 a_266_n161# 0 0.110061f
C18 a_108_n161# 0 0.110061f
C19 a_n50_n161# 0 0.110061f
C20 a_n208_n161# 0 0.110061f
C21 a_n366_n161# 0 0.110061f
C22 a_n524_n161# 0 0.110061f
C23 a_n682_n161# 0 0.110061f
C24 a_n840_n161# 0 0.110061f
C25 a_n998_n161# 0 0.126262f
C26 w_n1194_n284# 0 5.57362f
.ends

.subckt schmitt_trigger in out dvdd dvss m
Xsky130_fd_pr__nfet_01v8_SCV3UK_1 m out dvss dvss m dvss dvss dvss in out m in sky130_fd_pr__nfet_01v8_SCV3UK
Xsky130_fd_pr__pfet_01v8_BZXTE7_0 dvdd dvdd out m out m in out dvdd dvdd m in dvdd
+ in m m in m out dvdd dvdd in dvss m out m in dvdd dvdd sky130_fd_pr__pfet_01v8_BZXTE7
C0 out dvdd 0.796706f
C1 out m 1.859932f
C2 in out 0.107481f
C3 dvdd m 1.037752f
C4 in dvdd 0.663292f
C5 in m 0.720533f
C6 out dvss 1.64006f
C7 m dvss 2.034164f
C8 in dvss 1.214657f
C9 dvdd dvss 6.619973f
.ends

.subckt sky130_fd_sc_hvl__lsbuflv2hv_1 A LVPWR VGND VNB VPB VPWR X
X0 VGND a_404_1133# a_504_1221# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X1 a_504_1221# a_404_1133# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X2 X a_1711_885# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.24375 ps=1.825 w=1.5 l=0.5
X3 X a_1711_885# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.121875 ps=1.075 w=0.75 l=0.5
X4 VGND A a_404_1133# VNB sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X5 a_1197_107# a_772_151# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X6 VPWR a_1197_107# a_504_1221# VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.2142 pd=1.99 as=0.2142 ps=1.99 w=0.42 l=1
X7 a_504_1221# a_404_1133# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X8 a_1197_107# a_772_151# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X9 a_772_151# a_404_1133# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X10 a_504_1221# a_404_1133# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X11 VGND a_404_1133# a_504_1221# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X12 LVPWR A a_404_1133# LVPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X13 VGND a_772_151# a_1197_107# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X14 VPWR a_504_1221# a_1711_885# VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.24375 pd=1.825 as=0.3975 ps=3.53 w=1.5 l=0.5
X15 VGND a_504_1221# a_1711_885# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.121875 pd=1.075 as=0.19875 ps=2.03 w=0.75 l=0.5
X16 VGND a_772_151# a_1197_107# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X17 a_772_151# a_404_1133# LVPWR LVPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X18 a_1197_107# a_772_151# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X19 VPWR a_504_1221# a_1197_107# VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.1365 ps=1.49 w=0.42 l=1
C0 VPWR a_1197_107# 0.247134f
C1 VPWR a_1711_885# 0.262393f
C2 a_504_1221# VGND 0.702325f
C3 LVPWR a_1197_107# 0.103614f
C4 a_504_1221# VPB 0.570551f
C5 a_772_151# VGND 0.646883f
C6 LVPWR VPWR 1.310519f
C7 a_772_151# VPB 0.116911f
C8 VPWR a_404_1133# 0.120704f
C9 a_1197_107# a_504_1221# 0.264594f
C10 a_504_1221# a_1711_885# 0.28899f
C11 VPWR a_504_1221# 0.272656f
C12 a_1197_107# a_772_151# 0.460766f
C13 a_1197_107# VGND 0.634871f
C14 LVPWR a_404_1133# 0.378765f
C15 a_1711_885# VGND 0.164303f
C16 a_1197_107# VPB 0.336238f
C17 VPWR VGND 0.168962f
C18 X a_1711_885# 0.108338f
C19 a_1711_885# VPB 0.154759f
C20 A a_404_1133# 0.182372f
C21 VPWR X 0.120607f
C22 VPWR VPB 2.72025f
C23 a_404_1133# a_504_1221# 0.40546f
C24 LVPWR a_772_151# 0.168977f
C25 LVPWR VGND 0.193471f
C26 LVPWR VPB 0.11581f
C27 a_404_1133# a_772_151# 0.138963f
C28 a_404_1133# VGND 0.578546f
C29 VGND VNB 3.86422f
C30 A VNB 0.261789f
C31 VPWR VNB 0.273779f
C32 X VNB 0.143785f
C33 LVPWR VNB 0.577555f
C34 VPB VNB 2.88904f
C35 a_772_151# VNB 1.04864f
C36 a_1197_107# VNB 0.25514f
C37 a_1711_885# VNB 0.339894f
C38 a_504_1221# VNB 0.834376f
C39 a_404_1133# VNB 1.44294f
.ends

.subckt sky130_fd_pr__pfet_01v8_MA8JJJ a_18_n136# a_n33_95# w_n112_n198# a_n76_n136#
X0 a_18_n136# a_n33_95# a_n76_n136# w_n112_n198# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.18
C0 a_18_n136# a_n76_n136# 0.151817f
C1 a_18_n136# 0 0.109283f
C2 a_n76_n136# 0 0.109283f
C3 a_n33_95# 0 0.15012f
C4 w_n112_n198# 0 0.243264f
.ends

.subckt sky130_fd_pr__res_xhigh_po_1p41_ZB8LT7 a_1560_11084# a_48_n11516# a_n1972_n11646#
+ a_804_n11516# a_1560_n11516# a_48_11084# a_n330_11084# a_n708_11084# a_426_n11516#
+ a_n1086_11084# a_n1464_11084# a_1182_n11516# a_n1842_11084# a_n330_n11516# a_n1842_n11516#
+ a_n708_n11516# a_426_11084# a_804_11084# a_n1464_n11516# a_1182_11084# a_n1086_n11516#
X0 a_804_11084# a_804_n11516# a_n1972_n11646# sky130_fd_pr__res_xhigh_po_1p41 l=111
X1 a_n1464_11084# a_n1464_n11516# a_n1972_n11646# sky130_fd_pr__res_xhigh_po_1p41 l=111
X2 a_426_11084# a_426_n11516# a_n1972_n11646# sky130_fd_pr__res_xhigh_po_1p41 l=111
X3 a_n708_11084# a_n708_n11516# a_n1972_n11646# sky130_fd_pr__res_xhigh_po_1p41 l=111
X4 a_1560_11084# a_1560_n11516# a_n1972_n11646# sky130_fd_pr__res_xhigh_po_1p41 l=111
X5 a_n1086_11084# a_n1086_n11516# a_n1972_n11646# sky130_fd_pr__res_xhigh_po_1p41 l=111
X6 a_n1842_11084# a_n1842_n11516# a_n1972_n11646# sky130_fd_pr__res_xhigh_po_1p41 l=111
X7 a_n330_11084# a_n330_n11516# a_n1972_n11646# sky130_fd_pr__res_xhigh_po_1p41 l=111
X8 a_1182_11084# a_1182_n11516# a_n1972_n11646# sky130_fd_pr__res_xhigh_po_1p41 l=111
X9 a_48_11084# a_48_n11516# a_n1972_n11646# sky130_fd_pr__res_xhigh_po_1p41 l=111
C0 a_n330_n11516# a_n708_n11516# 0.296258f
C1 a_426_n11516# a_48_n11516# 0.296258f
C2 a_1560_n11516# a_1182_n11516# 0.296258f
C3 a_1182_11084# a_804_11084# 0.296258f
C4 a_n1464_n11516# a_n1842_n11516# 0.296258f
C5 a_n708_n11516# a_n1086_n11516# 0.296258f
C6 a_48_11084# a_426_11084# 0.296258f
C7 a_n330_n11516# a_48_n11516# 0.296258f
C8 a_n330_11084# a_n708_11084# 0.296258f
C9 a_n1842_11084# a_n1464_11084# 0.296258f
C10 a_426_11084# a_804_11084# 0.296258f
C11 a_804_n11516# a_426_n11516# 0.296258f
C12 a_n1086_11084# a_n708_11084# 0.296258f
C13 a_n1464_11084# a_n1086_11084# 0.296258f
C14 a_1560_11084# a_1182_11084# 0.296258f
C15 a_n1086_n11516# a_n1464_n11516# 0.296258f
C16 a_804_n11516# a_1182_n11516# 0.296258f
C17 a_48_11084# a_n330_11084# 0.296258f
C18 a_1560_n11516# a_n1972_n11646# 0.62945f
C19 a_1560_11084# a_n1972_n11646# 0.62945f
C20 a_1182_n11516# a_n1972_n11646# 0.419137f
C21 a_1182_11084# a_n1972_n11646# 0.419137f
C22 a_804_n11516# a_n1972_n11646# 0.419137f
C23 a_804_11084# a_n1972_n11646# 0.419137f
C24 a_426_n11516# a_n1972_n11646# 0.419137f
C25 a_426_11084# a_n1972_n11646# 0.419137f
C26 a_48_n11516# a_n1972_n11646# 0.419137f
C27 a_48_11084# a_n1972_n11646# 0.419137f
C28 a_n330_n11516# a_n1972_n11646# 0.419137f
C29 a_n330_11084# a_n1972_n11646# 0.419137f
C30 a_n708_n11516# a_n1972_n11646# 0.419137f
C31 a_n708_11084# a_n1972_n11646# 0.419137f
C32 a_n1086_n11516# a_n1972_n11646# 0.419137f
C33 a_n1086_11084# a_n1972_n11646# 0.419137f
C34 a_n1464_n11516# a_n1972_n11646# 0.419137f
C35 a_n1464_11084# a_n1972_n11646# 0.419137f
C36 a_n1842_n11516# a_n1972_n11646# 0.62945f
C37 a_n1842_11084# a_n1972_n11646# 0.62945f
.ends

.subckt sky130_fd_pr__pfet_01v8_LAUYMQ w_n161_n200# a_n125_n100# a_66_n100# a_15_131#
+ a_n30_n100# a_n81_n197#
X0 a_n30_n100# a_n81_n197# a_n125_n100# w_n161_n200# sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.295 ps=2.59 w=1 l=0.18
X1 a_66_n100# a_15_131# a_n30_n100# w_n161_n200# sky130_fd_pr__pfet_01v8 ad=0.295 pd=2.59 as=0.15 ps=1.3 w=1 l=0.18
C0 a_n30_n100# a_n125_n100# 0.148887f
C1 a_n30_n100# a_66_n100# 0.148887f
C2 a_66_n100# 0 0.109727f
C3 a_n125_n100# 0 0.109727f
C4 a_n81_n197# 0 0.137231f
C5 a_15_131# 0 0.137231f
C6 w_n161_n200# 0 0.364512f
.ends

.subckt sky130_fd_pr__pfet_01v8_C64SS5 a_287_n64# a_n187_n64# a_129_n64# w_n539_n164#
+ a_29_n161# a_n129_n161# a_187_n161# a_n29_n64# a_n287_n161# a_n503_n64# a_345_n161#
+ a_n345_n64# a_445_n64# a_n445_n161#
X0 a_129_n64# a_29_n161# a_n29_n64# w_n539_n164# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X1 a_n187_n64# a_n287_n161# a_n345_n64# w_n539_n164# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X2 a_n345_n64# a_n445_n161# a_n503_n64# w_n539_n164# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X3 a_n29_n64# a_n129_n161# a_n187_n64# w_n539_n164# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X4 a_287_n64# a_187_n161# a_129_n64# w_n539_n164# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X5 a_445_n64# a_345_n161# a_287_n64# w_n539_n164# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
C0 a_445_n64# 0 0.114157f
C1 a_n503_n64# 0 0.114157f
C2 a_345_n161# 0 0.199722f
C3 a_187_n161# 0 0.169394f
C4 a_29_n161# 0 0.169394f
C5 a_n129_n161# 0 0.169394f
C6 a_n287_n161# 0 0.169394f
C7 a_n445_n161# 0 0.199722f
C8 w_n539_n164# 0 1.17071f
.ends

.subckt sky130_fd_pr__cap_mim_m3_2_LUWKLG c2_n3269_n19000# m4_n3349_n19080#
X0 c2_n3269_n19000# m4_n3349_n19080# sky130_fd_pr__cap_mim_m3_2 l=30 w=30
X1 c2_n3269_n19000# m4_n3349_n19080# sky130_fd_pr__cap_mim_m3_2 l=30 w=30
X2 c2_n3269_n19000# m4_n3349_n19080# sky130_fd_pr__cap_mim_m3_2 l=30 w=30
X3 c2_n3269_n19000# m4_n3349_n19080# sky130_fd_pr__cap_mim_m3_2 l=30 w=30
X4 c2_n3269_n19000# m4_n3349_n19080# sky130_fd_pr__cap_mim_m3_2 l=30 w=30
X5 c2_n3269_n19000# m4_n3349_n19080# sky130_fd_pr__cap_mim_m3_2 l=30 w=30
C0 m4_n3349_n19080# c2_n3269_n19000# 0.407926p
C1 c2_n3269_n19000# 0 10.8139f
C2 m4_n3349_n19080# 0 77.859604f
.ends

.subckt sky130_fd_pr__pfet_01v8_2XUZHN a_n73_n100# w_n109_n162# a_15_n100# a_n15_n126#
X0 a_15_n100# a_n15_n126# a_n73_n100# w_n109_n162# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
C0 a_15_n100# a_n73_n100# 0.162113f
C1 a_15_n100# 0 0.111398f
C2 a_n73_n100# 0 0.111398f
C3 w_n109_n162# 0 0.211896f
.ends

.subckt sky130_fd_pr__pfet_01v8_C68ZY6 a_208_n64# a_n108_n64# a_108_n161# w_n618_n164#
+ a_50_n64# a_n208_n161# a_266_n161# a_n424_n64# a_524_n64# a_n366_n161# a_424_n161#
+ a_n266_n64# a_366_n64# a_n524_n161# a_n50_n161# a_n582_n64#
X0 a_50_n64# a_n50_n161# a_n108_n64# w_n618_n164# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X1 a_n266_n64# a_n366_n161# a_n424_n64# w_n618_n164# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X2 a_n424_n64# a_n524_n161# a_n582_n64# w_n618_n164# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X3 a_n108_n64# a_n208_n161# a_n266_n64# w_n618_n164# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X4 a_366_n64# a_266_n161# a_208_n64# w_n618_n164# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X5 a_524_n64# a_424_n161# a_366_n64# w_n618_n164# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X6 a_208_n64# a_108_n161# a_50_n64# w_n618_n164# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
C0 a_524_n64# 0 0.114157f
C1 a_n582_n64# 0 0.114157f
C2 a_424_n161# 0 0.199722f
C3 a_266_n161# 0 0.169394f
C4 a_108_n161# 0 0.169394f
C5 a_n50_n161# 0 0.169394f
C6 a_n208_n161# 0 0.169394f
C7 a_n366_n161# 0 0.169394f
C8 a_n524_n161# 0 0.199722f
C9 w_n618_n164# 0 1.3423f
.ends

.subckt sky130_fd_pr__pfet_01v8_C6GQGA w_n154_n164# a_n118_n64# a_60_n64# a_n60_n161#
X0 a_60_n64# a_n60_n161# a_n118_n64# w_n154_n164# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.6
C0 a_60_n64# 0 0.115203f
C1 a_n118_n64# 0 0.115203f
C2 a_n60_n161# 0 0.265217f
C3 w_n154_n164# 0 0.334488f
.ends

.subckt sky130_fd_pr__pfet_01v8_9QCJ55 a_358_n64# a_n158_n64# a_158_n161# a_n358_n161#
+ a_n100_n161# w_n452_n164# a_100_n64# a_n416_n64#
X0 a_100_n64# a_n100_n161# a_n158_n64# w_n452_n164# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1 a_358_n64# a_158_n161# a_100_n64# w_n452_n164# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2 a_n158_n64# a_n358_n161# a_n416_n64# w_n452_n164# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
C0 w_n452_n164# a_158_n161# 0.114821f
C1 w_n452_n164# a_n358_n161# 0.114821f
C2 w_n452_n164# a_n100_n161# 0.10872f
C3 a_358_n64# 0 0.119027f
C4 a_n416_n64# 0 0.119027f
C5 a_158_n161# 0 0.375556f
C6 a_n100_n161# 0 0.345228f
C7 a_n358_n161# 0 0.375556f
C8 w_n452_n164# 0 0.981744f
.ends

.subckt sky130_fd_pr__pfet_01v8_MLERZ7 a_50_n136# a_n108_n136# a_n50_n162# w_n144_n198#
X0 a_50_n136# a_n50_n162# a_n108_n136# w_n144_n198# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
C0 a_50_n136# 0 0.114157f
C1 a_n108_n136# 0 0.114157f
C2 a_n50_n162# 0 0.23005f
C3 w_n144_n198# 0 0.312768f
.ends

.subckt rc_osc dvdd out ena vr dvss
Xsky130_fd_pr__pfet_01v8_MA8JJJ_0 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_MA8JJJ
Xsky130_fd_pr__res_xhigh_po_1p41_ZB8LT7_0 m1_25146_n1894# m1_2270_n760# dvss m1_2270_n1516#
+ in m1_25146_n382# m1_25146_n382# m1_25146_374# m1_2270_n760# m1_25146_374# m1_25146_1130#
+ m1_2270_n1516# m1_25146_1130# m1_2270_n4# vr m1_2270_n4# m1_25146_n1138# m1_25146_n1138#
+ m1_2270_752# m1_25146_n1894# m1_2270_752# sky130_fd_pr__res_xhigh_po_1p41_ZB8LT7
Xsky130_fd_pr__pfet_01v8_LAUYMQ_0 dvdd dvdd vr ena_b out dvdd sky130_fd_pr__pfet_01v8_LAUYMQ
Xsky130_fd_pr__pfet_01v8_C64SS5_0 m dvdd dvdd dvdd in in in m in dvdd in m dvdd in
+ sky130_fd_pr__pfet_01v8_C64SS5
Xsky130_fd_pr__cap_mim_m3_2_LUWKLG_0 in dvss sky130_fd_pr__cap_mim_m3_2_LUWKLG
Xsky130_fd_pr__pfet_01v8_2XUZHN_0 in dvdd dvdd ena sky130_fd_pr__pfet_01v8_2XUZHN
Xsky130_fd_pr__pfet_01v8_C68ZY6_0 out n n dvdd dvdd m n n out m n dvdd dvdd dvdd m
+ m sky130_fd_pr__pfet_01v8_C68ZY6
Xsky130_fd_pr__pfet_01v8_C6GQGA_0 dvdd dvdd ena_b ena sky130_fd_pr__pfet_01v8_C6GQGA
Xsky130_fd_pr__pfet_01v8_9QCJ55_0 m m n n n dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_9QCJ55
Xsky130_fd_pr__pfet_01v8_MLERZ7_0 vr ena_b dvdd dvdd sky130_fd_pr__pfet_01v8_MLERZ7
X0 dvss dvss m dvss sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X1 m n dvss dvss sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2 dvss ena ena_b dvss sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.6
X3 out ena vr dvss sky130_fd_pr__nfet_01v8 ad=0.15 pd=1.3 as=0.1475 ps=1.295 w=1 l=0.18
X4 dvss dvss n dvss sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X5 dvss in m dvss sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X6 n m dvss dvss sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X7 dvss dvss out dvss sky130_fd_pr__nfet_01v8 ad=0.1475 pd=1.295 as=0.15 ps=1.3 w=1 l=0.18
X8 m in dvss dvss sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.1475 ps=1.295 w=1 l=0.5
X9 vr dvss dvss dvss sky130_fd_pr__nfet_01v8 ad=0.1475 pd=1.295 as=0.145 ps=1.29 w=1 l=0.6
X10 out n dvss dvss sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
C0 dvss vr 3.277629f
C1 in n 0.388742f
C2 dvss m 2.895181f
C3 dvss m1_2270_752# 0.474378f
C4 dvss m1_2270_n4# 0.474206f
C5 ena dvdd 0.633745f
C6 in ena_b 0.13356f
C7 m1_2270_n1516# in 0.474451f
C8 dvdd out 0.790288f
C9 ena out 0.143309f
C10 in dvdd 4.603239f
C11 ena in 0.155847f
C12 vr n 0.101782f
C13 n m 1.771966f
C14 vr ena_b 0.643266f
C15 in out 1.056859f
C16 dvss n 2.848999f
C17 dvss ena_b 1.209955f
C18 in m1_2270_n760# 0.516433f
C19 vr dvdd 1.140019f
C20 dvdd m 1.307017f
C21 ena vr 0.245726f
C22 ena m 0.252627f
C23 m1_2270_n1516# dvss 0.439492f
C24 dvss m1_25146_n382# 0.302983f
C25 dvss m1_25146_374# 0.305194f
C26 dvss dvdd 0.357331p
C27 vr out 0.537831f
C28 ena dvss 1.84657f
C29 m out 1.092154f
C30 in vr 0.495731f
C31 in m 1.009668f
C32 dvss out 3.041751f
C33 dvss m1_25146_n1894# 0.447179f
C34 in dvss 22.095154f
C35 m1_25146_1130# dvss 0.44257f
C36 dvss m1_2270_n760# 0.441536f
C37 dvdd n 1.849724f
C38 vr m 0.559422f
C39 dvss m1_25146_n1138# 0.303066f
C40 dvdd ena_b 0.30526f
C41 ena ena_b 0.469291f
C42 n out 0.92079f
C43 n 0 0.962242f
C44 ena_b 0 0.185393f
C45 ena 0 0.348082f
C46 dvdd 0 0.205349p
C47 dvss 0 79.7988f
C48 m 0 0.458106f
C49 in 0 17.843658f
C50 vr 0 0.974916f
C51 out 0 0.241293f
C52 m1_25146_n1894# 0 0.830903f
C53 m1_2270_n1516# 0 0.690318f
C54 m1_25146_n1138# 0 0.687159f
C55 m1_2270_n760# 0 0.690318f
C56 m1_25146_n382# 0 0.687159f
C57 m1_2270_n4# 0 0.690318f
C58 m1_25146_374# 0 0.687159f
C59 m1_2270_752# 0 0.690318f
C60 m1_25146_1130# 0 0.830903f
.ends

.subckt sky130_fd_sc_hvl__inv_16 A VGND VNB VPB VPWR Y
X0 VPWR A Y VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X1 Y A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X2 Y A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X3 VGND A Y VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X4 VPWR A Y VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X5 Y A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X6 VGND A Y VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X7 VPWR A Y VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X8 Y A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X9 VGND A Y VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X10 Y A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X11 VPWR A Y VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X12 VPWR A Y VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X13 VGND A Y VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X14 VGND A Y VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X15 VPWR A Y VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X16 Y A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X17 VGND A Y VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X18 Y A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X19 VPWR A Y VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X20 Y A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X21 Y A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X22 VGND A Y VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.2025 pd=2.04 as=0.105 ps=1.03 w=0.75 l=0.5
X23 Y A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X24 Y A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X25 Y A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X26 VPWR A Y VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X27 Y A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.19875 ps=2.03 w=0.75 l=0.5
X28 Y A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X29 VGND A Y VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X30 Y A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X31 Y A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
C0 Y VPB 0.243556f
C1 VPB A 1.28194f
C2 Y VPWR 3.23737f
C3 VPWR A 1.67031f
C4 Y A 2.32857f
C5 Y VGND 0.943812f
C6 VGND A 1.84449f
C7 VPB VPWR 2.19858f
C8 VGND VNB 2.40673f
C9 Y VNB 0.148266f
C10 VPWR VNB 0.105937f
C11 A VNB 3.49591f
C12 VPB VNB 5.44152f
.ends

.subckt sky130_fd_pr__res_xhigh_po_1p41_DVQADA a_48_n3916# a_n330_n3916# a_n708_n3916#
+ a_1182_3484# a_n2598_3484# a_n3354_n3916# a_n1086_n3916# a_n3732_n3916# a_n1464_n3916#
+ a_2694_n3916# a_n1842_n3916# a_n3862_n4046# a_1938_3484# a_48_3484# a_n1842_3484#
+ a_n2220_3484# a_2316_3484# a_426_n3916# a_1560_3484# a_n2976_3484# a_804_n3916#
+ a_n3354_3484# a_3072_n3916# a_426_3484# a_n2220_n3916# a_3450_n3916# a_n708_3484#
+ a_2694_3484# a_1182_n3916# a_1938_n3916# a_1560_n3916# a_3072_3484# a_n1086_3484#
+ a_n330_3484# a_n2598_n3916# a_n3732_3484# a_804_3484# a_n2976_n3916# a_2316_n3916#
+ a_3450_3484# a_n1464_3484#
X0 a_n330_3484# a_n330_n3916# a_n3862_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X1 a_3072_3484# a_3072_n3916# a_n3862_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X2 a_2316_3484# a_2316_n3916# a_n3862_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X3 a_n1086_3484# a_n1086_n3916# a_n3862_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X4 a_n3354_3484# a_n3354_n3916# a_n3862_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X5 a_n2220_3484# a_n2220_n3916# a_n3862_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X6 a_1938_3484# a_1938_n3916# a_n3862_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X7 a_2694_3484# a_2694_n3916# a_n3862_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X8 a_1560_3484# a_1560_n3916# a_n3862_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X9 a_n2976_3484# a_n2976_n3916# a_n3862_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X10 a_48_3484# a_48_n3916# a_n3862_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X11 a_n1842_3484# a_n1842_n3916# a_n3862_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X12 a_804_3484# a_804_n3916# a_n3862_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X13 a_n708_3484# a_n708_n3916# a_n3862_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X14 a_1182_3484# a_1182_n3916# a_n3862_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X15 a_n2598_3484# a_n2598_n3916# a_n3862_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X16 a_3450_3484# a_3450_n3916# a_n3862_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X17 a_n3732_3484# a_n3732_n3916# a_n3862_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X18 a_n1464_3484# a_n1464_n3916# a_n3862_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X19 a_426_3484# a_426_n3916# a_n3862_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
C0 a_2316_3484# a_1938_3484# 0.296258f
C1 a_2694_3484# a_2316_3484# 0.296258f
C2 a_n3354_3484# a_n3732_3484# 0.296258f
C3 a_426_n3916# a_48_n3916# 0.296258f
C4 a_n2220_3484# a_n2598_3484# 0.296258f
C5 a_n3354_3484# a_n2976_3484# 0.296258f
C6 a_48_3484# a_n330_3484# 0.296258f
C7 a_426_n3916# a_804_n3916# 0.296258f
C8 a_n1086_3484# a_n1464_3484# 0.296258f
C9 a_1560_n3916# a_1182_n3916# 0.296258f
C10 a_n1464_3484# a_n1842_3484# 0.296258f
C11 a_n2220_n3916# a_n1842_n3916# 0.296258f
C12 a_1560_n3916# a_1938_n3916# 0.296258f
C13 a_1938_n3916# a_2316_n3916# 0.296258f
C14 a_n2220_n3916# a_n2598_n3916# 0.296258f
C15 a_1182_3484# a_1560_3484# 0.296258f
C16 a_48_3484# a_426_3484# 0.296258f
C17 a_2694_n3916# a_3072_n3916# 0.296258f
C18 a_n3732_n3916# a_n3354_n3916# 0.296258f
C19 a_n1086_n3916# a_n708_n3916# 0.296258f
C20 a_n1086_n3916# a_n1464_n3916# 0.296258f
C21 a_3072_n3916# a_3450_n3916# 0.296258f
C22 a_n2220_3484# a_n1842_3484# 0.296258f
C23 a_n1464_n3916# a_n1842_n3916# 0.296258f
C24 a_n330_n3916# a_n708_n3916# 0.296258f
C25 a_n1086_3484# a_n708_3484# 0.296258f
C26 a_2694_n3916# a_2316_n3916# 0.296258f
C27 a_804_3484# a_426_3484# 0.296258f
C28 a_n708_3484# a_n330_3484# 0.296258f
C29 a_1560_3484# a_1938_3484# 0.296258f
C30 a_n2598_3484# a_n2976_3484# 0.296258f
C31 a_2694_3484# a_3072_3484# 0.296258f
C32 a_n2976_n3916# a_n3354_n3916# 0.296258f
C33 a_n2598_n3916# a_n2976_n3916# 0.296258f
C34 a_48_n3916# a_n330_n3916# 0.296258f
C35 a_3450_3484# a_3072_3484# 0.296258f
C36 a_1182_3484# a_804_3484# 0.296258f
C37 a_804_n3916# a_1182_n3916# 0.296258f
C38 a_3450_n3916# a_n3862_n4046# 0.62945f
C39 a_3450_3484# a_n3862_n4046# 0.62945f
C40 a_3072_n3916# a_n3862_n4046# 0.419137f
C41 a_3072_3484# a_n3862_n4046# 0.419137f
C42 a_2694_n3916# a_n3862_n4046# 0.419137f
C43 a_2694_3484# a_n3862_n4046# 0.419137f
C44 a_2316_n3916# a_n3862_n4046# 0.419137f
C45 a_2316_3484# a_n3862_n4046# 0.419137f
C46 a_1938_n3916# a_n3862_n4046# 0.419137f
C47 a_1938_3484# a_n3862_n4046# 0.419137f
C48 a_1560_n3916# a_n3862_n4046# 0.419137f
C49 a_1560_3484# a_n3862_n4046# 0.419137f
C50 a_1182_n3916# a_n3862_n4046# 0.419137f
C51 a_1182_3484# a_n3862_n4046# 0.419137f
C52 a_804_n3916# a_n3862_n4046# 0.419137f
C53 a_804_3484# a_n3862_n4046# 0.419137f
C54 a_426_n3916# a_n3862_n4046# 0.419137f
C55 a_426_3484# a_n3862_n4046# 0.419137f
C56 a_48_n3916# a_n3862_n4046# 0.419137f
C57 a_48_3484# a_n3862_n4046# 0.419137f
C58 a_n330_n3916# a_n3862_n4046# 0.419137f
C59 a_n330_3484# a_n3862_n4046# 0.419137f
C60 a_n708_n3916# a_n3862_n4046# 0.419137f
C61 a_n708_3484# a_n3862_n4046# 0.419137f
C62 a_n1086_n3916# a_n3862_n4046# 0.419137f
C63 a_n1086_3484# a_n3862_n4046# 0.419137f
C64 a_n1464_n3916# a_n3862_n4046# 0.419137f
C65 a_n1464_3484# a_n3862_n4046# 0.419137f
C66 a_n1842_n3916# a_n3862_n4046# 0.419137f
C67 a_n1842_3484# a_n3862_n4046# 0.419137f
C68 a_n2220_n3916# a_n3862_n4046# 0.419137f
C69 a_n2220_3484# a_n3862_n4046# 0.419137f
C70 a_n2598_n3916# a_n3862_n4046# 0.419137f
C71 a_n2598_3484# a_n3862_n4046# 0.419137f
C72 a_n2976_n3916# a_n3862_n4046# 0.419137f
C73 a_n2976_3484# a_n3862_n4046# 0.419137f
C74 a_n3354_n3916# a_n3862_n4046# 0.419137f
C75 a_n3354_3484# a_n3862_n4046# 0.419137f
C76 a_n3732_n3916# a_n3862_n4046# 0.62945f
C77 a_n3732_3484# a_n3862_n4046# 0.62945f
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_XZ4X25 a_n887_n588# a_n429_n588# a_487_n588#
+ a_n945_n500# a_29_n588# a_n487_n500# a_n1079_n722# a_n29_n500# a_887_n500# a_429_n500#
X0 a_n29_n500# a_n429_n588# a_n487_n500# a_n1079_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X1 a_429_n500# a_29_n588# a_n29_n500# a_n1079_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X2 a_887_n500# a_487_n588# a_429_n500# a_n1079_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=2
X3 a_n487_n500# a_n887_n588# a_n945_n500# a_n1079_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=2
C0 a_487_n588# a_429_n500# 0.161415f
C1 a_n887_n588# a_n487_n500# 0.161415f
C2 a_n29_n500# a_429_n500# 0.154106f
C3 a_n945_n500# a_n487_n500# 0.154106f
C4 a_n429_n588# a_n29_n500# 0.161415f
C5 a_29_n588# a_487_n588# 0.104496f
C6 a_n887_n588# a_n945_n500# 0.161415f
C7 a_n429_n588# a_n487_n500# 0.161415f
C8 a_29_n588# a_429_n500# 0.161415f
C9 a_n29_n500# a_n487_n500# 0.154106f
C10 a_n429_n588# a_n887_n588# 0.104496f
C11 a_887_n500# a_487_n588# 0.161415f
C12 a_n429_n588# a_29_n588# 0.104496f
C13 a_887_n500# a_429_n500# 0.154106f
C14 a_29_n588# a_n29_n500# 0.161415f
C15 a_887_n500# a_n1079_n722# 0.592008f
C16 a_429_n500# a_n1079_n722# 0.243437f
C17 a_n29_n500# a_n1079_n722# 0.243437f
C18 a_n487_n500# a_n1079_n722# 0.243437f
C19 a_n945_n500# a_n1079_n722# 0.592008f
C20 a_487_n588# a_n1079_n722# 1.21272f
C21 a_29_n588# a_n1079_n722# 1.14992f
C22 a_n429_n588# a_n1079_n722# 1.14992f
C23 a_n887_n588# a_n1079_n722# 1.21272f
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_Y9S9FP a_n1174_n500# a_n200_n597# a_200_n500#
+ a_n1116_n597# a_n716_n500# 0 a_n258_n500# w_n1374_n797# a_1116_n500# a_n658_n597#
+ a_658_n500# a_716_n597# a_258_n597#
X0 a_1116_n500# a_716_n597# a_658_n500# w_n1374_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=2
X1 a_200_n500# a_n200_n597# a_n258_n500# w_n1374_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X2 a_n716_n500# a_n1116_n597# a_n1174_n500# w_n1374_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=2
X3 a_658_n500# a_258_n597# a_200_n500# w_n1374_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X4 a_n258_n500# a_n658_n597# a_n716_n500# w_n1374_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
C0 a_658_n500# a_716_n597# 0.161415f
C1 a_n658_n597# a_n1116_n597# 0.109462f
C2 a_n1116_n597# a_n716_n500# 0.161415f
C3 w_n1374_n797# a_716_n597# 0.682905f
C4 a_n658_n597# a_n716_n500# 0.161415f
C5 a_200_n500# a_n200_n597# 0.161415f
C6 a_716_n597# a_1116_n500# 0.161415f
C7 a_n200_n597# w_n1374_n797# 0.640116f
C8 a_n1174_n500# a_n1116_n597# 0.161415f
C9 a_716_n597# a_258_n597# 0.109462f
C10 a_n258_n500# a_n200_n597# 0.161415f
C11 a_n200_n597# a_258_n597# 0.109462f
C12 a_n1116_n597# w_n1374_n797# 0.682905f
C13 a_n1174_n500# a_n716_n500# 0.154106f
C14 a_n658_n597# w_n1374_n797# 0.640116f
C15 a_n658_n597# a_n258_n500# 0.161415f
C16 a_200_n500# a_658_n500# 0.154106f
C17 a_n258_n500# a_n716_n500# 0.154106f
C18 a_658_n500# a_1116_n500# 0.154106f
C19 a_n1174_n500# w_n1374_n797# 0.305433f
C20 a_658_n500# a_258_n597# 0.161415f
C21 a_200_n500# a_n258_n500# 0.154106f
C22 a_200_n500# a_258_n597# 0.161415f
C23 w_n1374_n797# a_1116_n500# 0.305433f
C24 w_n1374_n797# a_258_n597# 0.640116f
C25 a_n658_n597# a_n200_n597# 0.109462f
C26 a_1116_n500# 0 0.288363f
C27 a_658_n500# 0 0.221345f
C28 a_200_n500# 0 0.221345f
C29 a_n258_n500# 0 0.221345f
C30 a_n716_n500# 0 0.221345f
C31 a_n1174_n500# 0 0.288363f
C32 a_716_n597# 0 0.557987f
C33 a_258_n597# 0 0.53443f
C34 a_n200_n597# 0 0.53443f
C35 a_n658_n597# 0 0.53443f
C36 a_n1116_n597# 0 0.557987f
C37 w_n1374_n797# 0 15.1963f
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_62W3XE a_358_n500# a_158_n588# a_100_n500# a_n158_n500#
+ a_n358_n588# a_n100_n588# a_n550_n722# a_n416_n500#
X0 a_100_n500# a_n100_n588# a_n158_n500# a_n550_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X1 a_n158_n500# a_n358_n588# a_n416_n500# a_n550_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=1
X2 a_358_n500# a_158_n588# a_100_n500# a_n550_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=1
C0 a_n358_n588# a_n158_n500# 0.112293f
C1 a_n158_n500# a_n416_n500# 0.273876f
C2 a_100_n500# a_n158_n500# 0.273876f
C3 a_158_n588# a_358_n500# 0.112293f
C4 a_n100_n588# a_158_n588# 0.104496f
C5 a_158_n588# a_100_n500# 0.112293f
C6 a_n100_n588# a_n358_n588# 0.104496f
C7 a_100_n500# a_358_n500# 0.273876f
C8 a_n100_n588# a_100_n500# 0.112293f
C9 a_n358_n588# a_n416_n500# 0.112293f
C10 a_n100_n588# a_n158_n500# 0.112293f
C11 a_358_n500# a_n550_n722# 0.553437f
C12 a_100_n500# a_n550_n722# 0.166296f
C13 a_n158_n500# a_n550_n722# 0.166296f
C14 a_n416_n500# a_n550_n722# 0.553437f
C15 a_158_n588# a_n550_n722# 0.651749f
C16 a_n100_n588# a_n550_n722# 0.588947f
C17 a_n358_n588# a_n550_n722# 0.651749f
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_EC8RE7 a_416_n500# a_n1364_n500# a_830_n588#
+ a_n1676_n722# a_n118_n500# a_1186_n588# a_n594_n588# a_238_n500# a_n1186_n500# a_652_n588#
+ a_1484_n500# a_n830_n500# a_n60_n588# a_950_n500# a_1008_n588# a_n416_n588# a_n1008_n500#
+ a_474_n588# a_n1484_n588# a_n652_n500# a_772_n500# a_n238_n588# a_296_n588# a_n474_n500#
+ a_1128_n500# a_n1306_n588# a_n950_n588# a_594_n500# a_n1542_n500# a_n296_n500# a_118_n588#
+ a_60_n500# a_1364_n588# a_n1128_n588# a_n772_n588#
X0 a_416_n500# a_296_n588# a_238_n500# a_n1676_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X1 a_n296_n500# a_n416_n588# a_n474_n500# a_n1676_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X2 a_1306_n500# a_1186_n588# a_1128_n500# a_n1676_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X3 a_n1364_n500# a_n1484_n588# a_n1542_n500# a_n1676_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=0.6
X4 a_238_n500# a_118_n588# a_60_n500# a_n1676_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X5 a_1128_n500# a_1008_n588# a_950_n500# a_n1676_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X6 a_n1186_n500# a_n1306_n588# a_n1364_n500# a_n1676_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X7 a_772_n500# a_652_n588# a_594_n500# a_n1676_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X8 a_n118_n500# a_n238_n588# a_n296_n500# a_n1676_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X9 a_n652_n500# a_n772_n588# a_n830_n500# a_n1676_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X10 a_n1008_n500# a_n1128_n588# a_n1186_n500# a_n1676_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X11 a_594_n500# a_474_n588# a_416_n500# a_n1676_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X12 a_60_n500# a_n60_n588# a_n118_n500# a_n1676_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X13 a_1484_n500# a_1364_n588# a_1306_n500# a_n1676_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=0.6
X14 a_950_n500# a_830_n588# a_772_n500# a_n1676_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X15 a_n830_n500# a_n950_n588# a_n1008_n500# a_n1676_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X16 a_n474_n500# a_n594_n588# a_n652_n500# a_n1676_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
C0 a_416_n500# a_238_n500# 0.396241f
C1 a_594_n500# a_772_n500# 0.396241f
C2 a_n1128_n588# a_n1306_n588# 0.104496f
C3 a_652_n588# a_830_n588# 0.104496f
C4 a_n772_n588# a_n950_n588# 0.104496f
C5 a_1306_n500# a_1128_n500# 0.396241f
C6 a_n652_n500# a_n474_n500# 0.396241f
C7 a_n1128_n588# a_n950_n588# 0.104496f
C8 a_n238_n588# a_n60_n588# 0.104496f
C9 a_830_n588# a_1008_n588# 0.104496f
C10 a_n416_n588# a_n238_n588# 0.104496f
C11 a_652_n588# a_474_n588# 0.104496f
C12 a_n296_n500# a_n474_n500# 0.396241f
C13 a_n830_n500# a_n652_n500# 0.396241f
C14 a_n772_n588# a_n594_n588# 0.104496f
C15 a_772_n500# a_950_n500# 0.396241f
C16 a_60_n500# a_238_n500# 0.396241f
C17 a_1364_n588# a_1186_n588# 0.104496f
C18 a_n296_n500# a_n118_n500# 0.396241f
C19 a_118_n588# a_n60_n588# 0.104496f
C20 a_n1186_n500# a_n1008_n500# 0.396241f
C21 a_296_n588# a_474_n588# 0.104496f
C22 a_1008_n588# a_1186_n588# 0.104496f
C23 a_n830_n500# a_n1008_n500# 0.396241f
C24 a_118_n588# a_296_n588# 0.104496f
C25 a_n594_n588# a_n416_n588# 0.104496f
C26 a_n1542_n500# a_n1364_n500# 0.396241f
C27 a_1128_n500# a_950_n500# 0.396241f
C28 a_594_n500# a_416_n500# 0.396241f
C29 a_1306_n500# a_1484_n500# 0.396241f
C30 a_n1484_n588# a_n1306_n588# 0.104496f
C31 a_n1186_n500# a_n1364_n500# 0.396241f
C32 a_n118_n500# a_60_n500# 0.396241f
C33 a_1484_n500# a_n1676_n722# 0.532243f
C34 a_1306_n500# a_n1676_n722# 0.123908f
C35 a_1128_n500# a_n1676_n722# 0.123908f
C36 a_950_n500# a_n1676_n722# 0.123908f
C37 a_772_n500# a_n1676_n722# 0.123908f
C38 a_594_n500# a_n1676_n722# 0.123908f
C39 a_416_n500# a_n1676_n722# 0.123908f
C40 a_238_n500# a_n1676_n722# 0.123908f
C41 a_60_n500# a_n1676_n722# 0.123908f
C42 a_n118_n500# a_n1676_n722# 0.123908f
C43 a_n296_n500# a_n1676_n722# 0.123908f
C44 a_n474_n500# a_n1676_n722# 0.123908f
C45 a_n652_n500# a_n1676_n722# 0.123908f
C46 a_n830_n500# a_n1676_n722# 0.123908f
C47 a_n1008_n500# a_n1676_n722# 0.123908f
C48 a_n1186_n500# a_n1676_n722# 0.123908f
C49 a_n1364_n500# a_n1676_n722# 0.123908f
C50 a_n1542_n500# a_n1676_n722# 0.532243f
C51 a_1364_n588# a_n1676_n722# 0.427362f
C52 a_1186_n588# a_n1676_n722# 0.364559f
C53 a_1008_n588# a_n1676_n722# 0.364559f
C54 a_830_n588# a_n1676_n722# 0.364559f
C55 a_652_n588# a_n1676_n722# 0.364559f
C56 a_474_n588# a_n1676_n722# 0.364559f
C57 a_296_n588# a_n1676_n722# 0.364559f
C58 a_118_n588# a_n1676_n722# 0.364559f
C59 a_n60_n588# a_n1676_n722# 0.364559f
C60 a_n238_n588# a_n1676_n722# 0.364559f
C61 a_n416_n588# a_n1676_n722# 0.364559f
C62 a_n594_n588# a_n1676_n722# 0.364559f
C63 a_n772_n588# a_n1676_n722# 0.364559f
C64 a_n950_n588# a_n1676_n722# 0.364559f
C65 a_n1128_n588# a_n1676_n722# 0.364559f
C66 a_n1306_n588# a_n1676_n722# 0.364559f
C67 a_n1484_n588# a_n1676_n722# 0.427362f
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_Y9J9EP a_n358_n597# a_358_n500# a_n100_n597#
+ a_100_n500# a_n158_n500# 0 a_158_n597# w_n616_n797# a_n416_n500#
X0 a_358_n500# a_158_n597# a_100_n500# w_n616_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=1
X1 a_100_n500# a_n100_n597# a_n158_n500# w_n616_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X2 a_n158_n500# a_n358_n597# a_n416_n500# w_n616_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=1
C0 a_n358_n597# a_n158_n500# 0.112293f
C1 a_n358_n597# w_n616_n797# 0.386009f
C2 a_100_n500# a_n100_n597# 0.112293f
C3 a_n158_n500# a_n100_n597# 0.112293f
C4 w_n616_n797# a_n100_n597# 0.34322f
C5 a_n158_n500# a_n416_n500# 0.273876f
C6 a_100_n500# a_n158_n500# 0.273876f
C7 w_n616_n797# a_n416_n500# 0.305447f
C8 a_158_n597# a_n100_n597# 0.109462f
C9 a_100_n500# a_158_n597# 0.112293f
C10 a_100_n500# a_358_n500# 0.273876f
C11 a_158_n597# w_n616_n797# 0.386009f
C12 a_n358_n597# a_n100_n597# 0.109462f
C13 w_n616_n797# a_358_n500# 0.305447f
C14 a_n358_n597# a_n416_n500# 0.112293f
C15 a_158_n597# a_358_n500# 0.112293f
C16 a_358_n500# 0 0.249778f
C17 a_100_n500# 0 0.144174f
C18 a_n158_n500# 0 0.144174f
C19 a_n416_n500# 0 0.249778f
C20 a_158_n597# 0 0.283364f
C21 a_n100_n597# 0 0.259807f
C22 a_n358_n597# 0 0.283364f
C23 w_n616_n797# 0 7.15269f
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_QZVU2P a_2974_n500# a_2116_n500# a_n458_n500#
+ a_n2974_n588# a_n3032_n500# a_n2116_n588# a_n400_n588# a_1258_n500# a_2174_n588#
+ a_n2174_n500# a_n3166_n722# a_n1258_n588# a_1316_n588# a_458_n588# a_400_n500# a_n1316_n500#
X0 a_n2174_n500# a_n2974_n588# a_n3032_n500# a_n3166_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=4
X1 a_1258_n500# a_458_n588# a_400_n500# a_n3166_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X2 a_n1316_n500# a_n2116_n588# a_n2174_n500# a_n3166_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X3 a_n458_n500# a_n1258_n588# a_n1316_n500# a_n3166_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X4 a_2116_n500# a_1316_n588# a_1258_n500# a_n3166_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X5 a_2974_n500# a_2174_n588# a_2116_n500# a_n3166_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=4
X6 a_400_n500# a_n400_n588# a_n458_n500# a_n3166_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
C0 a_n458_n500# a_n400_n588# 0.196631f
C1 a_1316_n588# a_2116_n500# 0.196631f
C2 a_n2974_n588# a_n3032_n500# 0.196631f
C3 a_1316_n588# a_2174_n588# 0.104496f
C4 a_458_n588# a_n400_n588# 0.104496f
C5 a_400_n500# a_n400_n588# 0.196631f
C6 a_n2974_n588# a_n2174_n500# 0.196631f
C7 a_1316_n588# a_458_n588# 0.104496f
C8 a_458_n588# a_400_n500# 0.196631f
C9 a_n2974_n588# a_n2116_n588# 0.104496f
C10 a_2174_n588# a_2974_n500# 0.196631f
C11 a_n1258_n588# a_n1316_n500# 0.196631f
C12 a_2174_n588# a_2116_n500# 0.196631f
C13 a_n1258_n588# a_n458_n500# 0.196631f
C14 a_1316_n588# a_1258_n500# 0.196631f
C15 a_458_n588# a_1258_n500# 0.196631f
C16 a_n1258_n588# a_n400_n588# 0.104496f
C17 a_n1316_n500# a_n2116_n588# 0.196631f
C18 a_n2174_n500# a_n2116_n588# 0.196631f
C19 a_n1258_n588# a_n2116_n588# 0.104496f
C20 a_2974_n500# a_n3166_n722# 0.629934f
C21 a_2116_n500# a_n3166_n722# 0.319289f
C22 a_1258_n500# a_n3166_n722# 0.319289f
C23 a_400_n500# a_n3166_n722# 0.319289f
C24 a_n458_n500# a_n3166_n722# 0.319289f
C25 a_n1316_n500# a_n3166_n722# 0.319289f
C26 a_n2174_n500# a_n3166_n722# 0.319289f
C27 a_n3032_n500# a_n3166_n722# 0.629934f
C28 a_2174_n588# a_n3166_n722# 2.33466f
C29 a_1316_n588# a_n3166_n722# 2.27186f
C30 a_458_n588# a_n3166_n722# 2.27186f
C31 a_n400_n588# a_n3166_n722# 2.27186f
C32 a_n1258_n588# a_n3166_n722# 2.27186f
C33 a_n2116_n588# a_n3166_n722# 2.27186f
C34 a_n2974_n588# a_n3166_n722# 2.33466f
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_7JLQGA a_416_n500# a_n238_n597# a_n118_n500#
+ a_296_n597# a_238_n500# a_n830_n500# a_118_n597# a_n652_n500# a_n772_n597# w_n1030_n797#
+ a_772_n500# 0 a_n474_n500# a_n594_n597# a_652_n597# a_594_n500# a_n60_n597# a_n296_n500#
+ a_60_n500# a_n416_n597# a_474_n597#
X0 a_n474_n500# a_n594_n597# a_n652_n500# w_n1030_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X1 a_416_n500# a_296_n597# a_238_n500# w_n1030_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X2 a_n296_n500# a_n416_n597# a_n474_n500# w_n1030_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X3 a_238_n500# a_118_n597# a_60_n500# w_n1030_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X4 a_772_n500# a_652_n597# a_594_n500# w_n1030_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=0.6
X5 a_n118_n500# a_n238_n597# a_n296_n500# w_n1030_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X6 a_n652_n500# a_n772_n597# a_n830_n500# w_n1030_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=0.6
X7 a_594_n500# a_474_n597# a_416_n500# w_n1030_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X8 a_60_n500# a_n60_n597# a_n118_n500# w_n1030_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
C0 a_n296_n500# a_n474_n500# 0.396241f
C1 w_n1030_n797# a_n772_n597# 0.26725f
C2 a_594_n500# a_772_n500# 0.396241f
C3 a_n296_n500# a_n118_n500# 0.396241f
C4 w_n1030_n797# a_118_n597# 0.224461f
C5 a_652_n597# a_474_n597# 0.109462f
C6 w_n1030_n797# a_n830_n500# 0.305456f
C7 a_n830_n500# a_n652_n500# 0.396241f
C8 a_n60_n597# a_n238_n597# 0.109462f
C9 w_n1030_n797# a_n416_n597# 0.224461f
C10 w_n1030_n797# a_296_n597# 0.224461f
C11 a_n474_n500# a_n652_n500# 0.396241f
C12 a_n594_n597# a_n772_n597# 0.109462f
C13 a_416_n500# a_594_n500# 0.396241f
C14 a_n238_n597# a_n416_n597# 0.109462f
C15 a_n60_n597# a_118_n597# 0.109462f
C16 a_474_n597# a_296_n597# 0.109462f
C17 a_238_n500# a_60_n500# 0.396241f
C18 a_n594_n597# a_n416_n597# 0.109462f
C19 w_n1030_n797# a_n238_n597# 0.224461f
C20 a_60_n500# a_n118_n500# 0.396241f
C21 w_n1030_n797# a_474_n597# 0.224461f
C22 a_118_n597# a_296_n597# 0.109462f
C23 a_416_n500# a_238_n500# 0.396241f
C24 w_n1030_n797# a_652_n597# 0.26725f
C25 w_n1030_n797# a_n594_n597# 0.224461f
C26 w_n1030_n797# a_772_n500# 0.305456f
C27 w_n1030_n797# a_n60_n597# 0.224461f
C28 a_772_n500# 0 0.228576f
C29 a_594_n500# 0 0.101769f
C30 a_416_n500# 0 0.101769f
C31 a_238_n500# 0 0.101769f
C32 a_60_n500# 0 0.101769f
C33 a_n118_n500# 0 0.101769f
C34 a_n296_n500# 0 0.101769f
C35 a_n474_n500# 0 0.101769f
C36 a_n652_n500# 0 0.101769f
C37 a_n830_n500# 0 0.228576f
C38 a_652_n597# 0 0.173515f
C39 a_474_n597# 0 0.149958f
C40 a_296_n597# 0 0.149958f
C41 a_118_n597# 0 0.149958f
C42 a_n60_n597# 0 0.149958f
C43 a_n238_n597# 0 0.149958f
C44 a_n416_n597# 0 0.149958f
C45 a_n594_n597# 0 0.149958f
C46 a_n772_n597# 0 0.173515f
C47 w_n1030_n797# 0 11.5938f
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_3DCHX4 a_n1687_n1687# a_n3287_n557# a_29_599#
+ a_1629_1781# a_1687_n2869# a_n3287_n1713# a_3287_n2843# a_3287_n531# a_n1629_1755#
+ a_1687_n1713# a_n1687_n531# a_n1687_625# a_29_n2869# a_n3345_n2843# a_n1687_n2843#
+ a_1687_1755# a_29_n1713# a_n29_n531# a_3287_1781# a_29_1755# a_n29_n1687# a_n3345_625#
+ a_n3479_n3003# a_n1687_1781# a_1629_n1687# a_n29_625# a_n3287_1755# a_n1629_n557#
+ a_3287_625# a_1687_599# a_n3345_n531# a_1629_n531# a_n3287_599# a_n1629_n2869# a_3287_n1687#
+ a_n29_1781# a_1629_625# a_n29_n2843# a_1687_n557# a_n1629_n1713# a_n1629_599# a_1629_n2843#
+ a_29_n557# a_n3287_n2869# a_n3345_n1687# a_n3345_1781#
X0 a_n1687_625# a_n3287_599# a_n3345_625# a_n3479_n3003# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=8
X1 a_1629_n531# a_29_n557# a_n29_n531# a_n3479_n3003# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=8
X2 a_1629_1781# a_29_1755# a_n29_1781# a_n3479_n3003# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=8
X3 a_3287_n531# a_1687_n557# a_1629_n531# a_n3479_n3003# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=8
X4 a_3287_1781# a_1687_1755# a_1629_1781# a_n3479_n3003# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=8
X5 a_n1687_n531# a_n3287_n557# a_n3345_n531# a_n3479_n3003# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=8
X6 a_n29_625# a_n1629_599# a_n1687_625# a_n3479_n3003# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=8
X7 a_n1687_n1687# a_n3287_n1713# a_n3345_n1687# a_n3479_n3003# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=8
X8 a_n1687_1781# a_n3287_1755# a_n3345_1781# a_n3479_n3003# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=8
X9 a_1629_n1687# a_29_n1713# a_n29_n1687# a_n3479_n3003# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=8
X10 a_n1687_n2843# a_n3287_n2869# a_n3345_n2843# a_n3479_n3003# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=8
X11 a_3287_n1687# a_1687_n1713# a_1629_n1687# a_n3479_n3003# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=8
X12 a_1629_n2843# a_29_n2869# a_n29_n2843# a_n3479_n3003# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=8
X13 a_1629_625# a_29_599# a_n29_625# a_n3479_n3003# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=8
X14 a_3287_625# a_1687_599# a_1629_625# a_n3479_n3003# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=8
X15 a_n29_n531# a_n1629_n557# a_n1687_n531# a_n3479_n3003# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=8
X16 a_3287_n2843# a_1687_n2869# a_1629_n2843# a_n3479_n3003# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=8
X17 a_n29_1781# a_n1629_1755# a_n1687_1781# a_n3479_n3003# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=8
X18 a_n29_n1687# a_n1629_n1713# a_n1687_n1687# a_n3479_n3003# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=8
X19 a_n29_n2843# a_n1629_n2869# a_n1687_n2843# a_n3479_n3003# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=8
C0 a_29_599# a_1629_625# 0.216528f
C1 a_n3345_n531# a_n3287_n557# 0.216528f
C2 a_1687_599# a_1629_625# 0.216528f
C3 a_n3287_599# a_n3287_n557# 0.981682f
C4 a_n1687_625# a_n3287_599# 0.216528f
C5 a_n1629_n2869# a_n1687_n2843# 0.216528f
C6 a_n1629_n557# a_n1629_n1713# 0.981682f
C7 a_1629_1781# a_1687_1755# 0.216528f
C8 a_29_n2869# a_n29_n2843# 0.216528f
C9 a_1629_n2843# a_1687_n2869# 0.216528f
C10 a_29_n557# a_29_n1713# 0.981682f
C11 a_n3287_n2869# a_n1687_n2843# 0.216528f
C12 a_3287_1781# a_1687_1755# 0.216528f
C13 a_1687_n557# a_1687_n1713# 0.981682f
C14 a_29_n1713# a_1629_n1687# 0.216528f
C15 a_n1629_n2869# a_n1629_n1713# 0.981682f
C16 a_1687_n557# a_3287_n531# 0.216528f
C17 a_29_n557# a_29_599# 0.981682f
C18 a_n1629_599# a_n29_625# 0.216528f
C19 a_n1629_1755# a_n29_1781# 0.216528f
C20 a_n3287_1755# a_n3345_1781# 0.216528f
C21 a_29_n557# a_1629_n531# 0.216528f
C22 a_3287_625# a_1687_599# 0.216528f
C23 a_n3287_n1713# a_n3287_n557# 0.981682f
C24 a_n29_n1687# a_n1629_n1713# 0.216528f
C25 a_n1629_n2869# a_n29_n2843# 0.216528f
C26 a_29_n1713# a_n29_n1687# 0.216528f
C27 a_n1687_1781# a_n3287_1755# 0.216528f
C28 a_3287_n2843# a_1687_n2869# 0.216528f
C29 a_n1687_n1687# a_n1629_n1713# 0.216528f
C30 a_n3345_n1687# a_n3287_n1713# 0.216528f
C31 a_1687_n1713# a_1629_n1687# 0.216528f
C32 a_1687_n2869# a_1687_n1713# 0.981682f
C33 a_29_1755# a_29_599# 0.981682f
C34 a_n1629_n557# a_n29_n531# 0.216528f
C35 a_29_n557# a_n29_n531# 0.216528f
C36 a_n1629_1755# a_n1687_1781# 0.216528f
C37 a_29_599# a_n29_625# 0.216528f
C38 a_n3287_n2869# a_n3287_n1713# 0.981682f
C39 a_29_1755# a_n29_1781# 0.216528f
C40 a_n1629_n557# a_n1687_n531# 0.216528f
C41 a_n1687_n531# a_n3287_n557# 0.216528f
C42 a_1629_n2843# a_29_n2869# 0.216528f
C43 a_n3345_n2843# a_n3287_n2869# 0.216528f
C44 a_n3287_1755# a_n3287_599# 0.981682f
C45 a_n1629_1755# a_n1629_599# 0.981682f
C46 a_1687_599# a_1687_1755# 0.981682f
C47 a_29_n1713# a_29_n2869# 0.981682f
C48 a_n1629_n557# a_n1629_599# 0.981682f
C49 a_3287_n1687# a_1687_n1713# 0.216528f
C50 a_29_1755# a_1629_1781# 0.216528f
C51 a_1687_n557# a_1687_599# 0.981682f
C52 a_n1687_625# a_n1629_599# 0.216528f
C53 a_n1687_n1687# a_n3287_n1713# 0.216528f
C54 a_1687_n557# a_1629_n531# 0.216528f
C55 a_n3287_599# a_n3345_625# 0.216528f
C56 a_3287_n2843# a_n3479_n3003# 0.706465f
C57 a_1629_n2843# a_n3479_n3003# 0.482688f
C58 a_n29_n2843# a_n3479_n3003# 0.482688f
C59 a_n1687_n2843# a_n3479_n3003# 0.482688f
C60 a_n3345_n2843# a_n3479_n3003# 0.706465f
C61 a_1687_n2869# a_n3479_n3003# 2.64477f
C62 a_29_n2869# a_n3479_n3003# 2.6085f
C63 a_n1629_n2869# a_n3479_n3003# 2.6085f
C64 a_n3287_n2869# a_n3479_n3003# 2.64477f
C65 a_3287_n1687# a_n3479_n3003# 0.692968f
C66 a_1629_n1687# a_n3479_n3003# 0.469191f
C67 a_n29_n1687# a_n3479_n3003# 0.469191f
C68 a_n1687_n1687# a_n3479_n3003# 0.469191f
C69 a_n3345_n1687# a_n3479_n3003# 0.692968f
C70 a_1687_n1713# a_n3479_n3003# 2.19493f
C71 a_29_n1713# a_n3479_n3003# 2.15867f
C72 a_n1629_n1713# a_n3479_n3003# 2.15867f
C73 a_n3287_n1713# a_n3479_n3003# 2.19493f
C74 a_3287_n531# a_n3479_n3003# 0.692968f
C75 a_1629_n531# a_n3479_n3003# 0.469191f
C76 a_n29_n531# a_n3479_n3003# 0.469191f
C77 a_n1687_n531# a_n3479_n3003# 0.469191f
C78 a_n3345_n531# a_n3479_n3003# 0.692968f
C79 a_1687_n557# a_n3479_n3003# 2.19493f
C80 a_29_n557# a_n3479_n3003# 2.15867f
C81 a_n1629_n557# a_n3479_n3003# 2.15867f
C82 a_n3287_n557# a_n3479_n3003# 2.19493f
C83 a_3287_625# a_n3479_n3003# 0.692968f
C84 a_1629_625# a_n3479_n3003# 0.469191f
C85 a_n29_625# a_n3479_n3003# 0.469191f
C86 a_n1687_625# a_n3479_n3003# 0.469191f
C87 a_n3345_625# a_n3479_n3003# 0.692968f
C88 a_1687_599# a_n3479_n3003# 2.19493f
C89 a_29_599# a_n3479_n3003# 2.15867f
C90 a_n1629_599# a_n3479_n3003# 2.15867f
C91 a_n3287_599# a_n3479_n3003# 2.19493f
C92 a_3287_1781# a_n3479_n3003# 0.704885f
C93 a_1629_1781# a_n3479_n3003# 0.481108f
C94 a_n29_1781# a_n3479_n3003# 0.481108f
C95 a_n1687_1781# a_n3479_n3003# 0.481108f
C96 a_n3345_1781# a_n3479_n3003# 0.704885f
C97 a_1687_1755# a_n3479_n3003# 2.97499f
C98 a_29_1755# a_n3479_n3003# 2.93872f
C99 a_n1629_1755# a_n3479_n3003# 2.93872f
C100 a_n3287_1755# a_n3479_n3003# 2.97499f
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_75J6LY a_n3403_n597# a_5977_n500# a_5177_n597#
+ a_29_n597# a_n2603_n500# a_5119_n500# a_n6893_n500# a_3461_n597# a_3403_n500# a_n6035_n500#
+ a_n2545_n597# w_n7093_n797# a_n1745_n500# a_4319_n597# a_n6835_n597# a_2545_n500#
+ a_2603_n597# a_n5177_n500# a_n1687_n597# a_n4261_n597# a_n887_n500# 0 a_6835_n500#
+ a_n3461_n500# a_6035_n597# a_n5977_n597# a_n29_n500# a_n5119_n597# a_1687_n500#
+ a_1745_n597# a_n829_n597# a_4261_n500# a_887_n597# a_829_n500# a_n4319_n500#
X0 a_n6035_n500# a_n6835_n597# a_n6893_n500# w_n7093_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=4
X1 a_3403_n500# a_2603_n597# a_2545_n500# w_n7093_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X2 a_n29_n500# a_n829_n597# a_n887_n500# w_n7093_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X3 a_n5177_n500# a_n5977_n597# a_n6035_n500# w_n7093_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X4 a_2545_n500# a_1745_n597# a_1687_n500# w_n7093_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X5 a_4261_n500# a_3461_n597# a_3403_n500# w_n7093_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X6 a_n4319_n500# a_n5119_n597# a_n5177_n500# w_n7093_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X7 a_829_n500# a_29_n597# a_n29_n500# w_n7093_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X8 a_n2603_n500# a_n3403_n597# a_n3461_n500# w_n7093_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X9 a_1687_n500# a_887_n597# a_829_n500# w_n7093_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X10 a_6835_n500# a_6035_n597# a_5977_n500# w_n7093_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=4
X11 a_5119_n500# a_4319_n597# a_4261_n500# w_n7093_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X12 a_n3461_n500# a_n4261_n597# a_n4319_n500# w_n7093_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X13 a_n1745_n500# a_n2545_n597# a_n2603_n500# w_n7093_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X14 a_5977_n500# a_5177_n597# a_5119_n500# w_n7093_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X15 a_n887_n500# a_n1687_n597# a_n1745_n500# w_n7093_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
C0 a_n5177_n500# a_n5119_n597# 0.196631f
C1 a_4319_n597# a_5177_n597# 0.109462f
C2 a_6035_n597# a_5977_n500# 0.196631f
C3 a_n29_n500# a_29_n597# 0.196631f
C4 a_1745_n597# a_2545_n500# 0.196631f
C5 w_n7093_n797# a_n3403_n597# 1.23391f
C6 a_4261_n500# a_3461_n597# 0.196631f
C7 a_n3403_n597# a_n2603_n500# 0.196631f
C8 a_n5119_n597# a_n4319_n500# 0.196631f
C9 a_4319_n597# a_3461_n597# 0.109462f
C10 a_5119_n500# a_5177_n597# 0.196631f
C11 w_n7093_n797# a_5177_n597# 1.23391f
C12 a_1745_n597# a_2603_n597# 0.109462f
C13 a_n6835_n597# a_n5977_n597# 0.109462f
C14 a_n6835_n597# a_n6893_n500# 0.196631f
C15 w_n7093_n797# a_3461_n597# 1.23391f
C16 a_887_n597# a_29_n597# 0.109462f
C17 a_6035_n597# a_6835_n500# 0.196631f
C18 a_n5119_n597# a_n5977_n597# 0.109462f
C19 w_n7093_n797# a_n6835_n597# 1.2767f
C20 a_n6035_n500# a_n5977_n597# 0.196631f
C21 w_n7093_n797# a_6035_n597# 1.2767f
C22 a_n5177_n500# a_n5977_n597# 0.196631f
C23 w_n7093_n797# a_n2545_n597# 1.23391f
C24 w_n7093_n797# a_n829_n597# 1.23391f
C25 a_n5119_n597# a_n4261_n597# 0.109462f
C26 a_n2545_n597# a_n2603_n500# 0.196631f
C27 a_1745_n597# a_887_n597# 0.109462f
C28 a_n4261_n597# a_n3461_n500# 0.196631f
C29 a_n3403_n597# a_n2545_n597# 0.109462f
C30 w_n7093_n797# a_2603_n597# 1.23391f
C31 w_n7093_n797# a_n5119_n597# 1.23391f
C32 a_6035_n597# a_5177_n597# 0.109462f
C33 w_n7093_n797# a_29_n597# 1.23391f
C34 a_n4261_n597# a_n4319_n500# 0.196631f
C35 a_n829_n597# a_n887_n500# 0.196631f
C36 a_n3403_n597# a_n3461_n500# 0.196631f
C37 a_829_n500# a_29_n597# 0.196631f
C38 w_n7093_n797# a_n1687_n597# 1.23391f
C39 a_n1745_n500# a_n2545_n597# 0.196631f
C40 w_n7093_n797# a_1745_n597# 1.23391f
C41 w_n7093_n797# a_887_n597# 1.23391f
C42 a_4261_n500# a_4319_n597# 0.196631f
C43 a_2603_n597# a_3461_n597# 0.109462f
C44 a_829_n500# a_887_n597# 0.196631f
C45 a_n887_n500# a_n1687_n597# 0.196631f
C46 a_3461_n597# a_3403_n500# 0.196631f
C47 a_5177_n597# a_5977_n500# 0.196631f
C48 a_2603_n597# a_2545_n500# 0.196631f
C49 w_n7093_n797# a_n5977_n597# 1.23391f
C50 w_n7093_n797# a_n6893_n500# 0.305424f
C51 a_4319_n597# a_5119_n500# 0.196631f
C52 w_n7093_n797# a_4319_n597# 1.23391f
C53 a_1745_n597# a_1687_n500# 0.196631f
C54 a_n1745_n500# a_n1687_n597# 0.196631f
C55 a_n6835_n597# a_n6035_n500# 0.196631f
C56 a_n829_n597# a_n29_n500# 0.196631f
C57 a_1687_n500# a_887_n597# 0.196631f
C58 w_n7093_n797# a_n4261_n597# 1.23391f
C59 w_n7093_n797# a_6835_n500# 0.305424f
C60 a_n829_n597# a_29_n597# 0.109462f
C61 a_n4261_n597# a_n3403_n597# 0.109462f
C62 a_n2545_n597# a_n1687_n597# 0.109462f
C63 a_2603_n597# a_3403_n500# 0.196631f
C64 a_n829_n597# a_n1687_n597# 0.109462f
C65 a_6835_n500# 0 0.326298f
C66 a_5977_n500# 0 0.297214f
C67 a_5119_n500# 0 0.297214f
C68 a_4261_n500# 0 0.297214f
C69 a_3403_n500# 0 0.297214f
C70 a_2545_n500# 0 0.297214f
C71 a_1687_n500# 0 0.297214f
C72 a_829_n500# 0 0.297214f
C73 a_n29_n500# 0 0.297214f
C74 a_n887_n500# 0 0.297214f
C75 a_n1745_n500# 0 0.297214f
C76 a_n2603_n500# 0 0.297214f
C77 a_n3461_n500# 0 0.297214f
C78 a_n4319_n500# 0 0.297214f
C79 a_n5177_n500# 0 0.297214f
C80 a_n6035_n500# 0 0.297214f
C81 a_n6893_n500# 0 0.326298f
C82 a_6035_n597# 0 1.10723f
C83 a_5177_n597# 0 1.08368f
C84 a_4319_n597# 0 1.08368f
C85 a_3461_n597# 0 1.08368f
C86 a_2603_n597# 0 1.08368f
C87 a_1745_n597# 0 1.08368f
C88 a_887_n597# 0 1.08368f
C89 a_29_n597# 0 1.08368f
C90 a_n829_n597# 0 1.08368f
C91 a_n1687_n597# 0 1.08368f
C92 a_n2545_n597# 0 1.08368f
C93 a_n3403_n597# 0 1.08368f
C94 a_n4261_n597# 0 1.08368f
C95 a_n5119_n597# 0 1.08368f
C96 a_n5977_n597# 0 1.08368f
C97 a_n6835_n597# 0 1.10723f
C98 w_n7093_n797# 0 75.727005f
.ends

.subckt ibias_gen ibias0 itest ibias1 ibg_200n vbg_1v2 ve m1_7189_119# m1_1897_119#
+ vstart vr isrc_sel_b m1_5677_119# vp1 m1_1141_119# ena_b vp ena m1_385_119# m1_2653_119#
+ m1_4165_119# isrc_sel vn0 avdd avss m1_763_7518# vp0 vn1
Xsky130_fd_pr__nfet_g5v0d10v5_XZ4X25_0 isrc_sel_b ena_b isrc_sel avss ena_b vn1 avss
+ avss avss vn0 sky130_fd_pr__nfet_g5v0d10v5_XZ4X25
Xsky130_fd_pr__pfet_g5v0d10v5_Y9S9FP_0 avdd ena vp0 isrc_sel vp1 avss avdd avdd vp
+ ena avdd ena isrc_sel_b sky130_fd_pr__pfet_g5v0d10v5_Y9S9FP
Xsky130_fd_pr__nfet_g5v0d10v5_62W3XE_0 avss isrc_sel isrc_sel_b ena_b ena avss avss
+ avss sky130_fd_pr__nfet_g5v0d10v5_62W3XE
Xsky130_fd_pr__nfet_g5v0d10v5_EC8RE7_1 vp0 vstart isrc_sel avss vn0 isrc_sel vbg_1v2
+ vn0 vn0 avss ibg_200n vn0 vbg_1v2 vp1 avss vbg_1v2 vstart isrc_sel_b vbg_1v2 vstart
+ vp vbg_1v2 avss vn0 vn1 vbg_1v2 vbg_1v2 vp vn0 vstart vbg_1v2 vstart ena vbg_1v2
+ vbg_1v2 sky130_fd_pr__nfet_g5v0d10v5_EC8RE7
Xsky130_fd_pr__pfet_g5v0d10v5_Y9J9EP_0 ena avdd avdd isrc_sel_b ena_b avss isrc_sel
+ avdd avdd sky130_fd_pr__pfet_g5v0d10v5_Y9J9EP
Xsky130_fd_pr__nfet_g5v0d10v5_QZVU2P_1 avss vr ve avss avss vn0 avss vp0 avss ve avss
+ vn0 vn0 vn0 vr vn0 sky130_fd_pr__nfet_g5v0d10v5_QZVU2P
Xsky130_fd_pr__res_xhigh_po_1p41_DVQADA_0 m1_4165_119# m1_3409_119# m1_3409_119# m1_5299_7518#
+ m1_1519_7518# m1_385_119# m1_2653_119# m1_385_119# m1_2653_119# m1_6433_119# m1_1897_119#
+ avss m1_6055_7518# m1_3787_7518# m1_2275_7518# m1_1519_7518# m1_6055_7518# m1_4165_119#
+ m1_5299_7518# m1_763_7518# m1_4921_119# m1_763_7518# m1_7189_119# m1_4543_7518#
+ m1_1897_119# m1_7189_119# m1_3031_7518# m1_6811_7518# m1_4921_119# m1_5677_119#
+ m1_5677_119# m1_6811_7518# m1_3031_7518# m1_3787_7518# m1_1141_119# avss m1_4543_7518#
+ m1_1141_119# m1_6433_119# vr m1_2275_7518# sky130_fd_pr__res_xhigh_po_1p41_DVQADA
Xsky130_fd_pr__pfet_g5v0d10v5_7JLQGA_0 vn1 isrc_sel vp avdd vp1 vstart isrc_sel_b
+ sky130_fd_pr__pfet_g5v0d10v5_7JLQGA_0/a_n652_n500# ena_b avdd ibg_200n avss avdd
+ isrc_sel ena_b sky130_fd_pr__pfet_g5v0d10v5_7JLQGA_0/a_594_n500# avdd vp0 vp avdd
+ isrc_sel_b sky130_fd_pr__pfet_g5v0d10v5_7JLQGA
Xsky130_fd_pr__nfet_g5v0d10v5_3DCHX4_0 avss avss vn1 avss avss avss avss avss vn1
+ avss avss avss vn1 avss avss avss vn1 vn1 avss vn1 vp1 avss avss avss avss vp1 avss
+ vn1 avss avss avss avss avss vn1 avss vp1 avss vp1 avss vn1 vn1 avss vn1 avss avss
+ avss sky130_fd_pr__nfet_g5v0d10v5_3DCHX4
Xsky130_fd_pr__pfet_g5v0d10v5_75J6LY_0 vp0 avdd vp vp vp0 ibias1 avdd vp1 vp1 avdd
+ vp0 avdd avdd vp avdd avdd vp1 vn0 avdd avdd avdd avss avdd avdd avdd vp0 ibias0
+ vp0 itest vp vp avdd vp avdd avdd sky130_fd_pr__pfet_g5v0d10v5_75J6LY
C0 avdd vn1 0.262267f
C1 ibg_200n ena_b 0.390945f
C2 vn0 ena_b 0.266557f
C3 vn0 isrc_sel_b 0.143624f
C4 vbg_1v2 vstart 1.118679f
C5 vn1 vp1 3.923848f
C6 vp0 isrc_sel 0.934617f
C7 vp0 vn0 1.62642f
C8 vp ena_b 0.254339f
C9 vp isrc_sel_b 0.469384f
C10 avdd ena_b 2.027189f
C11 isrc_sel sky130_fd_pr__pfet_g5v0d10v5_7JLQGA_0/a_n652_n500# 0.214977f
C12 avdd isrc_sel_b 1.376188f
C13 vp1 ena_b 0.142844f
C14 vn1 ena_b 0.154982f
C15 vp0 vp 0.551044f
C16 vp1 isrc_sel_b 0.336179f
C17 vn1 isrc_sel_b 0.337926f
C18 vp0 avdd 5.945743f
C19 vn0 vstart 0.887914f
C20 vp0 vp1 0.638232f
C21 m1_6811_7518# vn0 0.355414f
C22 vp vstart 0.101897f
C23 avdd vstart 0.54807f
C24 ena_b isrc_sel_b 2.308393f
C25 vp0 ena_b 0.494665f
C26 vp0 isrc_sel_b 0.229707f
C27 vp ibias0 0.210362f
C28 avdd ibias0 0.268708f
C29 vn0 vr 1.46054f
C30 isrc_sel ena 0.721356f
C31 ibg_200n ena 0.132599f
C32 vn0 ena 0.137245f
C33 vp0 vstart 0.337717f
C34 vbg_1v2 vn0 0.956591f
C35 vp0 m1_6811_7518# 0.114722f
C36 vp ena 0.308627f
C37 avdd ena 2.021183f
C38 vn1 ena 0.265105f
C39 avdd vbg_1v2 0.157961f
C40 vn0 isrc_sel 0.128091f
C41 vp0 vr 0.268135f
C42 ena_b ena 0.934834f
C43 vn0 ve 0.624897f
C44 ena isrc_sel_b 1.263019f
C45 vp isrc_sel 0.95764f
C46 avdd isrc_sel 4.496557f
C47 vp0 ena 0.224792f
C48 avdd ibg_200n 0.389983f
C49 avdd vn0 0.685485f
C50 isrc_sel vp1 0.427275f
C51 vn1 isrc_sel 0.467679f
C52 vn1 vn0 0.500783f
C53 vp0 vbg_1v2 0.126912f
C54 sky130_fd_pr__pfet_g5v0d10v5_7JLQGA_0/a_594_n500# ena_b 0.167441f
C55 vp ibias1 0.19584f
C56 vp avdd 9.989226f
C57 vp0 m1_6055_7518# 0.130049f
C58 vp vp1 1.225315f
C59 isrc_sel ena_b 0.867415f
C60 vp itest 0.210886f
C61 avdd vp1 3.235997f
C62 isrc_sel isrc_sel_b 1.70543f
C63 ena_b avss 3.288525f
C64 ibias1 avss 0.327614f
C65 itest avss 0.328668f
C66 ibias0 avss 0.329553f
C67 vp1 avss 6.166458f
C68 vn1 avss 36.535187f
C69 sky130_fd_pr__pfet_g5v0d10v5_7JLQGA_0/a_594_n500# avss 0.101769f
C70 sky130_fd_pr__pfet_g5v0d10v5_7JLQGA_0/a_n652_n500# avss 0.101769f
C71 vr avss 2.928733f
C72 m1_7189_119# avss 1.272288f
C73 m1_6811_7518# avss 0.981981f
C74 m1_6433_119# avss 0.979081f
C75 m1_6055_7518# avss 0.974485f
C76 m1_5677_119# avss 0.975689f
C77 m1_5299_7518# avss 0.974316f
C78 m1_4921_119# avss 0.975688f
C79 m1_4543_7518# avss 0.977415f
C80 m1_4165_119# avss 0.975689f
C81 m1_3787_7518# avss 0.976793f
C82 m1_3409_119# avss 0.975688f
C83 m1_3031_7518# avss 0.974316f
C84 m1_2653_119# avss 0.975689f
C85 m1_2275_7518# avss 0.975664f
C86 m1_1897_119# avss 0.975689f
C87 m1_1519_7518# avss 0.988117f
C88 m1_1141_119# avss 0.975771f
C89 m1_763_7518# avss 0.989193f
C90 m1_385_119# avss 1.244357f
C91 ve avss 1.524327f
C92 avdd avss 0.133453p
C93 ibg_200n avss 0.758831f
C94 sky130_fd_pr__nfet_g5v0d10v5_EC8RE7_1/a_1306_n500# avss 0.1558f $ **FLOATING
C95 vp avss 6.160111f
C96 vp0 avss 7.048689f
C97 vstart avss 1.070337f
C98 vn0 avss 18.357258f
C99 ena avss 2.928483f
C100 isrc_sel avss 4.333301f
C101 vbg_1v2 avss 4.502666f
C102 isrc_sel_b avss 3.295646f
.ends

.subckt sky130_fd_pr__rf_pnp_05v5_W0p68L0p68 Base Collector Emitter avss m=1
X0 Collector Base Emitter avss sky130_fd_pr__pnp_05v5_W0p68L0p68
**devattr s=18496,544
C0 Emitter Base 0.243586f
C1 Emitter Collector 0.105343f
C2 Base Collector 0.495333f
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_T82T27 a_1629_47# a_1687_21# a_n1687_47# a_4945_n309#
+ a_n1629_n335# a_n5137_n469# a_n4945_n335# a_n29_47# a_29_21# a_n3287_21# a_1687_n335#
+ a_3287_n309# a_n5003_n309# a_29_n335# a_n1687_n309# a_n5003_47# a_n4945_21# a_n3287_n335#
+ a_n1629_21# a_3345_21# a_n29_n309# a_3287_47# a_n3345_47# a_3345_n335# a_n3345_n309#
+ a_1629_n309# a_4945_47#
X0 a_1629_47# a_29_21# a_n29_47# a_n5137_n469# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1 a_n1687_47# a_n3287_21# a_n3345_47# a_n5137_n469# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X2 a_4945_47# a_3345_21# a_3287_47# a_n5137_n469# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=8
X3 a_1629_n309# a_29_n335# a_n29_n309# a_n5137_n469# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X4 a_n3345_n309# a_n4945_n335# a_n5003_n309# a_n5137_n469# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=8
X5 a_3287_n309# a_1687_n335# a_1629_n309# a_n5137_n469# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X6 a_n1687_n309# a_n3287_n335# a_n3345_n309# a_n5137_n469# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X7 a_n3345_47# a_n4945_21# a_n5003_47# a_n5137_n469# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=8
X8 a_n29_47# a_n1629_21# a_n1687_47# a_n5137_n469# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X9 a_4945_n309# a_3345_n335# a_3287_n309# a_n5137_n469# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=8
X10 a_3287_47# a_1687_21# a_1629_47# a_n5137_n469# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X11 a_n29_n309# a_n1629_n335# a_n1687_n309# a_n5137_n469# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
C0 a_n3287_21# a_n3287_n335# 1.09842f
C1 a_3345_n335# a_3345_21# 1.09842f
C2 a_29_n335# a_29_21# 1.09842f
C3 a_n4945_21# a_n4945_n335# 1.09842f
C4 a_1687_n335# a_1687_21# 1.09842f
C5 a_n1629_21# a_n1629_n335# 1.09842f
C6 a_4945_n309# a_n5137_n469# 0.157719f
C7 a_3287_n309# a_n5137_n469# 0.107936f
C8 a_1629_n309# a_n5137_n469# 0.107936f
C9 a_n29_n309# a_n5137_n469# 0.107936f
C10 a_n1687_n309# a_n5137_n469# 0.107936f
C11 a_n3345_n309# a_n5137_n469# 0.107936f
C12 a_n5003_n309# a_n5137_n469# 0.157719f
C13 a_3345_n335# a_n5137_n469# 2.63297f
C14 a_1687_n335# a_n5137_n469# 2.59671f
C15 a_29_n335# a_n5137_n469# 2.59671f
C16 a_n1629_n335# a_n5137_n469# 2.59671f
C17 a_n3287_n335# a_n5137_n469# 2.59671f
C18 a_n4945_n335# a_n5137_n469# 2.63297f
C19 a_4945_47# a_n5137_n469# 0.156139f
C20 a_3287_47# a_n5137_n469# 0.106356f
C21 a_1629_47# a_n5137_n469# 0.106356f
C22 a_n29_47# a_n5137_n469# 0.106356f
C23 a_n1687_47# a_n5137_n469# 0.106356f
C24 a_n3345_47# a_n5137_n469# 0.106356f
C25 a_n5003_47# a_n5137_n469# 0.156139f
C26 a_3345_21# a_n5137_n469# 2.87701f
C27 a_1687_21# a_n5137_n469# 2.84074f
C28 a_29_21# a_n5137_n469# 2.84074f
C29 a_n1629_21# a_n5137_n469# 2.84074f
C30 a_n3287_21# a_n5137_n469# 2.84074f
C31 a_n4945_21# a_n5137_n469# 2.87701f
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_3HV7M9 a_3345_n161# a_n1687_n64# a_n1629_n161#
+ a_n4945_n161# w_n5203_n362# a_1687_n161# a_n3345_n64# a_29_n161# 0 a_3287_n64# a_n29_n64#
+ a_n3287_n161# a_1629_n64# a_n5003_n64# a_4945_n64#
X0 a_n29_n64# a_n1629_n161# a_n1687_n64# w_n5203_n362# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1 a_n3345_n64# a_n4945_n161# a_n5003_n64# w_n5203_n362# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=8
X2 a_1629_n64# a_29_n161# a_n29_n64# w_n5203_n362# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X3 a_3287_n64# a_1687_n161# a_1629_n64# w_n5203_n362# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X4 a_4945_n64# a_3345_n161# a_3287_n64# w_n5203_n362# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=8
X5 a_n1687_n64# a_n3287_n161# a_n3345_n64# w_n5203_n362# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
C0 a_1687_n161# w_n5203_n362# 1.82215f
C1 a_n1629_n161# w_n5203_n362# 1.82215f
C2 a_n3287_n161# w_n5203_n362# 1.82215f
C3 a_3345_n161# w_n5203_n362# 1.84681f
C4 a_n4945_n161# w_n5203_n362# 1.84681f
C5 a_29_n161# w_n5203_n362# 1.82215f
C6 a_3345_n161# 0 1.7153f
C7 a_1687_n161# 0 1.70192f
C8 a_29_n161# 0 1.70192f
C9 a_n1629_n161# 0 1.70192f
C10 a_n3287_n161# 0 1.70192f
C11 a_n4945_n161# 0 1.7153f
C12 w_n5203_n362# 0 28.7441f
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_5H9LZ4 a_n100_n344# a_n158_118# a_n100_21# a_100_n612#
+ a_100_483# a_n100_n709# a_100_n247# 0 a_n158_n612# a_n100_386# a_n158_n247# a_100_118#
+ w_n358_n909# a_n158_483#
X0 a_100_118# a_n100_21# a_n158_118# w_n358_n909# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X1 a_100_483# a_n100_386# a_n158_483# w_n358_n909# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X2 a_100_n247# a_n100_n344# a_n158_n247# w_n358_n909# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X3 a_100_n612# a_n100_n709# a_n158_n612# w_n358_n909# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
C0 a_n100_n709# w_n358_n909# 0.256541f
C1 a_n100_21# a_n100_386# 0.138722f
C2 w_n358_n909# a_n100_386# 0.222637f
C3 a_n100_n344# a_n100_n709# 0.138722f
C4 a_n100_21# w_n358_n909# 0.176907f
C5 a_n100_21# a_n100_n344# 0.138722f
C6 a_n100_n344# w_n358_n909# 0.176907f
C7 a_n100_n709# 0 0.200574f
C8 a_n100_n344# 0 0.168079f
C9 a_n100_21# 0 0.168079f
C10 a_n100_386# 0 0.201694f
C11 w_n358_n909# 0 5.07037f
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_GG9S2Z a_n100_199# a_100_n487# a_100_581# a_100_n131#
+ a_n158_n487# a_n100_n157# a_n100_555# a_100_n843# a_n158_n131# a_n158_225# a_n100_n869#
+ a_n158_581# a_n158_n843# a_n100_n513# a_n292_n1003# a_100_225#
X0 a_100_n131# a_n100_n157# a_n158_n131# a_n292_n1003# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X1 a_100_581# a_n100_555# a_n158_581# a_n292_n1003# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X2 a_100_n843# a_n100_n869# a_n158_n843# a_n292_n1003# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X3 a_100_225# a_n100_199# a_n158_225# a_n292_n1003# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X4 a_100_n487# a_n100_n513# a_n158_n487# a_n292_n1003# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
C0 a_n100_n157# a_n100_199# 0.139254f
C1 a_n100_n869# a_n100_n513# 0.139254f
C2 a_n100_555# a_n100_199# 0.139254f
C3 a_n100_n157# a_n100_n513# 0.139254f
C4 a_100_n843# a_n292_n1003# 0.12711f
C5 a_n158_n843# a_n292_n1003# 0.12711f
C6 a_n100_n869# a_n292_n1003# 0.414462f
C7 a_100_n487# a_n292_n1003# 0.113612f
C8 a_n158_n487# a_n292_n1003# 0.113612f
C9 a_n100_n513# a_n292_n1003# 0.33438f
C10 a_100_n131# a_n292_n1003# 0.113612f
C11 a_n158_n131# a_n292_n1003# 0.113612f
C12 a_n100_n157# a_n292_n1003# 0.33438f
C13 a_100_225# a_n292_n1003# 0.113612f
C14 a_n158_225# a_n292_n1003# 0.113612f
C15 a_n100_199# a_n292_n1003# 0.33438f
C16 a_100_581# a_n292_n1003# 0.125529f
C17 a_n158_581# a_n292_n1003# 0.125529f
C18 a_n100_555# a_n292_n1003# 0.4464f
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_5HVT2F a_1629_n430# a_4945_n65# a_n3287_n1257#
+ a_n3287_n892# a_3345_n162# a_4945_665# a_n3287_568# w_n5203_n1457# a_3345_n1257#
+ a_3287_1030# a_n1629_933# a_n5003_1030# a_3287_n1160# a_n29_n795# a_n4945_n527#
+ a_n1687_1030# a_3345_933# a_n4945_933# a_1687_n1257# a_4945_n430# a_1687_n527# a_n1629_568#
+ a_29_933# a_29_n527# a_3345_568# a_n4945_568# a_n5003_n1160# a_3345_n892# a_n3345_300#
+ a_n3345_n1160# a_n3345_n795# a_n1687_n65# a_n1629_n162# a_29_568# a_29_n1257# a_1629_n795#
+ a_n3287_n527# a_3287_300# a_n29_300# a_n1687_665# a_n29_1030# a_n1687_n1160# a_3287_n430#
+ a_n5003_n430# a_n1687_n430# a_n4945_n162# a_4945_n795# a_1687_n162# a_1629_300#
+ a_n5003_300# a_n1629_n892# a_1687_203# a_4945_300# a_n3287_203# a_1629_1030# a_n3345_1030#
+ a_3345_n527# a_n3345_n65# a_29_n162# a_n3345_665# 0 a_n4945_n1257# a_n4945_n892#
+ a_n29_n430# a_3287_n65# a_n29_n65# a_n29_665# a_n3287_n162# a_3287_665# a_4945_n1160#
+ a_3287_n795# a_n5003_n795# a_1687_n892# a_n1629_203# a_4945_1030# a_n1629_n1257#
+ a_1687_933# a_n1687_n795# a_3345_203# a_n4945_203# a_n3287_933# a_n29_n1160# a_29_n892#
+ a_1629_n1160# a_n1629_n527# a_1629_n65# a_n5003_n65# a_1629_665# a_n5003_665# a_n3345_n430#
+ a_n1687_300# a_29_203# a_1687_568#
X0 a_n29_665# a_n1629_568# a_n1687_665# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1 a_n3345_n795# a_n4945_n892# a_n5003_n795# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=8
X2 a_n29_300# a_n1629_203# a_n1687_300# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X3 a_4945_n430# a_3345_n527# a_3287_n430# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=8
X4 a_3287_n795# a_1687_n892# a_1629_n795# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X5 a_n29_1030# a_n1629_933# a_n1687_1030# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X6 a_n1687_n795# a_n3287_n892# a_n3345_n795# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X7 a_n3345_665# a_n4945_568# a_n5003_665# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=8
X8 a_n3345_300# a_n4945_203# a_n5003_300# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=8
X9 a_n1687_n65# a_n3287_n162# a_n3345_n65# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X10 a_n29_n1160# a_n1629_n1257# a_n1687_n1160# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X11 a_1629_665# a_29_568# a_n29_665# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X12 a_4945_n795# a_3345_n892# a_3287_n795# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=8
X13 a_n29_n430# a_n1629_n527# a_n1687_n430# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X14 a_3287_665# a_1687_568# a_1629_665# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X15 a_1629_1030# a_29_933# a_n29_1030# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X16 a_1629_300# a_29_203# a_n29_300# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X17 a_4945_665# a_3345_568# a_3287_665# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=8
X18 a_3287_300# a_1687_203# a_1629_300# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X19 a_n29_n65# a_n1629_n162# a_n1687_n65# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X20 a_n3345_1030# a_n4945_933# a_n5003_1030# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=8
X21 a_4945_300# a_3345_203# a_3287_300# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=8
X22 a_3287_1030# a_1687_933# a_1629_1030# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X23 a_n3345_n65# a_n4945_n162# a_n5003_n65# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=8
X24 a_n1687_1030# a_n3287_933# a_n3345_1030# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X25 a_n29_n795# a_n1629_n892# a_n1687_n795# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X26 a_n3345_n1160# a_n4945_n1257# a_n5003_n1160# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=8
X27 a_1629_n430# a_29_n527# a_n29_n430# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X28 a_n1687_n1160# a_n3287_n1257# a_n3345_n1160# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X29 a_4945_n1160# a_3345_n1257# a_3287_n1160# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=8
X30 a_1629_n65# a_29_n162# a_n29_n65# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X31 a_n3345_n430# a_n4945_n527# a_n5003_n430# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=8
X32 a_4945_1030# a_3345_933# a_3287_1030# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=8
X33 a_n1687_665# a_n3287_568# a_n3345_665# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X34 a_3287_n65# a_1687_n162# a_1629_n65# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X35 a_3287_n430# a_1687_n527# a_1629_n430# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X36 a_1629_n1160# a_29_n1257# a_n29_n1160# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X37 a_n1687_n430# a_n3287_n527# a_n3345_n430# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X38 a_n1687_300# a_n3287_203# a_n3345_300# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X39 a_4945_n65# a_3345_n162# a_3287_n65# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=8
X40 a_1629_n795# a_29_n892# a_n29_n795# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X41 a_3287_n1160# a_1687_n1257# a_1629_n1160# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
C0 a_n1629_n892# a_n1629_n1257# 1.09385f
C1 w_n5203_n1457# a_3345_203# 0.847746f
C2 w_n5203_n1457# a_n3287_568# 0.823093f
C3 w_n5203_n1457# a_n4945_n527# 0.847746f
C4 a_n1629_n892# a_n1629_n527# 1.09385f
C5 a_n3287_203# a_n3287_n162# 1.09385f
C6 a_n4945_n527# a_n4945_n162# 1.09385f
C7 a_3345_203# a_3345_n162# 1.09385f
C8 a_1687_568# a_1687_933# 1.09385f
C9 w_n5203_n1457# a_n4945_n162# 0.847746f
C10 w_n5203_n1457# a_3345_n162# 0.847746f
C11 a_3345_n527# w_n5203_n1457# 0.847746f
C12 w_n5203_n1457# a_n1629_933# 1.18871f
C13 a_1687_n892# w_n5203_n1457# 0.823093f
C14 a_n4945_568# a_n4945_933# 1.09385f
C15 a_29_n527# w_n5203_n1457# 0.823093f
C16 a_3345_n527# a_3345_n162# 1.09385f
C17 a_1687_n162# a_1687_203# 1.09385f
C18 a_n3287_n892# a_n3287_n527# 1.09385f
C19 w_n5203_n1457# a_3345_n1257# 1.4835f
C20 a_29_n1257# a_29_n892# 1.09385f
C21 w_n5203_n1457# a_n4945_933# 1.21336f
C22 w_n5203_n1457# a_1687_n162# 0.823093f
C23 a_n4945_203# a_n4945_568# 1.09385f
C24 a_29_203# a_29_n162# 1.09385f
C25 w_n5203_n1457# a_n1629_n162# 0.823093f
C26 a_1687_203# a_1687_568# 1.09385f
C27 a_n1629_568# a_n1629_203# 1.09385f
C28 a_3345_203# a_3345_568# 1.09385f
C29 w_n5203_n1457# a_n3287_n162# 0.823093f
C30 w_n5203_n1457# a_3345_568# 0.847746f
C31 w_n5203_n1457# a_n4945_203# 0.847746f
C32 a_n4945_n527# a_n4945_n892# 1.09385f
C33 w_n5203_n1457# a_n1629_n1257# 1.45885f
C34 w_n5203_n1457# a_1687_568# 0.823093f
C35 a_29_203# a_29_568# 1.09385f
C36 a_n4945_203# a_n4945_n162# 1.09385f
C37 w_n5203_n1457# a_n3287_n527# 0.823093f
C38 w_n5203_n1457# a_n4945_n892# 0.847746f
C39 w_n5203_n1457# a_1687_n527# 0.823093f
C40 w_n5203_n1457# a_3345_n892# 0.847746f
C41 w_n5203_n1457# a_3345_933# 1.21336f
C42 w_n5203_n1457# a_1687_n1257# 1.45885f
C43 w_n5203_n1457# a_n4945_n1257# 1.4835f
C44 w_n5203_n1457# a_n1629_n527# 0.823093f
C45 a_3345_n527# a_3345_n892# 1.09385f
C46 w_n5203_n1457# a_n1629_n892# 0.823093f
C47 a_1687_n892# a_1687_n527# 1.09385f
C48 a_1687_n892# a_1687_n1257# 1.09385f
C49 a_29_933# a_29_568# 1.09385f
C50 a_n3287_568# a_n3287_203# 1.09385f
C51 a_3345_n1257# a_3345_n892# 1.09385f
C52 w_n5203_n1457# a_n1629_203# 0.823093f
C53 a_n3287_n1257# a_n3287_n892# 1.09385f
C54 w_n5203_n1457# a_29_n892# 0.823093f
C55 w_n5203_n1457# a_29_n1257# 1.45885f
C56 w_n5203_n1457# a_n3287_203# 0.823093f
C57 w_n5203_n1457# a_29_203# 0.823093f
C58 w_n5203_n1457# a_1687_933# 1.18871f
C59 w_n5203_n1457# a_29_n162# 0.823093f
C60 a_1687_n162# a_1687_n527# 1.09385f
C61 a_29_n527# a_29_n892# 1.09385f
C62 a_n3287_568# a_n3287_933# 1.09385f
C63 w_n5203_n1457# a_n3287_n892# 0.823093f
C64 w_n5203_n1457# a_n1629_568# 0.823093f
C65 w_n5203_n1457# a_29_933# 1.18871f
C66 a_n1629_n162# a_n1629_n527# 1.09385f
C67 w_n5203_n1457# a_n3287_933# 1.18871f
C68 a_29_n527# a_29_n162# 1.09385f
C69 a_n3287_n162# a_n3287_n527# 1.09385f
C70 w_n5203_n1457# a_29_568# 0.823093f
C71 a_n1629_933# a_n1629_568# 1.09385f
C72 a_3345_568# a_3345_933# 1.09385f
C73 a_n1629_n162# a_n1629_203# 1.09385f
C74 a_n3287_n1257# w_n5203_n1457# 1.45885f
C75 w_n5203_n1457# a_n4945_568# 0.847746f
C76 w_n5203_n1457# a_1687_203# 0.823093f
C77 a_n4945_n1257# a_n4945_n892# 1.09385f
C78 a_3345_n1257# 0 1.4406f
C79 a_1687_n1257# 0 1.42722f
C80 a_29_n1257# 0 1.42722f
C81 a_n1629_n1257# 0 1.42722f
C82 a_n3287_n1257# 0 1.42722f
C83 a_n4945_n1257# 0 1.4406f
C84 a_3345_n892# 0 1.18572f
C85 a_1687_n892# 0 1.17234f
C86 a_29_n892# 0 1.17234f
C87 a_n1629_n892# 0 1.17234f
C88 a_n3287_n892# 0 1.17234f
C89 a_n4945_n892# 0 1.18572f
C90 a_3345_n527# 0 1.18572f
C91 a_1687_n527# 0 1.17234f
C92 a_29_n527# 0 1.17234f
C93 a_n1629_n527# 0 1.17234f
C94 a_n3287_n527# 0 1.17234f
C95 a_n4945_n527# 0 1.18572f
C96 a_3345_n162# 0 1.18572f
C97 a_1687_n162# 0 1.17234f
C98 a_29_n162# 0 1.17234f
C99 a_n1629_n162# 0 1.17234f
C100 a_n3287_n162# 0 1.17234f
C101 a_n4945_n162# 0 1.18572f
C102 a_3345_203# 0 1.18572f
C103 a_1687_203# 0 1.17234f
C104 a_29_203# 0 1.17234f
C105 a_n1629_203# 0 1.17234f
C106 a_n3287_203# 0 1.17234f
C107 a_n4945_203# 0 1.18572f
C108 a_3345_568# 0 1.18572f
C109 a_1687_568# 0 1.17234f
C110 a_29_568# 0 1.17234f
C111 a_n1629_568# 0 1.17234f
C112 a_n3287_568# 0 1.17234f
C113 a_n4945_568# 0 1.18572f
C114 a_3345_933# 0 1.46042f
C115 a_1687_933# 0 1.44704f
C116 a_29_933# 0 1.44704f
C117 a_n1629_933# 0 1.44704f
C118 a_n3287_933# 0 1.44704f
C119 a_n4945_933# 0 1.46042f
C120 w_n5203_n1457# 0 98.4735f
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_HZHY2Z a_861_n131# a_207_n157# a_n861_n157# a_n563_n131#
+ a_683_n131# a_n919_n131# a_29_n157# a_n683_n157# a_n385_n131# a_n1053_n291# a_741_n157#
+ a_505_n131# a_n505_n157# a_563_n157# a_n207_n131# a_327_n131# a_n327_n157# a_385_n157#
+ a_n29_n131# a_149_n131# a_n741_n131# a_n149_n157#
X0 a_n563_n131# a_n683_n157# a_n741_n131# a_n1053_n291# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X1 a_505_n131# a_385_n157# a_327_n131# a_n1053_n291# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X2 a_n385_n131# a_n505_n157# a_n563_n131# a_n1053_n291# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X3 a_327_n131# a_207_n157# a_149_n131# a_n1053_n291# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X4 a_149_n131# a_29_n157# a_n29_n131# a_n1053_n291# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X5 a_861_n131# a_741_n157# a_683_n131# a_n1053_n291# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.6
X6 a_n207_n131# a_n327_n157# a_n385_n131# a_n1053_n291# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X7 a_n741_n131# a_n861_n157# a_n919_n131# a_n1053_n291# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.6
X8 a_683_n131# a_563_n157# a_505_n131# a_n1053_n291# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X9 a_n29_n131# a_n149_n157# a_n207_n131# a_n1053_n291# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
C0 a_861_n131# a_n1053_n291# 0.135212f
C1 a_n919_n131# a_n1053_n291# 0.135212f
C2 a_741_n157# a_n1053_n291# 0.316895f
C3 a_563_n157# a_n1053_n291# 0.280633f
C4 a_385_n157# a_n1053_n291# 0.280633f
C5 a_207_n157# a_n1053_n291# 0.280633f
C6 a_29_n157# a_n1053_n291# 0.280633f
C7 a_n149_n157# a_n1053_n291# 0.280633f
C8 a_n327_n157# a_n1053_n291# 0.280633f
C9 a_n505_n157# a_n1053_n291# 0.280633f
C10 a_n683_n157# a_n1053_n291# 0.280633f
C11 a_n861_n157# a_n1053_n291# 0.316895f
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_ZV8547 a_3345_439# a_3287_527# a_1687_21# a_n4945_439#
+ a_n5003_n1563# a_1629_n1145# a_3345_n815# a_3287_n727# a_29_439# a_n5003_n727# a_n3345_n1563#
+ a_n4945_1275# a_n29_1363# a_4945_n309# a_3345_n397# a_n1687_n727# a_1687_1275# a_n1687_n1563#
+ a_n5003_527# a_1629_527# a_n4945_n1651# a_29_n1233# a_3287_n1145# a_n3345_109# a_29_1275#
+ a_4945_527# a_n1687_945# a_n3287_21# a_n29_109# a_3287_109# a_n3345_1363# a_29_21#
+ a_n5003_n1145# a_n1629_n1651# a_n1629_n815# a_1629_1363# a_n3287_1275# a_1687_857#
+ a_3287_n309# a_n29_n727# a_n5003_n309# a_n3345_n1145# a_n3287_857# a_n1629_n397#
+ a_n1687_n309# a_n1687_n1145# a_n5003_109# a_1629_109# a_n4945_n815# a_n4945_n1233#
+ a_n3287_n1651# a_4945_1363# a_n4945_21# a_4945_n1563# a_n3345_945# a_1687_n815#
+ a_3345_n1651# a_n1629_21# a_4945_109# a_n1687_527# a_n4945_n397# a_n3345_n727# a_n1629_857#
+ a_3345_1275# a_n29_n1563# a_1629_n727# a_1687_n1651# a_29_n815# a_n29_945# a_n1629_n1233#
+ a_1687_n397# a_3345_857# a_3287_945# a_n4945_857# a_3345_21# a_1629_n1563# a_1687_439#
+ a_n29_n309# a_29_n397# a_29_857# a_n3287_439# a_n3287_n815# a_3287_1363# a_n5003_1363#
+ a_4945_n727# a_n5137_n1785# a_n3287_n1233# a_n1687_1363# a_n5003_945# a_1629_945#
+ a_4945_n1145# a_29_n1651# a_3287_n1563# a_n3345_527# a_n3287_n397# a_3345_n1233#
+ a_4945_945# a_n1687_109# a_n1629_1275# a_n3345_n309# a_n1629_439# a_n29_n1145# a_1629_n309#
+ a_1687_n1233# a_n29_527#
X0 a_n1687_527# a_n3287_439# a_n3345_527# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1 a_3287_n1563# a_1687_n1651# a_1629_n1563# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X2 a_3287_945# a_1687_857# a_1629_945# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X3 a_1629_109# a_29_21# a_n29_109# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X4 a_4945_945# a_3345_857# a_3287_945# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=8
X5 a_3287_109# a_1687_21# a_1629_109# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X6 a_4945_n727# a_3345_n815# a_3287_n727# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=8
X7 a_4945_109# a_3345_21# a_3287_109# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=8
X8 a_n29_527# a_n1629_439# a_n1687_527# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X9 a_n3345_n1145# a_n4945_n1233# a_n5003_n1145# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=8
X10 a_n29_1363# a_n1629_1275# a_n1687_1363# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X11 a_1629_n309# a_29_n397# a_n29_n309# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X12 a_n1687_n1145# a_n3287_n1233# a_n3345_n1145# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X13 a_n3345_527# a_n4945_439# a_n5003_527# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=8
X14 a_4945_n1145# a_3345_n1233# a_3287_n1145# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=8
X15 a_n29_n1563# a_n1629_n1651# a_n1687_n1563# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X16 a_n3345_n309# a_n4945_n397# a_n5003_n309# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=8
X17 a_3287_n309# a_1687_n397# a_1629_n309# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X18 a_n29_n727# a_n1629_n815# a_n1687_n727# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X19 a_1629_n1145# a_29_n1233# a_n29_n1145# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X20 a_n1687_n309# a_n3287_n397# a_n3345_n309# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X21 a_n1687_945# a_n3287_857# a_n3345_945# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X22 a_1629_527# a_29_439# a_n29_527# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X23 a_n1687_109# a_n3287_21# a_n3345_109# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X24 a_3287_n1145# a_1687_n1233# a_1629_n1145# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X25 a_1629_1363# a_29_1275# a_n29_1363# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X26 a_3287_527# a_1687_439# a_1629_527# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X27 a_4945_527# a_3345_439# a_3287_527# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=8
X28 a_4945_n309# a_3345_n397# a_3287_n309# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=8
X29 a_n3345_1363# a_n4945_1275# a_n5003_1363# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=8
X30 a_n29_945# a_n1629_857# a_n1687_945# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X31 a_3287_1363# a_1687_1275# a_1629_1363# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X32 a_n29_109# a_n1629_21# a_n1687_109# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X33 a_n3345_n1563# a_n4945_n1651# a_n5003_n1563# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=8
X34 a_n1687_1363# a_n3287_1275# a_n3345_1363# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X35 a_1629_n727# a_29_n815# a_n29_n727# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X36 a_n1687_n1563# a_n3287_n1651# a_n3345_n1563# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X37 a_4945_n1563# a_3345_n1651# a_3287_n1563# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=8
X38 a_n3345_945# a_n4945_857# a_n5003_945# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=8
X39 a_n3345_n727# a_n4945_n815# a_n5003_n727# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=8
X40 a_n3345_109# a_n4945_21# a_n5003_109# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=8
X41 a_3287_n727# a_1687_n815# a_1629_n727# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X42 a_n29_n1145# a_n1629_n1233# a_n1687_n1145# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X43 a_1629_n1563# a_29_n1651# a_n29_n1563# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X44 a_n1687_n727# a_n3287_n815# a_n3345_n727# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X45 a_n29_n309# a_n1629_n397# a_n1687_n309# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X46 a_4945_1363# a_3345_1275# a_3287_1363# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=8
X47 a_1629_945# a_29_857# a_n29_945# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
C0 a_3345_n397# a_1687_n397# 0.104496f
C1 a_1687_857# a_1687_439# 1.65624f
C2 a_n1629_n815# a_n3287_n815# 0.104496f
C3 a_29_n1651# a_29_n1233# 1.65624f
C4 a_n3287_857# a_n1629_857# 0.104496f
C5 a_29_n397# a_1687_n397# 0.104496f
C6 a_3345_n397# a_3345_n815# 1.65624f
C7 a_n3287_857# a_n3287_1275# 1.65624f
C8 a_29_1275# a_29_857# 1.65624f
C9 a_n3287_n397# a_n3287_n815# 1.65624f
C10 a_3345_n1233# a_1687_n1233# 0.104496f
C11 a_3345_857# a_3345_439# 1.65624f
C12 a_29_n397# a_29_21# 1.65624f
C13 a_n1629_857# a_29_857# 0.104496f
C14 a_n1629_439# a_n1629_857# 1.65624f
C15 a_n1629_1275# a_29_1275# 0.104496f
C16 a_1687_n1233# a_1687_n1651# 1.65624f
C17 a_n4945_857# a_n4945_1275# 1.65624f
C18 a_n1629_n1651# a_n1629_n1233# 1.65624f
C19 a_n1629_21# a_29_21# 0.104496f
C20 a_1687_21# a_3345_21# 0.104496f
C21 a_n1629_1275# a_n1629_857# 1.65624f
C22 a_3345_439# a_1687_439# 0.104496f
C23 a_n1629_1275# a_n3287_1275# 0.104496f
C24 a_n3287_n1233# a_n4945_n1233# 0.104496f
C25 a_29_n1233# a_1687_n1233# 0.104496f
C26 a_n4945_21# a_n3287_21# 0.104496f
C27 a_n3287_n815# a_n3287_n1233# 1.65624f
C28 a_29_n1233# a_n1629_n1233# 0.104496f
C29 a_1687_1275# a_1687_857# 1.65624f
C30 a_n1629_n815# a_n1629_n397# 1.65624f
C31 a_n4945_21# a_n4945_439# 1.65624f
C32 a_3345_n1233# a_3345_n815# 1.65624f
C33 a_29_439# a_29_857# 1.65624f
C34 a_29_439# a_n1629_439# 0.104496f
C35 a_n3287_n397# a_n3287_21# 1.65624f
C36 a_n4945_n815# a_n4945_n397# 1.65624f
C37 a_n3287_n397# a_n1629_n397# 0.104496f
C38 a_29_n815# a_29_n1233# 1.65624f
C39 a_n3287_n1651# a_n3287_n1233# 1.65624f
C40 a_1687_n1233# a_1687_n815# 1.65624f
C41 a_n1629_n815# a_n1629_n1233# 1.65624f
C42 a_n4945_1275# a_n3287_1275# 0.104496f
C43 a_3345_1275# a_1687_1275# 0.104496f
C44 a_29_n815# a_1687_n815# 0.104496f
C45 a_3345_n397# a_3345_21# 1.65624f
C46 a_n4945_439# a_n4945_857# 1.65624f
C47 a_n1629_n815# a_29_n815# 0.104496f
C48 a_29_n397# a_n1629_n397# 0.104496f
C49 a_n4945_21# a_n4945_n397# 1.65624f
C50 a_n3287_439# a_n3287_21# 1.65624f
C51 a_1687_21# a_1687_n397# 1.65624f
C52 a_n3287_n397# a_n4945_n397# 0.104496f
C53 a_29_857# a_1687_857# 0.104496f
C54 a_n3287_439# a_n4945_439# 0.104496f
C55 a_29_439# a_29_21# 1.65624f
C56 a_n4945_857# a_n3287_857# 0.104496f
C57 a_n1629_21# a_n3287_21# 0.104496f
C58 a_29_439# a_1687_439# 0.104496f
C59 a_29_1275# a_1687_1275# 0.104496f
C60 a_1687_21# a_29_21# 0.104496f
C61 a_n1629_21# a_n1629_n397# 1.65624f
C62 a_3345_439# a_3345_21# 1.65624f
C63 a_3345_n1651# a_3345_n1233# 1.65624f
C64 a_1687_n397# a_1687_n815# 1.65624f
C65 a_n4945_n1651# a_n4945_n1233# 1.65624f
C66 a_n3287_439# a_n3287_857# 1.65624f
C67 a_1687_21# a_1687_439# 1.65624f
C68 a_n1629_n1651# a_n3287_n1651# 0.104496f
C69 a_n4945_n815# a_n4945_n1233# 1.65624f
C70 a_3345_857# a_1687_857# 0.104496f
C71 a_3345_n815# a_1687_n815# 0.104496f
C72 a_n4945_n815# a_n3287_n815# 0.104496f
C73 a_29_n397# a_29_n815# 1.65624f
C74 a_29_n1651# a_n1629_n1651# 0.104496f
C75 a_29_n1651# a_1687_n1651# 0.104496f
C76 a_n1629_n1233# a_n3287_n1233# 0.104496f
C77 a_n3287_439# a_n1629_439# 0.104496f
C78 a_3345_n1651# a_1687_n1651# 0.104496f
C79 a_n3287_n1651# a_n4945_n1651# 0.104496f
C80 a_3345_857# a_3345_1275# 1.65624f
C81 a_n1629_21# a_n1629_439# 1.65624f
C82 a_4945_n1563# a_n5137_n1785# 0.157617f
C83 a_3287_n1563# a_n5137_n1785# 0.107833f
C84 a_1629_n1563# a_n5137_n1785# 0.107833f
C85 a_n29_n1563# a_n5137_n1785# 0.107833f
C86 a_n1687_n1563# a_n5137_n1785# 0.107833f
C87 a_n3345_n1563# a_n5137_n1785# 0.107833f
C88 a_n5003_n1563# a_n5137_n1785# 0.157617f
C89 a_3345_n1651# a_n5137_n1785# 3.34043f
C90 a_1687_n1651# a_n5137_n1785# 3.27762f
C91 a_29_n1651# a_n5137_n1785# 3.27762f
C92 a_n1629_n1651# a_n5137_n1785# 3.27762f
C93 a_n3287_n1651# a_n5137_n1785# 3.27762f
C94 a_n4945_n1651# a_n5137_n1785# 3.34043f
C95 a_4945_n1145# a_n5137_n1785# 0.147177f
C96 a_n5003_n1145# a_n5137_n1785# 0.147177f
C97 a_3345_n1233# a_n5137_n1785# 2.34788f
C98 a_1687_n1233# a_n5137_n1785# 2.28507f
C99 a_29_n1233# a_n5137_n1785# 2.28507f
C100 a_n1629_n1233# a_n5137_n1785# 2.28507f
C101 a_n3287_n1233# a_n5137_n1785# 2.28507f
C102 a_n4945_n1233# a_n5137_n1785# 2.34788f
C103 a_4945_n727# a_n5137_n1785# 0.147177f
C104 a_n5003_n727# a_n5137_n1785# 0.147177f
C105 a_3345_n815# a_n5137_n1785# 2.34788f
C106 a_1687_n815# a_n5137_n1785# 2.28507f
C107 a_29_n815# a_n5137_n1785# 2.28507f
C108 a_n1629_n815# a_n5137_n1785# 2.28507f
C109 a_n3287_n815# a_n5137_n1785# 2.28507f
C110 a_n4945_n815# a_n5137_n1785# 2.34788f
C111 a_4945_n309# a_n5137_n1785# 0.147177f
C112 a_n5003_n309# a_n5137_n1785# 0.147177f
C113 a_3345_n397# a_n5137_n1785# 2.34788f
C114 a_1687_n397# a_n5137_n1785# 2.28507f
C115 a_29_n397# a_n5137_n1785# 2.28507f
C116 a_n1629_n397# a_n5137_n1785# 2.28507f
C117 a_n3287_n397# a_n5137_n1785# 2.28507f
C118 a_n4945_n397# a_n5137_n1785# 2.34788f
C119 a_4945_109# a_n5137_n1785# 0.147177f
C120 a_n5003_109# a_n5137_n1785# 0.147177f
C121 a_3345_21# a_n5137_n1785# 2.34788f
C122 a_1687_21# a_n5137_n1785# 2.28507f
C123 a_29_21# a_n5137_n1785# 2.28507f
C124 a_n1629_21# a_n5137_n1785# 2.28507f
C125 a_n3287_21# a_n5137_n1785# 2.28507f
C126 a_n4945_21# a_n5137_n1785# 2.34788f
C127 a_4945_527# a_n5137_n1785# 0.147177f
C128 a_n5003_527# a_n5137_n1785# 0.147177f
C129 a_3345_439# a_n5137_n1785# 2.34788f
C130 a_1687_439# a_n5137_n1785# 2.28507f
C131 a_29_439# a_n5137_n1785# 2.28507f
C132 a_n1629_439# a_n5137_n1785# 2.28507f
C133 a_n3287_439# a_n5137_n1785# 2.28507f
C134 a_n4945_439# a_n5137_n1785# 2.34788f
C135 a_4945_945# a_n5137_n1785# 0.147177f
C136 a_n5003_945# a_n5137_n1785# 0.147177f
C137 a_3345_857# a_n5137_n1785# 2.34788f
C138 a_1687_857# a_n5137_n1785# 2.28507f
C139 a_29_857# a_n5137_n1785# 2.28507f
C140 a_n1629_857# a_n5137_n1785# 2.28507f
C141 a_n3287_857# a_n5137_n1785# 2.28507f
C142 a_n4945_857# a_n5137_n1785# 2.34788f
C143 a_4945_1363# a_n5137_n1785# 0.157617f
C144 a_3287_1363# a_n5137_n1785# 0.107833f
C145 a_1629_1363# a_n5137_n1785# 0.107833f
C146 a_n29_1363# a_n5137_n1785# 0.107833f
C147 a_n1687_1363# a_n5137_n1785# 0.107833f
C148 a_n3345_1363# a_n5137_n1785# 0.107833f
C149 a_n5003_1363# a_n5137_n1785# 0.157617f
C150 a_3345_1275# a_n5137_n1785# 3.34043f
C151 a_1687_1275# a_n5137_n1785# 3.27762f
C152 a_29_1275# a_n5137_n1785# 3.27762f
C153 a_n1629_1275# a_n5137_n1785# 3.27762f
C154 a_n3287_1275# a_n5137_n1785# 3.27762f
C155 a_n4945_1275# a_n5137_n1785# 3.34043f
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_5HV9F5 a_1629_118# a_n5003_118# a_1687_21# a_n29_n612#
+ a_n3287_n344# a_4945_118# a_29_386# a_n1687_483# a_n29_n247# a_n3345_n612# a_n1629_n709#
+ a_1629_n612# a_3345_n344# a_29_21# a_n3287_21# a_n3345_n247# a_n3345_483# w_n5203_n909#
+ a_n4945_n709# a_1629_n247# a_4945_n612# a_n1687_118# a_1687_n709# a_3287_483# a_n29_483#
+ a_29_n709# a_n4945_21# a_n1629_21# a_4945_n247# a_n1629_n344# a_n3287_n709# a_1629_483#
+ a_n5003_483# 0 a_3345_21# a_1687_386# a_3287_n612# a_n5003_n612# a_n3345_118# a_4945_483#
+ a_n3287_386# a_n1687_n612# a_n4945_n344# a_n29_118# a_3287_n247# a_n5003_n247# a_1687_n344#
+ a_3287_118# a_n1687_n247# a_n1629_386# a_3345_n709# a_29_n344# a_3345_386# a_n4945_386#
X0 a_4945_n247# a_3345_n344# a_3287_n247# w_n5203_n909# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=8
X1 a_4945_n612# a_3345_n709# a_3287_n612# w_n5203_n909# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=8
X2 a_n29_118# a_n1629_21# a_n1687_118# w_n5203_n909# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X3 a_n1687_483# a_n3287_386# a_n3345_483# w_n5203_n909# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X4 a_n3345_118# a_n4945_21# a_n5003_118# w_n5203_n909# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=8
X5 a_n29_483# a_n1629_386# a_n1687_483# w_n5203_n909# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X6 a_n29_n612# a_n1629_n709# a_n1687_n612# w_n5203_n909# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X7 a_n29_n247# a_n1629_n344# a_n1687_n247# w_n5203_n909# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X8 a_1629_118# a_29_21# a_n29_118# w_n5203_n909# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X9 a_n3345_483# a_n4945_386# a_n5003_483# w_n5203_n909# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=8
X10 a_3287_118# a_1687_21# a_1629_118# w_n5203_n909# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X11 a_4945_118# a_3345_21# a_3287_118# w_n5203_n909# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=8
X12 a_1629_483# a_29_386# a_n29_483# w_n5203_n909# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X13 a_1629_n247# a_29_n344# a_n29_n247# w_n5203_n909# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X14 a_1629_n612# a_29_n709# a_n29_n612# w_n5203_n909# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X15 a_3287_483# a_1687_386# a_1629_483# w_n5203_n909# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X16 a_n3345_n247# a_n4945_n344# a_n5003_n247# w_n5203_n909# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=8
X17 a_n3345_n612# a_n4945_n709# a_n5003_n612# w_n5203_n909# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=8
X18 a_4945_483# a_3345_386# a_3287_483# w_n5203_n909# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=8
X19 a_3287_n612# a_1687_n709# a_1629_n612# w_n5203_n909# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X20 a_3287_n247# a_1687_n344# a_1629_n247# w_n5203_n909# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X21 a_n1687_n247# a_n3287_n344# a_n3345_n247# w_n5203_n909# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X22 a_n1687_n612# a_n3287_n709# a_n3345_n612# w_n5203_n909# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X23 a_n1687_118# a_n3287_21# a_n3345_118# w_n5203_n909# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
C0 a_n3287_386# w_n5203_n909# 1.18842f
C1 a_n1629_21# a_n1629_n344# 1.09385f
C2 a_n4945_21# a_n4945_386# 1.09385f
C3 a_n3287_n344# w_n5203_n909# 0.823093f
C4 a_n3287_21# w_n5203_n909# 0.823093f
C5 a_3345_n344# w_n5203_n909# 0.847746f
C6 a_1687_n709# w_n5203_n909# 1.45885f
C7 a_3345_21# a_3345_386# 1.09385f
C8 a_n3287_n344# a_n3287_n709# 1.09385f
C9 a_3345_n344# a_3345_21# 1.09385f
C10 a_n4945_n344# w_n5203_n909# 0.847746f
C11 a_1687_21# w_n5203_n909# 0.823093f
C12 w_n5203_n909# a_29_386# 1.18842f
C13 a_n1629_21# a_n1629_386# 1.09385f
C14 w_n5203_n909# a_n1629_n344# 0.823093f
C15 a_3345_n344# a_3345_n709# 1.09385f
C16 w_n5203_n909# a_29_n344# 0.823093f
C17 a_n1629_n709# w_n5203_n909# 1.45885f
C18 w_n5203_n909# a_3345_21# 0.847746f
C19 a_n3287_n709# w_n5203_n909# 1.45885f
C20 a_n4945_386# w_n5203_n909# 1.21308f
C21 a_n3287_21# a_n3287_386# 1.09385f
C22 a_1687_n344# a_1687_n709# 1.09385f
C23 a_n4945_21# a_n4945_n344# 1.09385f
C24 a_1687_21# a_1687_386# 1.09385f
C25 a_n1629_n709# a_n1629_n344# 1.09385f
C26 a_29_21# a_29_386# 1.09385f
C27 a_29_21# w_n5203_n909# 0.823093f
C28 a_1687_386# w_n5203_n909# 1.18842f
C29 a_n4945_21# w_n5203_n909# 0.847746f
C30 a_n3287_n344# a_n3287_21# 1.09385f
C31 w_n5203_n909# a_3345_n709# 1.4835f
C32 a_29_n709# w_n5203_n909# 1.45885f
C33 a_n4945_n344# a_n4945_n709# 1.09385f
C34 w_n5203_n909# a_n4945_n709# 1.4835f
C35 w_n5203_n909# a_n1629_386# 1.18842f
C36 a_1687_21# a_1687_n344# 1.09385f
C37 a_1687_n344# w_n5203_n909# 0.823093f
C38 a_n1629_21# w_n5203_n909# 0.823093f
C39 a_29_21# a_29_n344# 1.09385f
C40 w_n5203_n909# a_3345_386# 1.21308f
C41 a_29_n709# a_29_n344# 1.09385f
C42 a_3345_n709# 0 1.4406f
C43 a_1687_n709# 0 1.42722f
C44 a_29_n709# 0 1.42722f
C45 a_n1629_n709# 0 1.42722f
C46 a_n3287_n709# 0 1.42722f
C47 a_n4945_n709# 0 1.4406f
C48 a_3345_n344# 0 1.18572f
C49 a_1687_n344# 0 1.17234f
C50 a_29_n344# 0 1.17234f
C51 a_n1629_n344# 0 1.17234f
C52 a_n3287_n344# 0 1.17234f
C53 a_n4945_n344# 0 1.18572f
C54 a_3345_21# 0 1.18572f
C55 a_1687_21# 0 1.17234f
C56 a_29_21# 0 1.17234f
C57 a_n1629_21# 0 1.17234f
C58 a_n3287_21# 0 1.17234f
C59 a_n4945_21# 0 1.18572f
C60 a_3345_386# 0 1.46089f
C61 a_1687_386# 0 1.44751f
C62 a_29_386# 0 1.44751f
C63 a_n1629_386# 0 1.44751f
C64 a_n3287_386# 0 1.44751f
C65 a_n4945_386# 0 1.46089f
C66 w_n5203_n909# 0 63.574802f
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_W8MWAU a_n741_n136# w_n1119_n362# a_861_n136#
+ a_n327_n162# a_385_n162# a_n563_n136# a_683_n136# a_n149_n162# a_n919_n136# a_207_n162#
+ a_n385_n136# a_n861_n162# a_505_n136# a_29_n162# 0 a_n207_n136# a_n683_n162# a_741_n162#
+ a_327_n136# a_n505_n162# a_n29_n136# a_563_n162# a_149_n136#
X0 a_861_n136# a_741_n162# a_683_n136# w_n1119_n362# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.6
X1 a_n207_n136# a_n327_n162# a_n385_n136# w_n1119_n362# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X2 a_n741_n136# a_n861_n162# a_n919_n136# w_n1119_n362# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.6
X3 a_683_n136# a_563_n162# a_505_n136# w_n1119_n362# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X4 a_n29_n136# a_n149_n162# a_n207_n136# w_n1119_n362# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X5 a_n563_n136# a_n683_n162# a_n741_n136# w_n1119_n362# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X6 a_505_n136# a_385_n162# a_327_n136# w_n1119_n362# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X7 a_n385_n136# a_n505_n162# a_n563_n136# w_n1119_n362# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X8 a_327_n136# a_207_n162# a_149_n136# w_n1119_n362# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X9 a_149_n136# a_29_n162# a_n29_n136# w_n1119_n362# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
C0 a_n861_n162# w_n1119_n362# 0.187694f
C1 w_n1119_n362# a_385_n162# 0.163041f
C2 a_n327_n162# w_n1119_n362# 0.163041f
C3 w_n1119_n362# a_741_n162# 0.187694f
C4 a_n505_n162# w_n1119_n362# 0.163041f
C5 a_563_n162# w_n1119_n362# 0.163041f
C6 a_207_n162# w_n1119_n362# 0.163041f
C7 w_n1119_n362# a_29_n162# 0.163041f
C8 a_n683_n162# w_n1119_n362# 0.163041f
C9 w_n1119_n362# a_n149_n162# 0.163041f
C10 a_741_n162# 0 0.13534f
C11 a_563_n162# 0 0.121959f
C12 a_385_n162# 0 0.121959f
C13 a_207_n162# 0 0.121959f
C14 a_29_n162# 0 0.121959f
C15 a_n149_n162# 0 0.121959f
C16 a_n327_n162# 0 0.121959f
C17 a_n505_n162# 0 0.121959f
C18 a_n683_n162# 0 0.121959f
C19 a_n861_n162# 0 0.13534f
C20 w_n1119_n362# 0 6.30984f
.ends

.subckt comparator ibias out ena ena_b vt vinp n0 avss vpp vinn avdd vm vn vnn n1
Xsky130_fd_pr__nfet_g5v0d10v5_T82T27_1 n0 vm vm avss vn avss avss avss vm vm vn avss
+ avss vn vn avss avss vn vm avss avss avss avss avss avss vt avss sky130_fd_pr__nfet_g5v0d10v5_T82T27
Xsky130_fd_pr__pfet_g5v0d10v5_3HV7M9_0 avdd vm vnn avdd avdd vpp avdd vpp avss avdd
+ avdd vnn n0 avdd avdd sky130_fd_pr__pfet_g5v0d10v5_3HV7M9
Xsky130_fd_pr__pfet_g5v0d10v5_5H9LZ4_0 ena avdd ena vn vpp ena_b ena_b avss ibias
+ ena avdd vnn avdd avdd sky130_fd_pr__pfet_g5v0d10v5_5H9LZ4
Xsky130_fd_pr__nfet_g5v0d10v5_GG9S2Z_0 ena vm vn vn avss ena_b ena n0 avss avss ena_b
+ ibias avss ena_b avss ena_b sky130_fd_pr__nfet_g5v0d10v5_GG9S2Z
Xsky130_fd_pr__pfet_g5v0d10v5_5HVT2F_0 vnn avdd vnn vnn avdd avdd vnn avdd avdd avdd
+ vnn avdd avdd avdd avdd vpp avdd avdd vpp avdd vpp vnn vpp vpp avdd avdd avdd avdd
+ avdd avdd avdd vpp vnn vpp vpp vnn vnn avdd avdd vpp avdd vpp avdd avdd vpp avdd
+ avdd vpp vnn avdd vnn vpp avdd vnn vnn avdd avdd avdd vpp avdd avss avdd avdd avdd
+ avdd avdd avdd vnn avdd avdd avdd avdd vpp vnn avdd vnn vpp vpp avdd avdd vnn avdd
+ vpp vnn vnn vnn avdd vnn avdd avdd vpp vpp vpp sky130_fd_pr__pfet_g5v0d10v5_5HVT2F
Xsky130_fd_pr__nfet_g5v0d10v5_HZHY2Z_0 avss n1 n1 avss n1 avss n1 n1 out avss n0 avss
+ n1 n0 avss out n1 n1 out avss out n1 sky130_fd_pr__nfet_g5v0d10v5_HZHY2Z
Xsky130_fd_pr__nfet_g5v0d10v5_ZV8547_0 avss vnn vinn avss vt vt avss vnn vinp vt vnn
+ avss vpp vt avss vt vinn vt vt vt avss vinp vnn vnn vinp vt vt vinn vpp vnn vnn
+ vinp vt vinp vinp vt vinn vinn vnn vpp vt vnn vinn vinp vt vt vt vt avss avss vinn
+ vt avss vt vnn vinn avss vinp vt vt avss vnn vinp avss vpp vt vinn vinp vpp vinp
+ vinn avss vnn avss avss vt vinn vpp vinp vinp vinn vinn vnn vt vt vt vinn vt vt
+ vt vt vinp vnn vnn vinn avss vt vt vinp vnn vinp vpp vt vinn vpp sky130_fd_pr__nfet_g5v0d10v5_ZV8547
Xsky130_fd_pr__pfet_g5v0d10v5_5HV9F5_0 vnn avdd vnn avdd vpp avdd vnn vpp avdd avdd
+ vpp vnn avdd vnn vpp avdd avdd avdd avdd vnn avdd vpp vnn avdd avdd vnn avdd vpp
+ avdd vpp vpp vnn avdd avss avdd vnn avdd avdd avdd avdd vpp vpp avdd avdd avdd avdd
+ vnn avdd vpp vpp avdd vnn avdd avdd sky130_fd_pr__pfet_g5v0d10v5_5HV9F5
Xsky130_fd_pr__pfet_g5v0d10v5_W8MWAU_0 out avdd avdd n1 n1 avdd n1 n1 avdd n1 out
+ n1 avdd n1 avss avdd n1 n0 out n1 out n0 avdd sky130_fd_pr__pfet_g5v0d10v5_W8MWAU
C0 vt vn 0.111311f
C1 vinp vnn 0.779798f
C2 n0 vinp 0.529892f
C3 n0 vnn 0.42855f
C4 vn ibias 0.175171f
C5 avdd ena 0.684847f
C6 vpp vm 0.636921f
C7 vinn avss 0.480122f
C8 avdd vt 0.142054p
C9 ena_b ena 0.288446f
C10 vm avss 3.978539f
C11 vinp vt 22.104887f
C12 vt vnn 4.270693f
C13 n1 avss 0.866082f
C14 avdd vinn 0.485544f
C15 vm vn 0.237962f
C16 vinp vinn 2.328362f
C17 avdd vm 0.366792f
C18 vpp avss 1.048114f
C19 vinn vnn 2.30985f
C20 ena ibias 0.627137f
C21 avdd n1 1.032601f
C22 out n1 1.388767f
C23 vpp vn 0.332307f
C24 vnn vm 0.474767f
C25 n0 vm 2.502012f
C26 n0 n1 0.730567f
C27 avdd vpp 9.440008f
C28 vt vinn 23.074863f
C29 vn avss 2.95165f
C30 vinp vpp 2.164735f
C31 avdd avss 12.92849f
C32 vpp vnn 6.630513f
C33 n0 vpp 0.258129f
C34 out avss 0.926372f
C35 ena_b avss 0.713504f
C36 avdd vn 0.689774f
C37 vinp avss 0.729608f
C38 vnn avss 1.947571f
C39 n0 avss 2.854966f
C40 ena_b vn 1.03509f
C41 vinp vn 0.72801f
C42 vt vpp 2.57115f
C43 avdd out 2.006841f
C44 vnn vn 0.298893f
C45 n0 vn 1.991385f
C46 avdd ena_b 0.614152f
C47 avdd vinp 1.780272f
C48 ena avss 0.112348f
C49 avdd vnn 9.45953f
C50 n0 avdd 0.680561f
C51 vt avss 26.043423f
C52 n0 out 0.388405f
C53 vinn vpp 2.498551f
C54 ena vn 0.113034f
C55 vt 0 -2.338832f
C56 vpp 0 30.489046f
C57 vnn 0 31.37283f
C58 vinp 0 21.601118f
C59 vinn 0 22.277264f
C60 avss 0 37.106976f
C61 out 0 0.395015f
C62 n1 0 3.166643f
C63 avdd 0 0.387077p
C64 n0 0 2.028785f
C65 ena_b 0 1.545081f
C66 vm 0 10.557391f
C67 ibias 0 0.276354f
C68 ena 0 1.670602f
C69 vn 0 10.521617f
.ends

.subckt por_ana vin otrip_decoded[7] otrip_decoded[6] otrip_decoded[5] otrip_decoded[4]
+ otrip_decoded[3] otrip_decoded[2] otrip_decoded[1] otrip_decoded[0] vbg_1v2 avdd
+ itest avss ibg_200n force_pdnb dvdd dvss dcomp isrc_sel pwup_filt osc_ck osc_ena
+ porb_h por_unbuf por porb
Xsky130_fd_sc_hd__inv_16_3 sky130_fd_sc_hd__inv_4_4/Y dvss dvss dvdd dvdd por sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hvl__lsbufhv2lv_1_0 dcomp3v3 dvdd dvss dvss avdd avdd vl sky130_fd_sc_hvl__lsbufhv2lv_1
Xsky130_fd_sc_hvl__lsbufhv2lv_1_1 dcomp3v3uv dvdd dvss dvss avdd avdd sky130_fd_sc_hvl__lsbufhv2lv_1_1/X
+ sky130_fd_sc_hvl__lsbufhv2lv_1
Xrstring_mux_0 vin ibias_gen_0/ena rstring_mux_0/otrip_decoded_avdd[7] rstring_mux_0/otrip_decoded_avdd[6]
+ rstring_mux_0/otrip_decoded_avdd[3] rstring_mux_0/otrip_decoded_avdd[1] rstring_mux_0/m1_10352_4059#
+ rstring_mux_0/m1_24716_4059# rstring_mux_0/m1_10730_n3340# rstring_mux_0/m1_6572_4059#
+ rstring_mux_0/m1_12998_n3340# rstring_mux_0/m1_25850_n3340# rstring_mux_0/m1_12242_n3340#
+ rstring_mux_0/m1_12620_4059# rstring_mux_0/m1_3548_4059# rstring_mux_0/m1_8840_4059#
+ rstring_mux_0/m1_23204_4059# rstring_mux_0/m1_6194_n3340# rstring_mux_0/vtrip_decoded_avdd[3]
+ rstring_mux_0/m1_5060_4059# rstring_mux_0/m1_13376_4059# rstring_mux_0/m1_22826_n3340#
+ rstring_mux_0/m1_20558_n3340# rstring_mux_0/vtrip_decoded_avdd[1] rstring_mux_0/vtrip_decoded_b_avdd[0]
+ rstring_mux_0/m1_902_n3340# rstring_mux_0/m1_17156_4059# rstring_mux_0/m1_2036_4059#
+ rstring_mux_0/m1_19046_n3340# rstring_mux_0/vtrip7 rstring_mux_0/ena_b rstring_mux_0/m1_24338_n3340#
+ rstring_mux_0/vtrip5 rstring_mux_0/m1_2414_n3340# rstring_mux_0/vtop rstring_mux_0/m1_11864_4059#
+ rstring_mux_0/m1_21692_4059# rstring_mux_0/m1_7706_n3340# rstring_mux_0/m1_8084_4059#
+ rstring_mux_0/otrip_decoded_avdd[2] rstring_mux_0/otrip_decoded_avdd[4] rstring_mux_0/otrip_decoded_avdd[0]
+ rstring_mux_0/m1_21314_n3340# rstring_mux_0/m1_9218_n3340# comparator_0/vinn rstring_mux_0/m1_7328_4059#
+ rstring_mux_0/m1_11486_n3340# rstring_mux_0/m1_19802_n3340# rstring_mux_0/m1_1658_n3340#
+ rstring_mux_0/vtrip0 rstring_mux_0/vtrip_decoded_avdd[5] rstring_mux_0/m1_17534_n3340#
+ rstring_mux_0/vtrip_decoded_avdd[7] rstring_mux_0/vtrip2 rstring_mux_0/vtrip4 rstring_mux_0/m1_4304_4059#
+ rstring_mux_0/vtrip6 rstring_mux_0/m1_9596_4059# rstring_mux_0/m1_4682_n3340# rstring_mux_0/m1_3170_n3340#
+ rstring_mux_0/vtrip_decoded_avdd[2] rstring_mux_0/vtrip_decoded_avdd[4] rstring_mux_0/m1_25472_4059#
+ rstring_mux_0/vtrip_decoded_avdd[6] rstring_mux_0/vtrip3 rstring_mux_0/m1_5816_4059#
+ rstring_mux_0/m1_22070_n3340# avdd rstring_mux_0/vtrip_decoded_b_avdd[7] rstring_mux_0/vtrip_decoded_avdd[0]
+ rstring_mux_0/otrip_decoded_avdd[5] rstring_mux_0/vtrip1 avss rstring_mux
Xsky130_fd_sc_hvl__inv_4_0 sky130_fd_sc_hvl__inv_4_0/A avss avss avdd avdd sky130_fd_sc_hvl__inv_4_0/Y
+ sky130_fd_sc_hvl__inv_4
Xsky130_fd_sc_hd__inv_4_0 schmitt_trigger_0/out dvss dvss dvdd dvdd sky130_fd_sc_hd__inv_4_0/Y
+ sky130_fd_sc_hd__inv_4
Xsky130_fd_sc_hd__inv_4_1 sky130_fd_sc_hd__inv_4_2/Y dvss dvss dvdd dvdd sky130_fd_sc_hd__inv_4_1/Y
+ sky130_fd_sc_hd__inv_4
Xsky130_fd_sc_hd__inv_4_2 por_unbuf dvss dvss dvdd dvdd sky130_fd_sc_hd__inv_4_2/Y
+ sky130_fd_sc_hd__inv_4
Xschmitt_trigger_0 schmitt_trigger_0/in schmitt_trigger_0/out dvdd dvss schmitt_trigger_0/m
+ schmitt_trigger
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[0|0] otrip_decoded[0] dvdd dvss dvss avdd avdd rstring_mux_0/otrip_decoded_avdd[0]
+ sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[1|0] otrip_decoded[1] dvdd dvss dvss avdd avdd rstring_mux_0/otrip_decoded_avdd[1]
+ sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[0|1] otrip_decoded[2] dvdd dvss dvss avdd avdd rstring_mux_0/otrip_decoded_avdd[2]
+ sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[1|1] otrip_decoded[3] dvdd dvss dvss avdd avdd rstring_mux_0/otrip_decoded_avdd[3]
+ sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[0|2] otrip_decoded[4] dvdd dvss dvss avdd avdd rstring_mux_0/otrip_decoded_avdd[4]
+ sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[1|2] otrip_decoded[5] dvdd dvss dvss avdd avdd rstring_mux_0/otrip_decoded_avdd[5]
+ sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[0|3] otrip_decoded[6] dvdd dvss dvss avdd avdd rstring_mux_0/otrip_decoded_avdd[6]
+ sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[1|3] otrip_decoded[7] dvdd dvss dvss avdd avdd rstring_mux_0/otrip_decoded_avdd[7]
+ sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[0|4] dvss dvdd dvss dvss avdd avdd rstring_mux_0/vtrip_decoded_avdd[0]
+ sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[1|4] dvss dvdd dvss dvss avdd avdd rstring_mux_0/vtrip_decoded_avdd[1]
+ sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[0|5] dvss dvdd dvss dvss avdd avdd rstring_mux_0/vtrip_decoded_avdd[2]
+ sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[1|5] dvss dvdd dvss dvss avdd avdd rstring_mux_0/vtrip_decoded_avdd[3]
+ sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[0|6] dvss dvdd dvss dvss avdd avdd rstring_mux_0/vtrip_decoded_avdd[4]
+ sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[1|6] dvss dvdd dvss dvss avdd avdd rstring_mux_0/vtrip_decoded_avdd[5]
+ sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[0|7] dvss dvdd dvss dvss avdd avdd rstring_mux_0/vtrip_decoded_avdd[6]
+ sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[1|7] dvss dvdd dvss dvss avdd avdd rstring_mux_0/vtrip_decoded_avdd[7]
+ sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[0|8] force_pdnb dvdd dvss dvss avdd avdd ibias_gen_0/ena
+ sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[1|8] isrc_sel dvdd dvss dvss avdd avdd ibias_gen_0/isrc_sel
+ sky130_fd_sc_hvl__lsbuflv2hv_1
Xrc_osc_0 dvdd osc_ck osc_ena rc_osc_0/vr dvss rc_osc
Xsky130_fd_sc_hvl__lsbuflv2hv_1_1 por_unbuf dvdd dvss dvss avdd avdd sky130_fd_sc_hvl__inv_1_0/A
+ sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hd__inv_4_3 vl dvss dvss dvdd dvdd sky130_fd_sc_hd__inv_4_3/Y sky130_fd_sc_hd__inv_4
Xsky130_fd_sc_hd__inv_4_4 por_unbuf dvss dvss dvdd dvdd sky130_fd_sc_hd__inv_4_4/Y
+ sky130_fd_sc_hd__inv_4
Xsky130_fd_sc_hvl__inv_16_0 sky130_fd_sc_hvl__inv_4_0/Y avss avss avdd avdd porb_h
+ sky130_fd_sc_hvl__inv_16
Xsky130_fd_pr__res_xhigh_po_1p41_DVQADA_0 m1_n11325_2001# m1_n11325_2001# m1_n12081_2001#
+ m1_n10191_9400# m1_n13971_9400# m1_n14349_2001# m1_n12081_2001# vl m1_n12837_2001#
+ m1_n8301_2001# m1_n12837_2001# avss m1_n9435_9400# m1_n10947_9400# m1_n13215_9400#
+ m1_n13215_9400# m1_n8679_9400# m1_n10569_2001# m1_n9435_9400# m1_n13971_9400# m1_n10569_2001#
+ m1_n14727_9400# m1_n8301_2001# m1_n10947_9400# m1_n13593_2001# schmitt_trigger_0/in
+ m1_n11703_9400# m1_n8679_9400# m1_n9813_2001# m1_n9057_2001# m1_n9813_2001# m1_n7923_9400#
+ m1_n12459_9400# m1_n11703_9400# m1_n13593_2001# m1_n14727_9400# m1_n10191_9400#
+ m1_n14349_2001# m1_n9057_2001# m1_n7923_9400# m1_n12459_9400# sky130_fd_pr__res_xhigh_po_1p41_DVQADA
Xsky130_fd_pr__cap_mim_m3_2_LUWKLG_0 schmitt_trigger_0/in dvss sky130_fd_pr__cap_mim_m3_2_LUWKLG
Xibias_gen_0 ibias_gen_0/ibias0 itest ibias_gen_0/ibias1 ibg_200n vbg_1v2 ibias_gen_0/ve
+ ibias_gen_0/m1_7189_119# ibias_gen_0/m1_1897_119# ibias_gen_0/vstart ibias_gen_0/vr
+ ibias_gen_0/isrc_sel_b ibias_gen_0/m1_5677_119# ibias_gen_0/vp1 ibias_gen_0/m1_1141_119#
+ ibias_gen_0/ena_b ibias_gen_0/vp ibias_gen_0/ena ibias_gen_0/m1_385_119# ibias_gen_0/m1_2653_119#
+ ibias_gen_0/m1_4165_119# ibias_gen_0/isrc_sel ibias_gen_0/vn0 avdd avss ibias_gen_0/m1_763_7518#
+ ibias_gen_0/vp0 ibias_gen_0/vn1 ibias_gen
Xsky130_fd_pr__rf_pnp_05v5_W0p68L0p68_0 avss avss ibias_gen_0/ve avss sky130_fd_pr__rf_pnp_05v5_W0p68L0p68 m=1
Xsky130_fd_sc_hvl__inv_1_0 sky130_fd_sc_hvl__inv_1_0/A avss avss avdd avdd sky130_fd_sc_hvl__inv_4_0/A
+ sky130_fd_sc_hvl__inv_1
Xcomparator_0 ibias_gen_0/ibias1 dcomp3v3uv avss comparator_0/ena_b comparator_0/vt
+ vbg_1v2 comparator_0/n0 avss comparator_0/vpp comparator_0/vinn avdd comparator_0/vm
+ comparator_0/vn comparator_0/vnn comparator_0/n1 comparator
Xcomparator_1 ibias_gen_0/ibias0 dcomp3v3 ibias_gen_0/ena comparator_1/ena_b comparator_1/vt
+ vin comparator_1/n0 avss comparator_1/vpp vbg_1v2 avdd comparator_1/vm comparator_1/vn
+ comparator_1/vnn comparator_1/n1 comparator
Xsky130_fd_sc_hd__inv_16_0 sky130_fd_sc_hd__inv_4_0/Y dvss dvss dvdd dvdd pwup_filt
+ sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__inv_16_1 sky130_fd_sc_hd__inv_4_1/Y dvss dvss dvdd dvdd porb sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__inv_16_2 sky130_fd_sc_hd__inv_4_3/Y dvss dvss dvdd dvdd dcomp sky130_fd_sc_hd__inv_16
C0 dvss rstring_mux_0/vtrip0 3.056463f
C1 rc_osc_0/in comparator_0/vt 0.164658f
C2 rstring_mux_0/m1_22070_n3340# dvss 0.11558f
C3 dvss rstring_mux_0/vtrip_decoded_avdd[4] 0.593277f
C4 dvss ibias_gen_0/m1_4165_119# 0.137031f
C5 dvss porb 0.17194f
C6 rstring_mux_0/m1_24716_4059# dvss 0.157062f
C7 comparator_0/vinn rstring_mux_0/m1_4304_4059# 0.159467f
C8 ibias_gen_0/isrc_sel dcomp3v3 10.963935f
C9 dvss rstring_mux_0/m1_7328_4059# 0.12405f
C10 dvss comparator_0/vm 0.18333f
C11 dvss sky130_fd_sc_hvl__lsbufhv2lv_1_1/X 1.539706f
C12 schmitt_trigger_0/in rstring_mux_0/otrip_decoded_avdd[1] 0.556852f
C13 dvss ibias_gen_0/isrc_sel 0.544029f
C14 dvdd rstring_mux_0/vtop 0.177166f
C15 dvss rstring_mux_0/m1_4304_4059# 0.1412f
C16 vin comparator_1/vt 0.36298f
C17 comparator_0/vnn ibias_gen_0/ibias1 0.116472f
C18 ibias_gen_0/vp1 avdd -0.119038f
C19 dvss rstring_mux_0/m1_2414_n3340# 0.112505f
C20 dvdd sky130_fd_sc_hd__inv_4_4/Y 0.137857f
C21 avdd rstring_mux_0/vtrip_decoded_avdd[1] 1.321368f
C22 comparator_0/vinn comparator_0/n0 0.103671f
C23 ibias_gen_0/ena ibias_gen_0/vstart 0.293802f
C24 comparator_0/vn ibias_gen_0/ibias1 0.137125f
C25 por_unbuf schmitt_trigger_0/out 0.131748f
C26 vl dvdd 1.374402f
C27 schmitt_trigger_0/out schmitt_trigger_0/m 0.142691f
C28 comparator_0/vinn rstring_mux_0/m1_13376_4059# 0.154012f
C29 dvss comparator_0/n0 0.148095f
C30 comparator_1/vpp avdd -0.198399f
C31 rstring_mux_0/m1_20180_4059# dvss 0.150927f
C32 dvss ibias_gen_0/m1_5677_119# 0.144124f
C33 rstring_mux_0/vtrip_decoded_avdd[7] dvdd 0.289581f
C34 comparator_0/vinn rstring_mux_0/vtop 1.24609f
C35 dvss ibias_gen_0/m1_385_119# 0.111767f
C36 dvss rstring_mux_0/m1_13376_4059# 0.132297f
C37 rstring_mux_0/m1_26606_n3340# dvss 0.110111f
C38 rstring_mux_0/otrip_decoded_avdd[7] avdd 1.172732f
C39 ibias_gen_0/ena comparator_0/vnn 0.298208f
C40 ibias_gen_0/ena dvdd 0.351058f
C41 dvss rstring_mux_0/m1_9218_n3340# 0.118906f
C42 rstring_mux_0/otrip_decoded_avdd[1] rstring_mux_0/otrip_decoded_avdd[0] 3.164846f
C43 rstring_mux_0/vtrip_decoded_avdd[2] rstring_mux_0/vtrip_decoded_avdd[3] 1.699062f
C44 comparator_1/vt avdd -0.299234f
C45 dvss rstring_mux_0/vtop 8.409122f
C46 avdd rstring_mux_0/vtrip_decoded_avdd[5] 1.608562f
C47 comparator_1/vt vbg_1v2 0.218707f
C48 comparator_0/vinn rstring_mux_0/m1_17156_4059# 0.329592f
C49 dvss ibias_gen_0/ibias1 0.949401f
C50 vl dcomp3v3 10.054001f
C51 rstring_mux_0/m1_18290_n3340# dvss 0.1105f
C52 dvss sky130_fd_sc_hd__inv_4_4/Y 0.901102f
C53 dvss rstring_mux_0/m1_6194_n3340# 0.1105f
C54 dvdd rstring_mux_0/otrip_decoded_avdd[5] 0.423139f
C55 ibias_gen_0/ve avdd 8.371976f
C56 dvss rstring_mux_0/m1_11486_n3340# 0.1105f
C57 dcomp3v3uv ibias_gen_0/ena 0.508881f
C58 ibias_gen_0/ve vbg_1v2 2.022147f
C59 vl dvss 2.50144f
C60 dvss rstring_mux_0/m1_17156_4059# 0.139446f
C61 rstring_mux_0/vtrip_decoded_avdd[5] rstring_mux_0/vtrip_decoded_avdd[6] 1.257583f
C62 por dvss 0.177774f
C63 rstring_mux_0/vtrip_decoded_avdd[4] rstring_mux_0/vtrip_decoded_avdd[5] 2.208645f
C64 schmitt_trigger_0/in avdd 4.444283f
C65 ibias_gen_0/ena comparator_0/vinn 0.229267f
C66 comparator_0/vinn rstring_mux_0/vtrip4 0.113272f
C67 ibias_gen_0/vp dcomp3v3 0.494701f
C68 ibias_gen_0/ibias0 comparator_1/vnn 1.847506f
C69 vin rstring_mux_0/otrip_decoded_avdd[0] 0.330246f
C70 dvss rstring_mux_0/vtrip_decoded_avdd[7] 0.804244f
C71 dcomp3v3uv rstring_mux_0/otrip_decoded_avdd[5] 0.213252f
C72 ibias_gen_0/ena comparator_0/vpp 0.429225f
C73 dvss ibias_gen_0/ena 1.503252f
C74 dvss rstring_mux_0/vtrip4 2.979705f
C75 avdd rstring_mux_0/otrip_decoded_avdd[2] 0.880362f
C76 schmitt_trigger_0/in rstring_mux_0/vtrip_decoded_avdd[6] 0.211299f
C77 comparator_0/vinn rstring_mux_0/m1_8084_4059# 0.128847f
C78 comparator_1/vnn ibias_gen_0/ena 0.641406f
C79 sky130_fd_sc_hvl__inv_1_0/A dvss 0.134844f
C80 vin ibias_gen_0/vn1 0.823593f
C81 rstring_mux_0/vtrip_decoded_avdd[4] schmitt_trigger_0/in 0.158489f
C82 rstring_mux_0/m1_22826_n3340# dvss 0.1105f
C83 avdd rstring_mux_0/otrip_decoded_avdd[3] 1.073604f
C84 vin ibias_gen_0/vn0 0.111328f
C85 rstring_mux_0/m1_25472_4059# dvss 0.157062f
C86 ibias_gen_0/vp1 ibias_gen_0/ibias1 0.389737f
C87 ibias_gen_0/ena rstring_mux_0/vtrip_decoded_b_avdd[0] 0.100519f
C88 dvss rstring_mux_0/otrip_decoded_avdd[5] 0.832834f
C89 comparator_0/vinn rstring_mux_0/m1_5060_4059# 0.159467f
C90 dvss rstring_mux_0/m1_8084_4059# 0.540776f
C91 comparator_0/vinn rstring_mux_0/m1_10352_4059# 0.159467f
C92 avdd rstring_mux_0/otrip_decoded_avdd[4] 0.882012f
C93 rstring_mux_0/otrip_decoded_avdd[6] avdd 0.981291f
C94 avdd rstring_mux_0/vtrip_decoded_avdd[0] 0.946822f
C95 avdd rstring_mux_0/otrip_decoded_avdd[0] 0.596861f
C96 dvss rstring_mux_0/m1_5060_4059# 0.1412f
C97 dvss rstring_mux_0/m1_10352_4059# 0.1412f
C98 dcomp3v3uv dvdd 1.091701f
C99 ibias_gen_0/vp0 ibias_gen_0/ve 0.462312f
C100 ibias_gen_0/ena ibias_gen_0/vp1 0.114022f
C101 sky130_fd_sc_hvl__lsbufhv2lv_1_1/X rstring_mux_0/otrip_decoded_avdd[3] 1.379306f
C102 vl por_unbuf 0.129633f
C103 dvdd comparator_0/vinn 0.119454f
C104 ibias_gen_0/ibias0 comparator_1/vpp 1.31426f
C105 dvss rstring_mux_0/m1_3170_n3340# 0.109428f
C106 rstring_mux_0/vtrip_decoded_b_avdd[7] ibias_gen_0/ena 0.1256f
C107 dvdd dcomp3v3 1.10492f
C108 rstring_mux_0/vtrip_decoded_avdd[2] avdd 1.01317f
C109 comparator_0/vnn comparator_0/vpp -0.215697f
C110 rstring_mux_0/m1_20936_4059# dvss 0.144948f
C111 dvss ibias_gen_0/m1_6433_119# 0.137031f
C112 dvss ibias_gen_0/m1_1141_119# 0.137031f
C113 dvss comparator_0/vnn 13.870564f
C114 dvss dvdd 78.327576f
C115 ibias_gen_0/ibias0 comparator_1/vt 0.504594f
C116 comparator_1/vpp ibias_gen_0/ena 0.744362f
C117 rstring_mux_0/m1_21692_4059# dvss 0.157062f
C118 ibias_gen_0/ibias0 comparator_1/vn 0.310222f
C119 dvss sky130_fd_sc_hd__inv_4_1/Y 0.965214f
C120 dvss comparator_0/vn 0.329439f
C121 avdd rstring_mux_0/vtrip_decoded_avdd[3] 1.229798f
C122 rc_osc_0/in avdd 0.210176f
C123 rstring_mux_0/m1_19046_n3340# dvss 0.1105f
C124 comparator_0/vinn rstring_mux_0/m1_2036_4059# 0.159695f
C125 comparator_1/vt ibias_gen_0/ena 0.306813f
C126 dvss dcomp3v3uv 4.379798f
C127 dvss rstring_mux_0/m1_12242_n3340# 0.110499f
C128 vl schmitt_trigger_0/in 0.503663f
C129 ibias_gen_0/ena comparator_1/vn 0.153582f
C130 ibias_gen_0/m1_763_7518# ibias_gen_0/ibias1 0.134538f
C131 dvss comparator_0/vinn 16.246464f
C132 dvss rstring_mux_0/m1_2036_4059# 0.1412f
C133 rstring_mux_0/vtrip_decoded_avdd[4] rstring_mux_0/vtrip_decoded_avdd[3] 0.96514f
C134 dvss dcomp3v3 0.108037f
C135 comparator_0/vinn rstring_mux_0/vtrip6 0.179683f
C136 dvss dcomp 0.17772f
C137 dvss comparator_0/vpp 8.892797f
C138 avdd rstring_mux_0/otrip_decoded_avdd[1] 1.088785f
C139 rstring_mux_0/vtrip_decoded_avdd[7] schmitt_trigger_0/in 0.377385f
C140 dvss comparator_0/ena_b 0.173573f
C141 ibias_gen_0/ena schmitt_trigger_0/in 1.1842f
C142 comparator_0/vinn rstring_mux_0/vtrip2 0.228545f
C143 dvss rstring_mux_0/vtrip6 2.883271f
C144 comparator_0/vinn rstring_mux_0/m1_8840_4059# 0.159467f
C145 dvdd rstring_mux_0/vtrip_decoded_avdd[1] 0.335417f
C146 rstring_mux_0/m1_23582_n3340# dvss 0.1105f
C147 dvdd rc_osc_0/vr 0.342728f
C148 itest ibias_gen_0/ibias1 0.10252f
C149 rstring_mux_0/m1_26228_4059# dvss 0.157061f
C150 dvss rstring_mux_0/vtrip2 2.513916f
C151 schmitt_trigger_0/in rstring_mux_0/otrip_decoded_avdd[5] 0.101776f
C152 comparator_0/vinn rstring_mux_0/m1_5816_4059# 0.159467f
C153 dvss rstring_mux_0/m1_8840_4059# 0.148613f
C154 comparator_0/vinn rstring_mux_0/m1_11108_4059# 0.159467f
C155 ibias_gen_0/vn1 rstring_mux_0/vtop 0.192959f
C156 dcomp3v3uv ibias_gen_0/vp1 0.195351f
C157 vin avdd 2.390318f
C158 dvdd por_unbuf 1.084255f
C159 dcomp3v3uv rstring_mux_0/vtrip_decoded_avdd[1] 0.100293f
C160 vin vbg_1v2 3.662411f
C161 sky130_fd_sc_hd__inv_4_0/Y schmitt_trigger_0/out 0.14029f
C162 rstring_mux_0/m1_17912_4059# dvss 0.154064f
C163 rstring_mux_0/otrip_decoded_avdd[7] dvdd 0.291769f
C164 dvss rstring_mux_0/m1_5816_4059# 0.1412f
C165 dvss rstring_mux_0/m1_11108_4059# 0.1412f
C166 ibias_gen_0/vp1 dcomp3v3 0.543408f
C167 dvss rstring_mux_0/m1_6950_n3340# 0.1105f
C168 dvdd rstring_mux_0/vtrip_decoded_avdd[5] 0.324294f
C169 ibias_gen_0/ibias0 comparator_1/vm 0.155341f
C170 ibias_gen_0/ena rstring_mux_0/otrip_decoded_avdd[0] 0.821959f
C171 dvss ibias_gen_0/vp1 0.15897f
C172 ibias_gen_0/ena itest 0.154848f
C173 dvss rstring_mux_0/vtrip_decoded_avdd[1] 1.07926f
C174 rstring_mux_0/otrip_decoded_avdd[4] rstring_mux_0/otrip_decoded_avdd[5] 1.071892f
C175 comparator_0/vinn rstring_mux_0/vtrip1 0.318627f
C176 rstring_mux_0/otrip_decoded_avdd[6] rstring_mux_0/otrip_decoded_avdd[5] 0.257867f
C177 dvss rc_osc_0/vr -0.113725f
C178 dvss rstring_mux_0/m1_3926_n3340# 0.1105f
C179 ibias_gen_0/vn1 ibias_gen_0/ena 1.243157f
C180 schmitt_trigger_0/in comparator_0/vnn 0.268371f
C181 dvss ibias_gen_0/m1_1897_119# 0.137031f
C182 dvdd schmitt_trigger_0/in 0.873131f
C183 ibias_gen_0/ena ibias_gen_0/vn0 0.139772f
C184 avdd vbg_1v2 4.391585f
C185 dvss rstring_mux_0/vtrip1 1.877567f
C186 porb_h sky130_fd_sc_hvl__inv_4_0/Y 0.117022f
C187 dvss por_unbuf 3.598459f
C188 rstring_mux_0/m1_22448_4059# dvss 0.157061f
C189 comparator_1/vpp comparator_1/vnn -0.111946f
C190 comparator_1/vt dcomp3v3 2.363666f
C191 dvss rc_osc_0/m1_2270_n4# 0.150408f
C192 dvss schmitt_trigger_0/m 0.565618f
C193 dvss rstring_mux_0/otrip_decoded_avdd[7] 0.863725f
C194 dvss ibias_gen_0/m1_7189_119# 0.13632f
C195 dvdd rstring_mux_0/otrip_decoded_avdd[2] 0.255577f
C196 avdd rstring_mux_0/vtrip_decoded_avdd[6] 1.287716f
C197 rstring_mux_0/m1_19802_n3340# dvss 0.110499f
C198 comparator_0/vinn rstring_mux_0/m1_2792_4059# 0.159467f
C199 rstring_mux_0/vtrip_decoded_avdd[4] avdd 0.966219f
C200 dcomp3v3uv schmitt_trigger_0/in 0.122613f
C201 comparator_1/vnn comparator_1/vt -0.116128f
C202 comparator_1/n0 avdd -0.120008f
C203 dvss rstring_mux_0/vtrip_decoded_avdd[5] 0.875311f
C204 dvss rstring_mux_0/m1_12998_n3340# 0.1105f
C205 dvdd rstring_mux_0/otrip_decoded_avdd[3] 0.382485f
C206 vl rstring_mux_0/otrip_decoded_avdd[1] 0.145097f
C207 dvss rstring_mux_0/m1_2792_4059# 0.1412f
C208 avdd sky130_fd_sc_hvl__lsbufhv2lv_1_1/X 3.011103f
C209 schmitt_trigger_0/in comparator_0/vpp 0.250959f
C210 comparator_1/vnn ibias_gen_0/ve 1.565198f
C211 ibias_gen_0/isrc_sel avdd 3.510198f
C212 dcomp3v3uv rstring_mux_0/otrip_decoded_avdd[2] 0.375655f
C213 osc_ck dvdd 0.110121f
C214 dvdd rstring_mux_0/otrip_decoded_avdd[4] 0.266092f
C215 rstring_mux_0/otrip_decoded_avdd[6] dvdd 0.257138f
C216 dvdd rstring_mux_0/vtrip_decoded_avdd[0] 0.275187f
C217 dvdd rstring_mux_0/otrip_decoded_avdd[0] 0.197825f
C218 dvss schmitt_trigger_0/in 2.534112f
C219 dvdd rstring_mux_0/m1_7706_n3340# 0.407976f
C220 dvss comparator_0/vt 7.298046f
C221 dcomp3v3uv rstring_mux_0/otrip_decoded_avdd[3] 0.156703f
C222 dvss rstring_mux_0/m1_16778_n3340# 0.1105f
C223 ibias_gen_0/ena rstring_mux_0/otrip_decoded_avdd[1] 0.173335f
C224 comparator_0/vinn rstring_mux_0/m1_9596_4059# 0.159467f
C225 rstring_mux_0/m1_24338_n3340# dvss 0.1105f
C226 rstring_mux_0/otrip_decoded_avdd[6] dcomp3v3uv 0.148623f
C227 dcomp3v3uv rstring_mux_0/vtrip_decoded_avdd[0] 0.497383f
C228 dvss rstring_mux_0/otrip_decoded_avdd[2] 0.518951f
C229 comparator_0/vinn rstring_mux_0/m1_6572_4059# 0.159467f
C230 dvss rstring_mux_0/m1_9596_4059# 0.142297f
C231 ibias_gen_0/ibias0 vin 0.543516f
C232 rstring_mux_0/ena_b dvss 0.574124f
C233 dvdd rstring_mux_0/vtrip_decoded_avdd[2] 0.279976f
C234 comparator_0/vinn rstring_mux_0/m1_11864_4059# 0.159467f
C235 comparator_0/n0 vbg_1v2 0.16272f
C236 dvss rstring_mux_0/otrip_decoded_avdd[3] 0.782358f
C237 ibias_gen_0/vp0 avdd -0.516263f
C238 rstring_mux_0/m1_18668_4059# dvss 0.154064f
C239 dvss rstring_mux_0/m1_6572_4059# 0.1412f
C240 por_unbuf schmitt_trigger_0/m 0.13807f
C241 dcomp3v3uv ibias_gen_0/vn1 1.835448f
C242 ibias_gen_0/vp vin 0.362615f
C243 dvss rstring_mux_0/otrip_decoded_avdd[4] 0.366785f
C244 dvss rstring_mux_0/otrip_decoded_avdd[6] 0.42164f
C245 dvss rstring_mux_0/m1_11864_4059# 0.1412f
C246 dvss ibias_gen_0/m1_3409_119# 0.137031f
C247 dvss rstring_mux_0/vtrip_decoded_avdd[0] 0.60324f
C248 vin ibias_gen_0/ena 2.348609f
C249 rstring_mux_0/m1_25094_n3340# dvss 0.1105f
C250 avdd rstring_mux_0/vtop 1.571107f
C251 dvss rstring_mux_0/otrip_decoded_avdd[0] 0.396704f
C252 dvss rstring_mux_0/m1_7706_n3340# 0.475412f
C253 avdd ibias_gen_0/ibias1 7.06357f
C254 dvdd rstring_mux_0/vtrip_decoded_avdd[3] 0.517826f
C255 dcomp3v3uv rstring_mux_0/vtrip_decoded_avdd[2] 0.359441f
C256 schmitt_trigger_0/in rstring_mux_0/vtrip_decoded_avdd[1] 0.133642f
C257 comparator_0/vinn rstring_mux_0/vtrip5 0.205628f
C258 comparator_1/vpp ibias_gen_0/ve 1.055305f
C259 vl avdd 2.826377f
C260 dvss rstring_mux_0/m1_4682_n3340# 0.1105f
C261 dvss ibias_gen_0/vn1 1.353608f
C262 dvss rstring_mux_0/m1_9974_n3340# 0.1105f
C263 ibias_gen_0/ibias0 avdd 1.930784f
C264 dvss ibias_gen_0/m1_2653_119# 0.137031f
C265 avdd sky130_fd_sc_hvl__inv_4_0/A 0.133985f
C266 dvss rstring_mux_0/vtrip5 2.392901f
C267 ibias_gen_0/ibias0 vbg_1v2 2.287594f
C268 dvss rstring_mux_0/vtrip_decoded_avdd[2] 0.89944f
C269 ibias_gen_0/ve comparator_1/vt 0.467296f
C270 rstring_mux_0/vtrip_decoded_avdd[7] avdd 1.166121f
C271 dvdd rstring_mux_0/otrip_decoded_avdd[1] 0.266224f
C272 rstring_mux_0/m1_23204_4059# dvss 0.157062f
C273 schmitt_trigger_0/in schmitt_trigger_0/m 0.105255f
C274 ibias_gen_0/ve comparator_1/vn 0.219066f
C275 ibias_gen_0/isrc_sel ibias_gen_0/isrc_sel_b -0.129258f
C276 ibias_gen_0/vp avdd -0.512519f
C277 rstring_mux_0/otrip_decoded_avdd[7] schmitt_trigger_0/in 0.12621f
C278 ibias_gen_0/ena avdd 9.272375f
C279 rc_osc_0/in comparator_0/vinn 0.174353f
C280 ibias_gen_0/vp vbg_1v2 0.379191f
C281 sky130_fd_sc_hvl__inv_1_0/A avdd 0.25195f
C282 ibias_gen_0/ena vbg_1v2 0.553772f
C283 rstring_mux_0/m1_20558_n3340# dvss 0.1105f
C284 ibias_gen_0/ibias0 comparator_1/n0 0.172673f
C285 comparator_0/vinn rstring_mux_0/m1_1280_4059# 0.161624f
C286 schmitt_trigger_0/in rstring_mux_0/vtrip_decoded_avdd[5] 0.174324f
C287 sky130_fd_sc_hd__inv_4_3/Y dvdd 0.127361f
C288 rstring_mux_0/vtrip_decoded_avdd[7] rstring_mux_0/vtrip_decoded_avdd[6] 2.980441f
C289 dvss rstring_mux_0/vtrip_decoded_avdd[3] 0.959662f
C290 rstring_mux_0/vtrip_decoded_avdd[1] rstring_mux_0/vtrip_decoded_avdd[0] 1.18814f
C291 vl sky130_fd_sc_hvl__lsbufhv2lv_1_1/X 0.799667f
C292 avdd rstring_mux_0/otrip_decoded_avdd[5] 1.176434f
C293 rstring_mux_0/m1_21314_n3340# dvss 0.1105f
C294 vl ibias_gen_0/isrc_sel 0.171709f
C295 dvss rstring_mux_0/m1_1280_4059# 0.126012f
C296 ibias_gen_0/ena comparator_1/n0 0.123113f
C297 vin dvdd 0.119455f
C298 comparator_0/vinn rstring_mux_0/m1_3548_4059# 0.159467f
C299 dvss rstring_mux_0/otrip_decoded_avdd[1] 0.75323f
C300 rstring_mux_0/otrip_decoded_avdd[7] rstring_mux_0/otrip_decoded_avdd[6] 1.047274f
C301 ibias_gen_0/vp ibias_gen_0/isrc_sel -0.287702f
C302 rstring_mux_0/otrip_decoded_avdd[7] rstring_mux_0/vtrip_decoded_avdd[0] 0.25154f
C303 dvss rstring_mux_0/m1_3548_4059# 0.1412f
C304 ibias_gen_0/m1_385_119# ibias_gen_0/ibias1 0.311542f
C305 ibias_gen_0/isrc_sel ibias_gen_0/ena 0.563816f
C306 dvss pwup_filt 0.14947f
C307 ibias_gen_0/vp0 ibias_gen_0/ibias1 0.954291f
C308 rstring_mux_0/vtrip_decoded_avdd[2] rstring_mux_0/vtrip_decoded_avdd[1] 0.535743f
C309 dvss rstring_mux_0/m1_1658_n3340# 0.1105f
C310 dvdd sky130_fd_sc_hd__inv_4_0/Y 0.168709f
C311 schmitt_trigger_0/in rstring_mux_0/otrip_decoded_avdd[2] 0.10426f
C312 dvss rstring_mux_0/m1_902_n3340# 0.110092f
C313 dvdd schmitt_trigger_0/out 0.368019f
C314 dvss sky130_fd_sc_hd__inv_4_3/Y 0.908573f
C315 schmitt_trigger_0/in rstring_mux_0/otrip_decoded_avdd[3] 0.117015f
C316 dvss sky130_fd_sc_hd__inv_4_2/Y 0.291792f
C317 comparator_0/vinn rstring_mux_0/m1_12620_4059# 0.157512f
C318 dvdd avdd 17.440788f
C319 rstring_mux_0/m1_19424_4059# dvss 0.154064f
C320 dvss ibias_gen_0/m1_4921_119# 0.137031f
C321 schmitt_trigger_0/in rstring_mux_0/otrip_decoded_avdd[4] 0.101976f
C322 vl ibias_gen_0/ibias1 0.261037f
C323 dvss vin 1.825811f
C324 rstring_mux_0/otrip_decoded_avdd[6] schmitt_trigger_0/in 0.105908f
C325 schmitt_trigger_0/in rstring_mux_0/vtrip_decoded_avdd[0] 0.128751f
C326 dvss rstring_mux_0/m1_12620_4059# 0.137708f
C327 rstring_mux_0/m1_25850_n3340# dvss 0.1105f
C328 ibias_gen_0/m1_385_119# ibias_gen_0/ena 0.294281f
C329 schmitt_trigger_0/in rstring_mux_0/otrip_decoded_avdd[0] 0.260407f
C330 rstring_mux_0/otrip_decoded_avdd[2] rstring_mux_0/otrip_decoded_avdd[3] 1.343758f
C331 ibias_gen_0/vp0 ibias_gen_0/ena 0.530637f
C332 ibias_gen_0/ve comparator_1/vm 0.263306f
C333 dvss rstring_mux_0/m1_8462_n3340# 0.142178f
C334 dvss comparator_0/n1 0.251619f
C335 dvdd rstring_mux_0/vtrip_decoded_avdd[6] 0.309916f
C336 ibias_gen_0/ena ibias_gen_0/isrc_sel_b 0.507252f
C337 ibias_gen_0/ve ibias_gen_0/vn0 0.428899f
C338 rstring_mux_0/vtrip_decoded_avdd[4] dvdd 0.669746f
C339 dcomp3v3uv avdd 2.796168f
C340 comparator_0/vinn rstring_mux_0/vtrip7 0.446279f
C341 ibias_gen_0/vp ibias_gen_0/ibias1 0.864109f
C342 dvss sky130_fd_sc_hd__inv_4_0/Y 0.880299f
C343 dcomp3v3uv vbg_1v2 0.3098f
C344 rstring_mux_0/m1_17534_n3340# dvss 0.1105f
C345 ibias_gen_0/ena ibias_gen_0/ibias1 2.329607f
C346 dvss rstring_mux_0/m1_5438_n3340# 0.1105f
C347 dvdd rstring_mux_0/m1_7328_4059# 0.431259f
C348 comparator_0/vinn avdd 1.437882f
C349 dvss schmitt_trigger_0/out 1.177791f
C350 dvss rstring_mux_0/m1_10730_n3340# 0.1105f
C351 rstring_mux_0/otrip_decoded_avdd[4] rstring_mux_0/otrip_decoded_avdd[3] 0.421114f
C352 comparator_0/vinn rstring_mux_0/vtrip3 0.342375f
C353 avdd dcomp3v3 3.699368f
C354 comparator_0/vinn vbg_1v2 0.304227f
C355 rstring_mux_0/vtrip_decoded_avdd[2] schmitt_trigger_0/in 0.137711f
C356 avdd comparator_0/vpp -0.101205f
C357 dvss rstring_mux_0/vtrip7 2.283851f
C358 vl ibias_gen_0/vp 0.599776f
C359 dvdd sky130_fd_sc_hvl__lsbufhv2lv_1_1/X 0.83762f
C360 dcomp3v3uv rstring_mux_0/vtrip_decoded_avdd[6] 0.194356f
C361 ibias_gen_0/isrc_sel dvdd 0.175734f
C362 dcomp3v3uv rstring_mux_0/vtrip_decoded_avdd[4] 0.249577f
C363 rstring_mux_0/m1_23960_4059# dvss 0.157061f
C364 dvss avdd 46.30195f
C365 ibias_gen_0/ibias0 ibias_gen_0/ena 1.050499f
C366 dvss rstring_mux_0/vtrip3 1.861528f
C367 ibias_gen_0/vp0 ibias_gen_0/vstart -0.124456f
C368 dvss vbg_1v2 5.71504f
C369 comparator_0/vinn rstring_mux_0/vtrip0 0.214256f
C370 rstring_mux_0/vtrip_decoded_avdd[7] ibias_gen_0/ena 1.915045f
C371 comparator_1/vnn vbg_1v2 0.46016f
C372 schmitt_trigger_0/in rstring_mux_0/vtrip_decoded_avdd[3] 0.14576f
C373 dcomp3v3uv sky130_fd_sc_hvl__lsbufhv2lv_1_1/X 2.568928f
C374 ibias_gen_0/vp ibias_gen_0/ena 0.600369f
C375 comparator_1/n0 dcomp3v3 0.556901f
C376 comparator_0/vinn rstring_mux_0/m1_7328_4059# 0.128847f
C377 dvss rstring_mux_0/vtrip_decoded_avdd[6] 0.490514f
C378 pwup_filt sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.104973f
C379 comparator_1/vt sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 -5.980006f
C380 comparator_1/vpp sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 31.232635f
C381 comparator_1/vnn sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 31.715967f
C382 vin sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 33.35816f
C383 dcomp3v3 sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 2.798703f
C384 comparator_1/n1 sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 4.68235f
C385 comparator_1/n0 sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 2.878679f
C386 comparator_1/ena_b sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 2.364393f
C387 comparator_1/vm sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 14.965508f
C388 ibias_gen_0/ibias0 sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 1.54151f
C389 comparator_1/vn sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 15.289467f
C390 comparator_0/vt sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 -5.846239f
C391 comparator_0/vpp sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 31.815475f
C392 comparator_0/vnn sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 32.259075f
C393 vbg_1v2 sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 53.08963f
C394 dcomp3v3uv sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 6.407106f
C395 comparator_0/n1 sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 4.683574f
C396 avdd sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 3.613298p
C397 comparator_0/n0 sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 3.13703f
C398 comparator_0/ena_b sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 2.354586f
C399 comparator_0/vm sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 15.008218f
C400 ibias_gen_0/ibias1 sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 5.208468f
C401 comparator_0/vn sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 15.363231f
C402 ibias_gen_0/ena_b sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 3.86876f
C403 itest sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.310141f
C404 ibias_gen_0/vp1 sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 4.795395f
C405 ibias_gen_0/vn1 sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 32.751534f
C406 ibias_gen_0/sky130_fd_pr__pfet_g5v0d10v5_7JLQGA_0/a_594_n500# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.101769f
C407 ibias_gen_0/sky130_fd_pr__pfet_g5v0d10v5_7JLQGA_0/a_n652_n500# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.101769f
C408 ibias_gen_0/vr sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 1.530451f
C409 ibias_gen_0/m1_7189_119# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 1.002334f
C410 ibias_gen_0/m1_6811_7518# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.862163f
C411 ibias_gen_0/m1_6433_119# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.861757f
C412 ibias_gen_0/m1_6055_7518# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.862163f
C413 ibias_gen_0/m1_5677_119# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.861757f
C414 ibias_gen_0/m1_5299_7518# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.862163f
C415 ibias_gen_0/m1_4921_119# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.861757f
C416 ibias_gen_0/m1_4543_7518# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.862163f
C417 ibias_gen_0/m1_4165_119# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.861757f
C418 ibias_gen_0/m1_3787_7518# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.862163f
C419 ibias_gen_0/m1_3409_119# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.861757f
C420 ibias_gen_0/m1_3031_7518# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.862163f
C421 ibias_gen_0/m1_2653_119# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.861757f
C422 ibias_gen_0/m1_2275_7518# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.862163f
C423 ibias_gen_0/m1_1897_119# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.861757f
C424 ibias_gen_0/m1_1519_7518# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.861301f
C425 ibias_gen_0/m1_1141_119# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.861757f
C426 ibias_gen_0/m1_763_7518# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.8557f
C427 ibias_gen_0/m1_385_119# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 1.021289f
C428 ibias_gen_0/ve sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 12.781865f
C429 ibg_200n sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.542864f
C430 ibias_gen_0/sky130_fd_pr__nfet_g5v0d10v5_EC8RE7_1/a_1306_n500# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.137397f $ **FLOATING
C431 ibias_gen_0/vp sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 6.523855f
C432 ibias_gen_0/vp0 sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 7.145138f
C433 ibias_gen_0/vstart sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 1.049887f
C434 ibias_gen_0/vn0 sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 15.506374f
C435 ibias_gen_0/ena sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 22.176567f
C436 ibias_gen_0/isrc_sel sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 5.129799f
C437 ibias_gen_0/isrc_sel_b sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 3.71774f
C438 m1_n7923_9400# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 1.224334f
C439 m1_n8301_2001# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.963111f
C440 m1_n8679_9400# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.962995f
C441 m1_n9057_2001# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.962942f
C442 m1_n9435_9400# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.962914f
C443 m1_n9813_2001# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.962914f
C444 m1_n10191_9400# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.962914f
C445 m1_n10569_2001# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.962914f
C446 m1_n10947_9400# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.962914f
C447 m1_n11325_2001# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.962914f
C448 m1_n11703_9400# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.962914f
C449 m1_n12081_2001# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.962914f
C450 m1_n12459_9400# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.962914f
C451 m1_n12837_2001# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.962914f
C452 m1_n13215_9400# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.962914f
C453 m1_n13593_2001# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.962942f
C454 m1_n13971_9400# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.965921f
C455 m1_n14349_2001# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.963111f
C456 m1_n14727_9400# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 1.247597f
C457 porb_h sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.193097f
C458 sky130_fd_sc_hvl__inv_4_0/Y sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 3.702777f
C459 sky130_fd_sc_hd__inv_4_4/Y sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.560331f
C460 sky130_fd_sc_hd__inv_4_3/Y sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.540491f
C461 sky130_fd_sc_hvl__inv_1_0/A sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 4.755877f
C462 sky130_fd_sc_hvl__lsbuflv2hv_1_1/a_772_151# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 1.04864f $ **FLOATING
C463 sky130_fd_sc_hvl__lsbuflv2hv_1_1/a_1197_107# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.25514f $ **FLOATING
C464 sky130_fd_sc_hvl__lsbuflv2hv_1_1/a_1711_885# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.339894f $ **FLOATING
C465 sky130_fd_sc_hvl__lsbuflv2hv_1_1/a_504_1221# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.834376f $ **FLOATING
C466 sky130_fd_sc_hvl__lsbuflv2hv_1_1/a_404_1133# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 1.44294f $ **FLOATING
C467 rc_osc_0/n sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.962242f
C468 rc_osc_0/ena_b sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.185393f
C469 osc_ena sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.348082f
C470 dvdd sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.312573p
C471 dvss sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.27171p
C472 rc_osc_0/m sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.458106f
C473 rc_osc_0/in sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 18.20599f
C474 rc_osc_0/vr sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.974916f
C475 osc_ck sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.231709f
C476 rc_osc_0/m1_25146_n1894# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.830903f
C477 rc_osc_0/m1_2270_n1516# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.690318f
C478 rc_osc_0/m1_25146_n1138# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.687159f
C479 rc_osc_0/m1_2270_n760# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.690318f
C480 rc_osc_0/m1_25146_n382# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.687159f
C481 rc_osc_0/m1_2270_n4# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.690318f
C482 rc_osc_0/m1_25146_374# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.687159f
C483 rc_osc_0/m1_2270_752# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.690318f
C484 rc_osc_0/m1_25146_1130# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.830903f
C485 isrc_sel sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.339407f
C486 sky130_fd_sc_hvl__lsbuflv2hv_1_0[1|8]/a_772_151# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 1.04864f $ **FLOATING
C487 sky130_fd_sc_hvl__lsbuflv2hv_1_0[1|8]/a_1197_107# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.25514f $ **FLOATING
C488 sky130_fd_sc_hvl__lsbuflv2hv_1_0[1|8]/a_1711_885# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.339894f $ **FLOATING
C489 sky130_fd_sc_hvl__lsbuflv2hv_1_0[1|8]/a_504_1221# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.834376f $ **FLOATING
C490 sky130_fd_sc_hvl__lsbuflv2hv_1_0[1|8]/a_404_1133# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 1.44294f $ **FLOATING
C491 force_pdnb sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.328995f
C492 sky130_fd_sc_hvl__lsbuflv2hv_1_0[0|8]/a_772_151# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 1.04864f $ **FLOATING
C493 sky130_fd_sc_hvl__lsbuflv2hv_1_0[0|8]/a_1197_107# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.25514f $ **FLOATING
C494 sky130_fd_sc_hvl__lsbuflv2hv_1_0[0|8]/a_1711_885# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.339894f $ **FLOATING
C495 sky130_fd_sc_hvl__lsbuflv2hv_1_0[0|8]/a_504_1221# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.834376f $ **FLOATING
C496 sky130_fd_sc_hvl__lsbuflv2hv_1_0[0|8]/a_404_1133# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 1.44294f $ **FLOATING
C497 sky130_fd_sc_hvl__lsbuflv2hv_1_0[1|7]/a_772_151# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 1.04864f $ **FLOATING
C498 sky130_fd_sc_hvl__lsbuflv2hv_1_0[1|7]/a_1197_107# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.25514f $ **FLOATING
C499 sky130_fd_sc_hvl__lsbuflv2hv_1_0[1|7]/a_1711_885# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.339894f $ **FLOATING
C500 sky130_fd_sc_hvl__lsbuflv2hv_1_0[1|7]/a_504_1221# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.834376f $ **FLOATING
C501 sky130_fd_sc_hvl__lsbuflv2hv_1_0[1|7]/a_404_1133# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 1.44294f $ **FLOATING
C502 sky130_fd_sc_hvl__lsbuflv2hv_1_0[0|7]/a_772_151# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 1.04864f $ **FLOATING
C503 sky130_fd_sc_hvl__lsbuflv2hv_1_0[0|7]/a_1197_107# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.25514f $ **FLOATING
C504 sky130_fd_sc_hvl__lsbuflv2hv_1_0[0|7]/a_1711_885# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.339894f $ **FLOATING
C505 sky130_fd_sc_hvl__lsbuflv2hv_1_0[0|7]/a_504_1221# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.834376f $ **FLOATING
C506 sky130_fd_sc_hvl__lsbuflv2hv_1_0[0|7]/a_404_1133# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 1.44294f $ **FLOATING
C507 sky130_fd_sc_hvl__lsbuflv2hv_1_0[1|6]/a_772_151# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 1.04864f $ **FLOATING
C508 sky130_fd_sc_hvl__lsbuflv2hv_1_0[1|6]/a_1197_107# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.25514f $ **FLOATING
C509 sky130_fd_sc_hvl__lsbuflv2hv_1_0[1|6]/a_1711_885# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.339894f $ **FLOATING
C510 sky130_fd_sc_hvl__lsbuflv2hv_1_0[1|6]/a_504_1221# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.834376f $ **FLOATING
C511 sky130_fd_sc_hvl__lsbuflv2hv_1_0[1|6]/a_404_1133# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 1.44294f $ **FLOATING
C512 sky130_fd_sc_hvl__lsbuflv2hv_1_0[0|6]/a_772_151# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 1.04864f $ **FLOATING
C513 sky130_fd_sc_hvl__lsbuflv2hv_1_0[0|6]/a_1197_107# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.25514f $ **FLOATING
C514 sky130_fd_sc_hvl__lsbuflv2hv_1_0[0|6]/a_1711_885# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.339894f $ **FLOATING
C515 sky130_fd_sc_hvl__lsbuflv2hv_1_0[0|6]/a_504_1221# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.834376f $ **FLOATING
C516 sky130_fd_sc_hvl__lsbuflv2hv_1_0[0|6]/a_404_1133# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 1.44294f $ **FLOATING
C517 sky130_fd_sc_hvl__lsbuflv2hv_1_0[1|5]/a_772_151# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 1.04864f $ **FLOATING
C518 sky130_fd_sc_hvl__lsbuflv2hv_1_0[1|5]/a_1197_107# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.25514f $ **FLOATING
C519 sky130_fd_sc_hvl__lsbuflv2hv_1_0[1|5]/a_1711_885# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.339894f $ **FLOATING
C520 sky130_fd_sc_hvl__lsbuflv2hv_1_0[1|5]/a_504_1221# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.834376f $ **FLOATING
C521 sky130_fd_sc_hvl__lsbuflv2hv_1_0[1|5]/a_404_1133# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 1.44294f $ **FLOATING
C522 sky130_fd_sc_hvl__lsbuflv2hv_1_0[0|5]/a_772_151# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 1.04864f $ **FLOATING
C523 sky130_fd_sc_hvl__lsbuflv2hv_1_0[0|5]/a_1197_107# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.25514f $ **FLOATING
C524 sky130_fd_sc_hvl__lsbuflv2hv_1_0[0|5]/a_1711_885# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.339894f $ **FLOATING
C525 sky130_fd_sc_hvl__lsbuflv2hv_1_0[0|5]/a_504_1221# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.834376f $ **FLOATING
C526 sky130_fd_sc_hvl__lsbuflv2hv_1_0[0|5]/a_404_1133# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 1.44294f $ **FLOATING
C527 sky130_fd_sc_hvl__lsbuflv2hv_1_0[1|4]/a_772_151# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 1.04864f $ **FLOATING
C528 sky130_fd_sc_hvl__lsbuflv2hv_1_0[1|4]/a_1197_107# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.25514f $ **FLOATING
C529 sky130_fd_sc_hvl__lsbuflv2hv_1_0[1|4]/a_1711_885# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.339894f $ **FLOATING
C530 sky130_fd_sc_hvl__lsbuflv2hv_1_0[1|4]/a_504_1221# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.834376f $ **FLOATING
C531 sky130_fd_sc_hvl__lsbuflv2hv_1_0[1|4]/a_404_1133# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 1.44294f $ **FLOATING
C532 sky130_fd_sc_hvl__lsbuflv2hv_1_0[0|4]/a_772_151# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 1.04864f $ **FLOATING
C533 sky130_fd_sc_hvl__lsbuflv2hv_1_0[0|4]/a_1197_107# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.25514f $ **FLOATING
C534 sky130_fd_sc_hvl__lsbuflv2hv_1_0[0|4]/a_1711_885# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.339894f $ **FLOATING
C535 sky130_fd_sc_hvl__lsbuflv2hv_1_0[0|4]/a_504_1221# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.834376f $ **FLOATING
C536 sky130_fd_sc_hvl__lsbuflv2hv_1_0[0|4]/a_404_1133# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 1.44294f $ **FLOATING
C537 otrip_decoded[7] sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.33104f
C538 sky130_fd_sc_hvl__lsbuflv2hv_1_0[1|3]/a_772_151# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 1.04864f $ **FLOATING
C539 sky130_fd_sc_hvl__lsbuflv2hv_1_0[1|3]/a_1197_107# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.25514f $ **FLOATING
C540 sky130_fd_sc_hvl__lsbuflv2hv_1_0[1|3]/a_1711_885# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.339894f $ **FLOATING
C541 sky130_fd_sc_hvl__lsbuflv2hv_1_0[1|3]/a_504_1221# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.834376f $ **FLOATING
C542 sky130_fd_sc_hvl__lsbuflv2hv_1_0[1|3]/a_404_1133# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 1.44294f $ **FLOATING
C543 otrip_decoded[6] sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.329592f
C544 sky130_fd_sc_hvl__lsbuflv2hv_1_0[0|3]/a_772_151# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 1.04864f $ **FLOATING
C545 sky130_fd_sc_hvl__lsbuflv2hv_1_0[0|3]/a_1197_107# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.25514f $ **FLOATING
C546 sky130_fd_sc_hvl__lsbuflv2hv_1_0[0|3]/a_1711_885# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.339894f $ **FLOATING
C547 sky130_fd_sc_hvl__lsbuflv2hv_1_0[0|3]/a_504_1221# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.834376f $ **FLOATING
C548 sky130_fd_sc_hvl__lsbuflv2hv_1_0[0|3]/a_404_1133# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 1.44294f $ **FLOATING
C549 otrip_decoded[5] sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.329062f
C550 sky130_fd_sc_hvl__lsbuflv2hv_1_0[1|2]/a_772_151# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 1.04864f $ **FLOATING
C551 sky130_fd_sc_hvl__lsbuflv2hv_1_0[1|2]/a_1197_107# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.25514f $ **FLOATING
C552 sky130_fd_sc_hvl__lsbuflv2hv_1_0[1|2]/a_1711_885# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.339894f $ **FLOATING
C553 sky130_fd_sc_hvl__lsbuflv2hv_1_0[1|2]/a_504_1221# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.834376f $ **FLOATING
C554 sky130_fd_sc_hvl__lsbuflv2hv_1_0[1|2]/a_404_1133# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 1.44294f $ **FLOATING
C555 otrip_decoded[4] sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.336087f
C556 sky130_fd_sc_hvl__lsbuflv2hv_1_0[0|2]/a_772_151# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 1.04864f $ **FLOATING
C557 sky130_fd_sc_hvl__lsbuflv2hv_1_0[0|2]/a_1197_107# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.25514f $ **FLOATING
C558 sky130_fd_sc_hvl__lsbuflv2hv_1_0[0|2]/a_1711_885# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.339894f $ **FLOATING
C559 sky130_fd_sc_hvl__lsbuflv2hv_1_0[0|2]/a_504_1221# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.834376f $ **FLOATING
C560 sky130_fd_sc_hvl__lsbuflv2hv_1_0[0|2]/a_404_1133# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 1.44294f $ **FLOATING
C561 otrip_decoded[3] sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.328176f
C562 sky130_fd_sc_hvl__lsbuflv2hv_1_0[1|1]/a_772_151# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 1.04864f $ **FLOATING
C563 sky130_fd_sc_hvl__lsbuflv2hv_1_0[1|1]/a_1197_107# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.25514f $ **FLOATING
C564 sky130_fd_sc_hvl__lsbuflv2hv_1_0[1|1]/a_1711_885# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.339894f $ **FLOATING
C565 sky130_fd_sc_hvl__lsbuflv2hv_1_0[1|1]/a_504_1221# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.834376f $ **FLOATING
C566 sky130_fd_sc_hvl__lsbuflv2hv_1_0[1|1]/a_404_1133# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 1.44294f $ **FLOATING
C567 otrip_decoded[2] sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.333543f
C568 sky130_fd_sc_hvl__lsbuflv2hv_1_0[0|1]/a_772_151# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 1.04864f $ **FLOATING
C569 sky130_fd_sc_hvl__lsbuflv2hv_1_0[0|1]/a_1197_107# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.25514f $ **FLOATING
C570 sky130_fd_sc_hvl__lsbuflv2hv_1_0[0|1]/a_1711_885# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.339894f $ **FLOATING
C571 sky130_fd_sc_hvl__lsbuflv2hv_1_0[0|1]/a_504_1221# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.834376f $ **FLOATING
C572 sky130_fd_sc_hvl__lsbuflv2hv_1_0[0|1]/a_404_1133# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 1.44294f $ **FLOATING
C573 otrip_decoded[1] sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.335439f
C574 sky130_fd_sc_hvl__lsbuflv2hv_1_0[1|0]/a_772_151# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 1.04864f $ **FLOATING
C575 sky130_fd_sc_hvl__lsbuflv2hv_1_0[1|0]/a_1197_107# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.25514f $ **FLOATING
C576 sky130_fd_sc_hvl__lsbuflv2hv_1_0[1|0]/a_1711_885# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.339913f $ **FLOATING
C577 sky130_fd_sc_hvl__lsbuflv2hv_1_0[1|0]/a_504_1221# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.83443f $ **FLOATING
C578 sky130_fd_sc_hvl__lsbuflv2hv_1_0[1|0]/a_404_1133# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 1.443208f $ **FLOATING
C579 otrip_decoded[0] sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.336251f
C580 sky130_fd_sc_hvl__lsbuflv2hv_1_0[0|0]/a_772_151# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 1.04864f $ **FLOATING
C581 sky130_fd_sc_hvl__lsbuflv2hv_1_0[0|0]/a_1197_107# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.25514f $ **FLOATING
C582 sky130_fd_sc_hvl__lsbuflv2hv_1_0[0|0]/a_1711_885# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.339894f $ **FLOATING
C583 sky130_fd_sc_hvl__lsbuflv2hv_1_0[0|0]/a_504_1221# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.834376f $ **FLOATING
C584 sky130_fd_sc_hvl__lsbuflv2hv_1_0[0|0]/a_404_1133# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 1.44294f $ **FLOATING
C585 schmitt_trigger_0/out sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.809398f
C586 schmitt_trigger_0/m sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 1.563827f
C587 schmitt_trigger_0/in sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 21.047577f
C588 por_unbuf sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 1.262839f
C589 sky130_fd_sc_hd__inv_4_1/Y sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.556998f
C590 sky130_fd_sc_hd__inv_4_2/Y sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.139892f
C591 sky130_fd_sc_hd__inv_4_0/Y sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.541678f
C592 sky130_fd_sc_hvl__inv_4_0/A sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 1.167166f
C593 rstring_mux_0/m1_26606_n3340# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 1.004901f
C594 rstring_mux_0/m1_26228_4059# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.864185f
C595 rstring_mux_0/m1_25850_n3340# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.863782f
C596 rstring_mux_0/m1_25472_4059# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.864185f
C597 rstring_mux_0/m1_25094_n3340# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.863782f
C598 rstring_mux_0/m1_24716_4059# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.864185f
C599 rstring_mux_0/m1_24338_n3340# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.863782f
C600 rstring_mux_0/m1_23960_4059# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.864185f
C601 rstring_mux_0/m1_23582_n3340# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.863782f
C602 rstring_mux_0/m1_23204_4059# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.864185f
C603 rstring_mux_0/m1_22826_n3340# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.863782f
C604 rstring_mux_0/m1_22448_4059# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.864185f
C605 rstring_mux_0/m1_22070_n3340# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.863782f
C606 rstring_mux_0/m1_21692_4059# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.864185f
C607 rstring_mux_0/m1_21314_n3340# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.863782f
C608 rstring_mux_0/m1_20936_4059# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.864185f
C609 rstring_mux_0/m1_20558_n3340# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.863782f
C610 rstring_mux_0/m1_20180_4059# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.864185f
C611 rstring_mux_0/m1_19802_n3340# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.863782f
C612 rstring_mux_0/m1_19424_4059# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.864185f
C613 rstring_mux_0/m1_19046_n3340# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.863782f
C614 rstring_mux_0/m1_18668_4059# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.864185f
C615 rstring_mux_0/m1_18290_n3340# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.863782f
C616 rstring_mux_0/m1_17912_4059# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.864185f
C617 rstring_mux_0/m1_17534_n3340# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.863782f
C618 rstring_mux_0/m1_17156_4059# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.864185f
C619 rstring_mux_0/m1_16778_n3340# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.863782f
C620 rstring_mux_0/vtrip7 sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 2.66344f
C621 rstring_mux_0/vtrip6 sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 3.339098f
C622 rstring_mux_0/vtrip5 sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 1.646662f
C623 rstring_mux_0/vtrip4 sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 2.752712f
C624 rstring_mux_0/vtrip3 sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 1.848688f
C625 rstring_mux_0/vtrip2 sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 2.952543f
C626 rstring_mux_0/vtrip1 sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 1.659759f
C627 rstring_mux_0/vtrip0 sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 3.67242f
C628 rstring_mux_0/m1_13376_4059# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.864185f
C629 rstring_mux_0/m1_12998_n3340# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.863782f
C630 rstring_mux_0/m1_12620_4059# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.864449f
C631 rstring_mux_0/m1_12242_n3340# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.863782f
C632 rstring_mux_0/m1_11864_4059# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.874226f
C633 rstring_mux_0/m1_11486_n3340# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.863782f
C634 rstring_mux_0/m1_11108_4059# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.864185f
C635 rstring_mux_0/m1_10730_n3340# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.863782f
C636 rstring_mux_0/m1_10352_4059# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.864185f
C637 rstring_mux_0/m1_9974_n3340# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.863782f
C638 rstring_mux_0/m1_9596_4059# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.864185f
C639 rstring_mux_0/m1_9218_n3340# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.863782f
C640 rstring_mux_0/m1_8840_4059# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.864185f
C641 rstring_mux_0/m1_8462_n3340# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.863782f
C642 rstring_mux_0/m1_8084_4059# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.864185f
C643 rstring_mux_0/m1_7706_n3340# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.863782f
C644 rstring_mux_0/m1_7328_4059# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.864185f
C645 rstring_mux_0/m1_6950_n3340# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.863782f
C646 rstring_mux_0/m1_6572_4059# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.864185f
C647 rstring_mux_0/m1_6194_n3340# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.863782f
C648 rstring_mux_0/m1_5816_4059# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.864185f
C649 rstring_mux_0/m1_5438_n3340# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.863782f
C650 rstring_mux_0/m1_5060_4059# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.864185f
C651 rstring_mux_0/m1_4682_n3340# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.863782f
C652 rstring_mux_0/m1_4304_4059# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.865582f
C653 rstring_mux_0/m1_3926_n3340# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.863782f
C654 rstring_mux_0/m1_3548_4059# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.865599f
C655 rstring_mux_0/m1_3170_n3340# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.863782f
C656 rstring_mux_0/m1_2792_4059# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.864381f
C657 rstring_mux_0/m1_2414_n3340# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.863782f
C658 rstring_mux_0/m1_2036_4059# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.864185f
C659 rstring_mux_0/m1_1658_n3340# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.863782f
C660 rstring_mux_0/m1_1280_4059# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.864185f
C661 rstring_mux_0/m1_902_n3340# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 1.005741f
C662 rstring_mux_0/vtop sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 5.554826f
C663 rstring_mux_0/ena_b sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 3.604659f
C664 rstring_mux_0/vtrip_decoded_b_avdd[7] sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.688611f
C665 rstring_mux_0/vtrip_decoded_b_avdd[6] sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.487044f
C666 rstring_mux_0/vtrip_decoded_b_avdd[5] sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.487044f
C667 rstring_mux_0/vtrip_decoded_b_avdd[4] sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.487044f
C668 rstring_mux_0/vtrip_decoded_b_avdd[3] sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.487035f
C669 rstring_mux_0/vtrip_decoded_b_avdd[2] sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.487041f
C670 rstring_mux_0/vtrip_decoded_b_avdd[1] sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.487044f
C671 rstring_mux_0/vtrip_decoded_b_avdd[0] sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.487044f
C672 rstring_mux_0/otrip_decoded_b_avdd[7] sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.487044f
C673 rstring_mux_0/otrip_decoded_b_avdd[6] sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.487034f
C674 rstring_mux_0/otrip_decoded_b_avdd[5] sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.487044f
C675 rstring_mux_0/otrip_decoded_b_avdd[4] sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.487044f
C676 rstring_mux_0/otrip_decoded_b_avdd[3] sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.487041f
C677 rstring_mux_0/otrip_decoded_b_avdd[2] sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.487041f
C678 rstring_mux_0/otrip_decoded_b_avdd[1] sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.487025f
C679 rstring_mux_0/otrip_decoded_b_avdd[0] sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.50765f
C680 comparator_0/vinn sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 31.27614f
C681 rstring_mux_0/vtrip_decoded_avdd[7] sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 2.111897f
C682 rstring_mux_0/vtrip_decoded_avdd[6] sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 1.97831f
C683 rstring_mux_0/vtrip_decoded_avdd[5] sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 2.103795f
C684 rstring_mux_0/vtrip_decoded_avdd[4] sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 1.967166f
C685 rstring_mux_0/vtrip_decoded_avdd[3] sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 2.090342f
C686 rstring_mux_0/vtrip_decoded_avdd[2] sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 1.925149f
C687 rstring_mux_0/vtrip_decoded_avdd[1] sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 2.034503f
C688 rstring_mux_0/vtrip_decoded_avdd[0] sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 1.976057f
C689 rstring_mux_0/otrip_decoded_avdd[7] sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 2.05949f
C690 rstring_mux_0/otrip_decoded_avdd[6] sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 1.890064f
C691 rstring_mux_0/otrip_decoded_avdd[5] sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 1.914958f
C692 rstring_mux_0/otrip_decoded_avdd[4] sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 1.743749f
C693 rstring_mux_0/otrip_decoded_avdd[3] sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 1.703108f
C694 rstring_mux_0/otrip_decoded_avdd[2] sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 2.020533f
C695 rstring_mux_0/otrip_decoded_avdd[1] sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 1.991324f
C696 rstring_mux_0/otrip_decoded_avdd[0] sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 1.991109f
C697 sky130_fd_sc_hvl__lsbufhv2lv_1_1/X sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.300918f
C698 sky130_fd_sc_hvl__lsbufhv2lv_1_1/a_30_207# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.665049f $ **FLOATING
C699 sky130_fd_sc_hvl__lsbufhv2lv_1_1/a_389_141# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.635783f $ **FLOATING
C700 sky130_fd_sc_hvl__lsbufhv2lv_1_1/a_389_1337# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.510776f $ **FLOATING
C701 sky130_fd_sc_hvl__lsbufhv2lv_1_1/a_30_1337# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 1.03613f $ **FLOATING
C702 vl sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 3.372648f
C703 sky130_fd_sc_hvl__lsbufhv2lv_1_0/a_30_207# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.665049f $ **FLOATING
C704 sky130_fd_sc_hvl__lsbufhv2lv_1_0/a_389_141# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.635783f $ **FLOATING
C705 sky130_fd_sc_hvl__lsbufhv2lv_1_0/a_389_1337# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 0.510776f $ **FLOATING
C706 sky130_fd_sc_hvl__lsbufhv2lv_1_0/a_30_1337# sky130_fd_pr__cap_mim_m3_2_LUWKLG_0/0 1.03613f $ **FLOATING
.ends

