magic
tech sky130A
magscale 1 2
timestamp 1713454396
<< error_s >>
rect 39827 23173 39828 23227
rect 39887 23123 39888 23173
rect 39887 22853 39888 22937
<< pwell >>
rect -1182 40391 42901 40527
rect -1182 -559 -1046 40391
rect 42765 -559 42901 40391
rect -1182 -695 42901 -559
<< psubdiff >>
rect -1146 40457 -1086 40491
rect 42805 40457 42865 40491
rect -1146 40431 -1112 40457
rect 42831 40431 42865 40457
rect 2221 27119 14128 27167
rect 2221 27058 2342 27119
rect 14001 27058 14128 27119
rect 2221 27022 14128 27058
rect 1136 1958 12732 1994
rect 1136 1899 1234 1958
rect 12612 1899 12732 1958
rect 1136 1857 12732 1899
rect -1146 -625 -1112 -599
rect 42831 -625 42865 -599
rect -1146 -659 -1086 -625
rect 42805 -659 42865 -625
<< psubdiffcont >>
rect -1086 40457 42805 40491
rect -1146 -599 -1112 40431
rect 2342 27058 14001 27119
rect 1234 1899 12612 1958
rect 42831 -599 42865 40431
rect -1086 -659 42805 -625
<< locali >>
rect -1146 40457 -1086 40491
rect 42805 40457 42865 40491
rect -1146 40431 -1112 40457
rect 42831 40431 42865 40457
rect -1146 -625 -1112 -599
rect 42831 -625 42865 -599
rect -1146 -659 -1086 -625
rect 42805 -659 42865 -625
<< viali >>
rect -1086 40457 42805 40491
rect -1146 -556 -1112 40404
rect 30169 38779 30234 38813
rect -704 32356 -670 32407
rect 2284 27058 2342 27119
rect 2342 27058 14001 27119
rect 14001 27058 14069 27119
rect 42460 26481 42494 26531
rect 1191 1899 1234 1958
rect 1234 1899 12612 1958
rect 12612 1899 12675 1958
rect 42831 -567 42865 40393
rect -1086 -659 42805 -625
<< metal1 >>
rect 41177 40531 41325 40612
rect -1186 40491 42905 40531
rect -1186 40457 -1086 40491
rect 42805 40457 42905 40491
rect -1186 40404 42905 40457
rect -1186 -556 -1146 40404
rect -1112 40393 42905 40404
rect -1112 40391 42831 40393
rect -1112 32422 -1046 40391
rect 30161 38813 30242 40391
rect 30161 38779 30169 38813
rect 30234 38779 30242 38813
rect 30161 38681 30242 38779
rect 29714 38635 31024 38681
rect 29714 38603 29760 38635
rect 30030 38603 30076 38635
rect 30346 38603 30392 38635
rect 30662 38603 30708 38635
rect 30978 38602 31024 38635
rect 29854 38541 29918 38547
rect 29854 38489 29860 38541
rect 29912 38489 29918 38541
rect 30808 38539 30872 38545
rect 29854 38483 29918 38489
rect 30171 38526 30235 38532
rect 30171 38474 30177 38526
rect 30229 38474 30235 38526
rect 30171 38468 30235 38474
rect 30483 38527 30547 38533
rect 30483 38475 30489 38527
rect 30541 38475 30547 38527
rect 30808 38487 30814 38539
rect 30866 38487 30872 38539
rect 30808 38481 30872 38487
rect 30483 38469 30547 38475
rect -433 32570 -361 32576
rect -433 32510 -427 32570
rect -367 32510 -361 32570
rect -433 32504 -361 32510
rect -576 32422 -530 32423
rect -1112 32407 -530 32422
rect -1112 32356 -704 32407
rect -670 32388 -530 32407
rect -260 32388 -214 32422
rect -670 32356 -214 32388
rect -1112 32342 -214 32356
rect -1112 -556 -1046 32342
rect 42284 27618 42362 27664
rect 42316 27608 42362 27618
rect 42118 27510 42182 27516
rect 42118 27458 42124 27510
rect 42176 27458 42182 27510
rect 42118 27452 42182 27458
rect 42316 27348 42362 27516
rect 42284 27302 42362 27348
rect 42180 27196 42244 27202
rect 2221 27119 14128 27167
rect 42180 27144 42186 27196
rect 42238 27144 42244 27196
rect 42180 27138 42244 27144
rect 2221 27118 2284 27119
rect 1695 27055 1701 27118
rect 1764 27058 2284 27118
rect 14069 27058 14128 27119
rect 1764 27055 14128 27058
rect 2221 27022 14128 27055
rect 42316 27032 42362 27302
rect 42284 26986 42362 27032
rect 42112 26882 42176 26888
rect 42112 26830 42118 26882
rect 42170 26830 42176 26882
rect 42112 26824 42176 26830
rect 42316 26716 42362 26986
rect 42284 26670 42362 26716
rect 42099 26566 42163 26572
rect 42099 26514 42105 26566
rect 42157 26514 42163 26566
rect 42099 26508 42163 26514
rect 42316 26543 42362 26670
rect 42765 26543 42831 40391
rect 42316 26531 42831 26543
rect 42316 26481 42460 26531
rect 42494 26481 42831 26531
rect 42316 26473 42831 26481
rect 42316 26400 42362 26473
rect 42284 26354 42362 26400
rect 42092 26256 42156 26262
rect 42092 26204 42098 26256
rect 42150 26204 42156 26256
rect 42092 26198 42156 26204
rect 42316 26186 42362 26354
rect 42316 26084 42362 26094
rect 42284 26038 42362 26084
rect 42765 25388 42831 26473
rect 42764 25281 42831 25388
rect 41034 24175 41174 24425
rect 41424 24175 41430 24425
rect 41158 24106 41256 24147
rect 41158 24091 41475 24106
rect 41256 24049 41475 24091
rect 41158 23987 41256 23993
rect 41078 23255 41084 23611
rect 41440 23255 41446 23611
rect 41020 22441 41224 22691
rect 41474 22441 41480 22691
rect 41193 22357 41716 22413
rect 41193 22313 41616 22357
rect 41616 22251 41716 22257
rect 41039 21567 41045 21877
rect 41355 21567 41361 21877
rect 39545 21372 40782 21511
rect 39545 21311 41108 21372
rect 39492 21055 40301 21255
rect 40582 21172 41108 21311
rect 41308 21172 41314 21372
rect 40101 21003 40301 21055
rect 40101 20803 41078 21003
rect 41278 20803 41284 21003
rect 34014 14819 34488 15019
rect 34688 14819 34694 15019
rect 6844 1994 6850 2004
rect 1136 1958 6850 1994
rect 6988 1994 6994 2004
rect 6988 1958 12732 1994
rect 1136 1899 1191 1958
rect 12675 1899 12732 1958
rect 1136 1866 6850 1899
rect 6988 1866 12732 1899
rect 1136 1857 12732 1866
rect 42252 127 42348 133
rect 42252 25 42348 31
rect -1186 -559 -1046 -556
rect 42765 -559 42831 25281
rect -1186 -567 42831 -559
rect 42865 -567 42905 40393
rect -1186 -625 42905 -567
rect -1186 -659 -1086 -625
rect 42805 -659 42905 -625
rect -1186 -699 42905 -659
<< via1 >>
rect 29860 38489 29912 38541
rect 30177 38474 30229 38526
rect 30489 38475 30541 38527
rect 30814 38487 30866 38539
rect -427 32510 -367 32570
rect 42124 27458 42176 27510
rect 42186 27144 42238 27196
rect 1701 27055 1764 27118
rect 42118 26830 42170 26882
rect 42105 26514 42157 26566
rect 42098 26204 42150 26256
rect 41266 24989 41414 25137
rect 41174 24175 41424 24425
rect 41158 23993 41256 24091
rect 41084 23255 41440 23611
rect 41224 22441 41474 22691
rect 41616 22257 41716 22357
rect 41045 21567 41355 21877
rect 41108 21172 41308 21372
rect 41078 20803 41278 21003
rect 34488 14819 34688 15019
rect 6850 1958 6988 2004
rect 6850 1899 6988 1958
rect 6850 1866 6988 1899
rect 42252 31 42348 127
<< metal2 >>
rect 1111 40272 1507 40292
rect 1111 39982 1131 40272
rect 1471 39982 1507 40272
rect 1111 39265 1507 39982
rect 1577 39865 1962 39896
rect 1577 39606 1599 39865
rect 1934 39606 1962 39865
rect 1577 39251 1962 39606
rect 10871 38396 10935 41282
rect 10858 38387 10935 38396
rect 10914 38331 10935 38387
rect 10858 38322 10935 38331
rect 10871 32731 10935 38322
rect 10871 32667 11144 32731
rect -425 32576 -369 32577
rect -433 32570 -361 32576
rect -433 32510 -427 32570
rect -367 32510 -361 32570
rect -433 32504 -361 32510
rect -425 32503 -369 32504
rect 11080 32217 11144 32667
rect 1701 27118 1764 27124
rect 1701 27049 1764 27055
rect 11841 26826 11850 26892
rect 11916 26826 11925 26892
rect 12255 26887 12321 41282
rect 12255 26831 12260 26887
rect 12316 26831 12321 26887
rect 12255 26826 12321 26831
rect 11850 26541 11916 26826
rect 12260 26822 12316 26826
rect 14078 23704 14142 23713
rect 14956 23700 15020 41282
rect 21267 37305 21331 41282
rect 24466 41110 24594 41119
rect 24057 40197 24185 40206
rect 19650 35406 19710 35408
rect 19643 35350 19652 35406
rect 19708 35350 19717 35406
rect 14956 23644 14960 23700
rect 15016 23644 15020 23700
rect 14956 23640 15020 23644
rect 14078 23631 14142 23640
rect 14960 23635 15016 23640
rect 15263 4251 15319 4258
rect 15261 4249 15321 4251
rect 15261 4193 15263 4249
rect 15319 4193 15321 4249
rect 15261 3490 15321 4193
rect 19650 3696 19710 35350
rect 24057 33041 24185 40069
rect 24466 32861 24594 40982
rect 24666 40637 24794 40646
rect 24666 33742 24794 40509
rect 25575 37439 25631 37446
rect 25573 37437 25633 37439
rect 25573 37381 25575 37437
rect 25631 37381 25633 37437
rect 25573 32795 25633 37381
rect 26348 30339 26414 41282
rect 26775 30842 26841 41282
rect 27432 33447 27496 41282
rect 28854 36088 28914 41282
rect 28854 35411 28914 36028
rect 28847 35406 28921 35411
rect 28847 35350 28856 35406
rect 28912 35350 28921 35406
rect 28847 35341 28921 35350
rect 27235 33383 27496 33447
rect 26348 30283 26353 30339
rect 26409 30283 26414 30339
rect 26348 30278 26414 30283
rect 26766 30278 26775 30344
rect 26841 30278 26850 30344
rect 26353 30274 26409 30278
rect 26775 29996 26841 30278
rect 26795 27891 26851 27900
rect 26795 27826 26851 27835
rect 21332 27605 21388 27612
rect 21330 27603 21390 27605
rect 21330 27547 21332 27603
rect 21388 27547 21390 27603
rect 21147 26295 21203 26302
rect 21145 26293 21205 26295
rect 21145 26237 21147 26293
rect 21203 26237 21205 26293
rect 19899 26133 19959 26142
rect 19899 4249 19959 26073
rect 21145 22193 21205 26237
rect 21330 23778 21390 27547
rect 23589 27323 23645 27330
rect 23587 27321 23647 27323
rect 23587 27265 23589 27321
rect 23645 27265 23647 27321
rect 23128 26451 23184 26458
rect 23126 26449 23186 26451
rect 23126 26393 23128 26449
rect 23184 26393 23186 26449
rect 23126 23796 23186 26393
rect 23126 23736 23490 23796
rect 23587 22311 23647 27265
rect 27235 27077 27299 33383
rect 29342 32686 29402 41282
rect 29921 39211 29981 41282
rect 30421 39463 30481 41282
rect 30421 39403 30724 39463
rect 29921 39155 29923 39211
rect 29979 39155 29981 39211
rect 29921 39153 29981 39155
rect 30471 39153 30480 39213
rect 30540 39153 30549 39213
rect 29923 39146 29979 39153
rect 30178 38758 30234 38765
rect 30176 38756 30236 38758
rect 30176 38700 30178 38756
rect 30234 38700 30236 38756
rect 29854 38541 29918 38547
rect 29854 38489 29860 38541
rect 29912 38489 29918 38541
rect 30176 38532 30236 38700
rect 29854 38483 29918 38489
rect 30171 38526 30236 38532
rect 29857 38389 29913 38483
rect 30171 38474 30177 38526
rect 30229 38475 30236 38526
rect 30480 38533 30540 39153
rect 30664 38758 30724 39403
rect 30480 38527 30547 38533
rect 30480 38475 30489 38527
rect 30541 38475 30547 38527
rect 30229 38474 30235 38475
rect 30171 38468 30235 38474
rect 30480 38469 30547 38475
rect 29846 38329 29855 38389
rect 29915 38329 29924 38389
rect 30250 37754 30306 37761
rect 30248 37752 30308 37754
rect 30248 37696 30250 37752
rect 30306 37696 30308 37752
rect 30248 34036 30308 37696
rect 30248 33967 30308 33976
rect 29342 32630 29344 32686
rect 29400 32630 29402 32686
rect 29342 32628 29402 32630
rect 29344 32621 29400 32628
rect 30480 32190 30540 38469
rect 30664 33374 30724 38698
rect 30879 38545 30939 41282
rect 30808 38539 30939 38545
rect 30808 38487 30814 38539
rect 30866 38487 30939 38539
rect 30808 38481 30939 38487
rect 30664 33305 30724 33314
rect 30354 32130 30540 32190
rect 30354 31322 30414 32130
rect 30354 31253 30414 31262
rect 30481 32014 30541 32023
rect 30336 30640 30396 30649
rect 30336 27893 30396 30580
rect 30336 27824 30396 27833
rect 25406 27025 25462 27032
rect 25404 27023 25464 27025
rect 25404 26967 25406 27023
rect 25462 26967 25464 27023
rect 25404 23416 25464 26967
rect 27864 26893 27920 26900
rect 27862 26891 27922 26893
rect 27862 26835 27864 26891
rect 27920 26835 27922 26891
rect 25564 26752 25620 26759
rect 25562 26750 25622 26752
rect 25562 26694 25564 26750
rect 25620 26694 25622 26750
rect 25562 23807 25622 26694
rect 27653 26590 27709 26597
rect 27651 26588 27711 26590
rect 27651 26532 27653 26588
rect 27709 26532 27711 26588
rect 27651 23763 27711 26532
rect 25404 23356 25603 23416
rect 23436 22251 23647 22311
rect 21145 22133 21389 22193
rect 23436 22068 23496 22251
rect 25543 22062 25603 23356
rect 27862 22350 27922 26835
rect 30481 26131 30541 31954
rect 30481 26075 30483 26131
rect 30539 26075 30541 26131
rect 30481 26073 30541 26075
rect 30662 29960 30722 29969
rect 30662 26124 30722 29900
rect 30879 29228 30939 38481
rect 40594 37754 40654 37763
rect 35756 37439 35834 37448
rect 35756 37379 35765 37439
rect 35825 37379 35834 37439
rect 35756 37370 35834 37379
rect 40594 33372 40654 37694
rect 40586 33366 40662 33372
rect 40586 33310 40596 33366
rect 40652 33310 40662 33366
rect 40586 33300 40662 33310
rect 41322 32008 41378 32015
rect 41320 32006 41380 32008
rect 41320 31950 41322 32006
rect 41378 31950 41380 32006
rect 41320 31324 41380 31950
rect 41899 32006 41973 32015
rect 41899 31950 41908 32006
rect 41964 31950 41973 32006
rect 41899 31945 41973 31950
rect 41320 31255 41380 31264
rect 33836 27603 33892 27612
rect 33836 27538 33892 27547
rect 39066 27467 39122 27476
rect 39066 27402 39122 27411
rect 35214 27321 35270 27330
rect 35214 27256 35270 27265
rect 33186 27152 33242 27161
rect 33186 27087 33242 27096
rect 41372 27073 41428 27080
rect 41370 27071 41430 27073
rect 34474 27023 34530 27032
rect 34474 26958 34530 26967
rect 41370 27015 41372 27071
rect 41428 27015 41430 27071
rect 38340 26891 38396 26900
rect 38340 26826 38396 26835
rect 37696 26750 37752 26759
rect 37696 26685 37752 26694
rect 35766 26588 35822 26597
rect 37713 26544 37741 26674
rect 35766 26523 35822 26532
rect 37054 26449 37110 26458
rect 37054 26384 37110 26393
rect 38357 26326 38385 26677
rect 36418 26293 36474 26302
rect 36418 26228 36474 26237
rect 38073 26126 38129 26133
rect 30483 26066 30539 26073
rect 30662 26068 30664 26124
rect 30720 26068 30722 26124
rect 30662 26066 30722 26068
rect 38071 26124 38131 26126
rect 38071 26068 38073 26124
rect 38129 26068 38131 26124
rect 30664 26059 30720 26066
rect 32548 25966 32604 25975
rect 32548 25901 32604 25910
rect 27666 22290 27922 22350
rect 27666 22067 27726 22290
rect 38071 22163 38131 26068
rect 41370 25968 41430 27015
rect 41906 26567 41966 31945
rect 42110 27460 42119 27516
rect 42175 27510 42184 27516
rect 42176 27460 42184 27510
rect 42118 27458 42124 27460
rect 42176 27458 42182 27460
rect 42118 27452 42182 27458
rect 42179 27202 42239 27204
rect 42179 27196 42244 27202
rect 42179 27144 42186 27196
rect 42238 27144 42244 27196
rect 42179 27138 42244 27144
rect 42179 27071 42239 27138
rect 42179 27015 42181 27071
rect 42237 27015 42239 27071
rect 42179 27013 42239 27015
rect 42181 27006 42237 27013
rect 42112 26888 42172 26890
rect 42112 26882 42176 26888
rect 42112 26830 42118 26882
rect 42170 26830 42176 26882
rect 42112 26824 42176 26830
rect 42112 26732 42172 26824
rect 42112 26676 42114 26732
rect 42170 26676 42172 26732
rect 42112 26674 42172 26676
rect 42114 26667 42170 26674
rect 42104 26572 42160 26574
rect 42099 26566 42163 26572
rect 42099 26565 42105 26566
rect 42157 26565 42163 26566
rect 42099 26509 42104 26565
rect 42160 26509 42163 26565
rect 42099 26508 42163 26509
rect 41906 26498 41966 26507
rect 42104 26500 42160 26508
rect 42093 26262 42157 26272
rect 42092 26256 42157 26262
rect 42092 26204 42098 26256
rect 42150 26204 42157 26256
rect 42092 26198 42157 26204
rect 41370 25899 41430 25908
rect 41257 25137 41423 25146
rect 41257 24989 41266 25137
rect 41414 24989 41423 25137
rect 41257 24980 41423 24989
rect 41165 24425 41433 24434
rect 41165 24175 41174 24425
rect 41424 24175 41433 24425
rect 41165 24166 41433 24175
rect 41149 24091 41265 24100
rect 41149 23993 41158 24091
rect 41256 23993 41265 24091
rect 41149 23984 41265 23993
rect 38223 23859 38286 23861
rect 42093 23860 42157 26198
rect 38223 23732 38286 23795
rect 42088 23855 42162 23860
rect 42088 23799 42097 23855
rect 42153 23799 42162 23855
rect 42088 23790 42162 23799
rect 41075 23611 41449 23620
rect 41075 23255 41084 23611
rect 41440 23255 41449 23611
rect 41075 23246 41449 23255
rect 41215 22691 41483 22700
rect 41215 22441 41224 22691
rect 41474 22441 41483 22691
rect 41215 22432 41483 22441
rect 41606 22357 41725 22366
rect 41606 22257 41616 22357
rect 41716 22257 41725 22357
rect 41606 22248 41725 22257
rect 38071 22103 38286 22163
rect 41036 21877 41364 21886
rect 41036 21567 41045 21877
rect 41355 21567 41364 21877
rect 41036 21558 41364 21567
rect 19899 4193 19901 4249
rect 19957 4193 19959 4249
rect 19899 4191 19959 4193
rect 19901 4184 19957 4191
rect 19650 3627 19710 3636
rect 15159 3430 15321 3490
rect 6850 2004 6988 2010
rect 10 -707 396 1690
rect 493 -110 893 1899
rect 493 -519 893 -510
rect 6850 1731 6988 1866
rect 6850 -379 6985 1731
rect 6850 -523 6985 -514
rect 10 -1039 28 -707
rect 383 -1039 396 -707
rect 10 -1056 396 -1039
rect 20121 -1717 20249 4106
rect 20321 -855 20449 21377
rect 41098 21372 41318 21381
rect 41098 21172 41108 21372
rect 41308 21172 41318 21372
rect 41098 21161 41318 21172
rect 41068 21003 41288 21012
rect 41068 20803 41078 21003
rect 41278 20803 41288 21003
rect 41068 20792 41288 20803
rect 34478 15019 34698 15029
rect 34478 14819 34488 15019
rect 34688 14819 34698 15019
rect 34478 14809 34698 14819
rect 41883 4260 41892 4404
rect 42036 4260 42310 4404
rect 20321 -992 20449 -983
rect 20521 -1286 20649 3055
rect 42246 31 42252 127
rect 42348 31 42960 127
rect 43056 31 43065 127
rect 20521 -1423 20649 -1414
rect 20121 -1854 20249 -1845
<< via2 >>
rect 1131 39982 1471 40272
rect 1599 39606 1934 39865
rect 10858 38331 10914 38387
rect -425 32512 -369 32568
rect 11850 26826 11916 26892
rect 12260 26831 12316 26887
rect 14078 23640 14142 23704
rect 24466 40982 24594 41110
rect 24057 40069 24185 40197
rect 19652 35350 19708 35406
rect 14960 23644 15016 23700
rect 15263 4193 15319 4249
rect 24666 40509 24794 40637
rect 25575 37381 25631 37437
rect 28854 36028 28914 36088
rect 28856 35350 28912 35406
rect 26353 30283 26409 30339
rect 26775 30278 26841 30344
rect 26795 27835 26851 27891
rect 21332 27547 21388 27603
rect 21147 26237 21203 26293
rect 19899 26073 19959 26133
rect 23589 27265 23645 27321
rect 23128 26393 23184 26449
rect 29923 39155 29979 39211
rect 30480 39153 30540 39213
rect 30178 38700 30234 38756
rect 30664 38698 30724 38758
rect 29855 38329 29915 38389
rect 30250 37696 30306 37752
rect 30248 33976 30308 34036
rect 29344 32630 29400 32686
rect 30664 33314 30724 33374
rect 30354 31262 30414 31322
rect 30481 31954 30541 32014
rect 30336 30580 30396 30640
rect 30336 27833 30396 27893
rect 25406 26967 25462 27023
rect 27864 26835 27920 26891
rect 25564 26694 25620 26750
rect 27653 26532 27709 26588
rect 30483 26075 30539 26131
rect 30662 29900 30722 29960
rect 40594 37694 40654 37754
rect 35765 37379 35825 37439
rect 40596 33310 40652 33366
rect 41322 31950 41378 32006
rect 41908 31950 41964 32006
rect 41320 31264 41380 31324
rect 33836 27547 33892 27603
rect 39066 27411 39122 27467
rect 35214 27265 35270 27321
rect 33186 27096 33242 27152
rect 34474 26967 34530 27023
rect 41372 27015 41428 27071
rect 38340 26835 38396 26891
rect 37696 26694 37752 26750
rect 35766 26532 35822 26588
rect 37054 26393 37110 26449
rect 36418 26237 36474 26293
rect 30664 26068 30720 26124
rect 38073 26068 38129 26124
rect 32548 25910 32604 25966
rect 42119 27510 42175 27516
rect 42119 27460 42124 27510
rect 42124 27460 42175 27510
rect 42181 27015 42237 27071
rect 42114 26676 42170 26732
rect 41906 26507 41966 26567
rect 42104 26514 42105 26565
rect 42105 26514 42157 26565
rect 42157 26514 42160 26565
rect 42104 26509 42160 26514
rect 41370 25908 41430 25968
rect 41266 24989 41414 25137
rect 41174 24175 41424 24425
rect 41158 23993 41256 24091
rect 38222 23795 38286 23859
rect 42097 23799 42153 23855
rect 41084 23255 41440 23611
rect 41224 22441 41474 22691
rect 41616 22257 41716 22357
rect 41045 21567 41355 21877
rect 19901 4193 19957 4249
rect 19650 3636 19710 3696
rect 493 -510 893 -110
rect 6850 -514 6985 -379
rect 28 -1039 383 -707
rect 41108 21172 41308 21372
rect 41078 20803 41278 21003
rect 34488 14819 34688 15019
rect 41892 4260 42036 4404
rect 20321 -983 20449 -855
rect 42960 31 43056 127
rect 20521 -1414 20649 -1286
rect 20121 -1845 20249 -1717
<< metal3 >>
rect -1604 41276 43293 41282
rect -1604 40888 -1598 41276
rect -1210 41248 42899 41276
rect -1210 41110 34162 41248
rect -1210 40982 24466 41110
rect 24594 40982 34162 41110
rect -1210 40930 34162 40982
rect 34480 40930 42899 41248
rect -1210 40888 42899 40930
rect 43287 40888 43293 41276
rect -1604 40882 43293 40888
rect -1604 40816 43293 40822
rect -1604 40428 -1138 40816
rect -750 40772 42439 40816
rect -750 40637 34822 40772
rect -750 40509 24666 40637
rect 24794 40509 34822 40637
rect -750 40454 34822 40509
rect 35140 40454 42439 40772
rect -750 40428 42439 40454
rect 42827 40428 43293 40816
rect -1604 40422 43293 40428
rect -1604 40356 43293 40362
rect -1604 39968 -678 40356
rect -290 40272 41979 40356
rect -290 39982 1131 40272
rect 1471 40197 41979 40272
rect 1471 40069 24057 40197
rect 24185 40069 41979 40197
rect 1471 39982 41979 40069
rect -290 39968 41979 39982
rect 42367 39968 43293 40356
rect -1604 39962 43293 39968
rect -1604 39896 43293 39902
rect -1604 39508 -218 39896
rect 170 39865 41519 39896
rect 170 39606 1599 39865
rect 1934 39606 41519 39865
rect 170 39508 41519 39606
rect 41907 39508 43293 39896
rect -1604 39502 43293 39508
rect 947 39492 1357 39502
rect 29918 39213 29984 39216
rect 30475 39213 30545 39218
rect 29918 39211 30480 39213
rect 29918 39155 29923 39211
rect 29979 39155 30480 39211
rect 29918 39153 30480 39155
rect 30540 39153 30545 39213
rect 29918 39150 29984 39153
rect 30475 39148 30545 39153
rect 30173 38758 30239 38761
rect 30659 38758 30729 38763
rect 30173 38756 30664 38758
rect 30173 38700 30178 38756
rect 30234 38700 30664 38756
rect 30173 38698 30664 38700
rect 30724 38698 30729 38758
rect 30173 38695 30239 38698
rect 30659 38693 30729 38698
rect 10853 38389 10919 38392
rect 29850 38389 29920 38394
rect 10853 38387 29855 38389
rect 10853 38331 10858 38387
rect 10914 38331 29855 38387
rect 10853 38329 29855 38331
rect 29915 38329 29920 38389
rect 10853 38326 10919 38329
rect 29850 38324 29920 38329
rect 30245 37754 30311 37757
rect 40589 37754 40659 37759
rect 30245 37752 40594 37754
rect 30245 37696 30250 37752
rect 30306 37696 40594 37752
rect 30245 37694 40594 37696
rect 40654 37694 40659 37754
rect 30245 37691 30311 37694
rect 40589 37689 40659 37694
rect 25570 37439 25636 37442
rect 35760 37439 35830 37444
rect 25570 37437 35765 37439
rect 25570 37381 25575 37437
rect 25631 37381 35765 37437
rect 25570 37379 35765 37381
rect 35825 37379 35830 37439
rect 25570 37376 25636 37379
rect 35760 37374 35830 37379
rect 28849 36088 28919 36093
rect 28849 36028 28854 36088
rect 28914 36028 30082 36088
rect 28849 36023 28919 36028
rect 19647 35408 19713 35411
rect 28851 35408 28917 35411
rect 19647 35406 28922 35408
rect 19647 35350 19652 35406
rect 19708 35350 28856 35406
rect 28912 35350 28922 35406
rect 19647 35348 28922 35350
rect 19647 35345 19713 35348
rect 28851 35345 28917 35348
rect 30243 34036 30313 34041
rect 30243 33976 30248 34036
rect 30308 33976 30313 34036
rect 30243 33971 30313 33976
rect 30659 33374 30729 33379
rect 30659 33314 30664 33374
rect 30724 33314 30729 33374
rect 40591 33368 40657 33371
rect 30659 33309 30729 33314
rect 40579 33366 43293 33368
rect 40579 33310 40596 33366
rect 40652 33310 43293 33366
rect 40579 33308 43293 33310
rect 40591 33305 40657 33308
rect 29339 32688 29405 32691
rect 29339 32686 30842 32688
rect 29339 32630 29344 32686
rect 29400 32630 30842 32686
rect 29339 32628 30842 32630
rect 29339 32625 29405 32628
rect -430 32570 -364 32573
rect -1604 32568 4716 32570
rect -1604 32512 -425 32568
rect -369 32512 4716 32568
rect -1604 32510 4716 32512
rect -430 32507 -364 32510
rect 30476 32014 30546 32019
rect 30476 31954 30481 32014
rect 30541 31954 30546 32014
rect 30476 31949 30546 31954
rect 41317 32008 41383 32011
rect 41903 32008 41969 32011
rect 41317 32006 43293 32008
rect 41317 31950 41322 32006
rect 41378 31950 41908 32006
rect 41964 31950 43293 32006
rect 41317 31948 43293 31950
rect 41317 31945 41383 31948
rect 41903 31945 41969 31948
rect 30349 31322 30419 31327
rect 30349 31262 30354 31322
rect 30414 31262 30419 31322
rect 30349 31257 30419 31262
rect 41315 31324 41385 31329
rect 41315 31264 41320 31324
rect 41380 31264 41385 31324
rect 41315 31259 41385 31264
rect 30331 30640 30401 30645
rect 30331 30580 30336 30640
rect 30396 30580 30401 30640
rect 30331 30575 30401 30580
rect 26770 30344 26846 30349
rect 26348 30339 26775 30344
rect 26348 30283 26353 30339
rect 26409 30283 26775 30339
rect 26348 30278 26775 30283
rect 26841 30278 26846 30344
rect 26770 30273 26846 30278
rect 30657 29960 30727 29965
rect 30657 29900 30662 29960
rect 30722 29900 30727 29960
rect 30657 29895 30727 29900
rect 26790 27893 26856 27896
rect 30331 27893 30401 27898
rect 26790 27891 30336 27893
rect 26790 27835 26795 27891
rect 26851 27835 30336 27891
rect 26790 27833 30336 27835
rect 30396 27833 34089 27893
rect 26790 27830 26856 27833
rect 30331 27828 30401 27833
rect 34029 27797 34089 27833
rect 34029 27737 43293 27797
rect 21327 27605 21393 27608
rect 33831 27605 33897 27608
rect 21327 27603 33897 27605
rect 21327 27547 21332 27603
rect 21388 27547 33836 27603
rect 33892 27547 33897 27603
rect 21327 27545 33897 27547
rect 21327 27542 21393 27545
rect 33831 27542 33897 27545
rect 42114 27516 42180 27521
rect 39061 27469 39127 27472
rect 42114 27469 42119 27516
rect 39061 27467 42119 27469
rect 39061 27411 39066 27467
rect 39122 27460 42119 27467
rect 42175 27469 42180 27516
rect 42175 27460 43293 27469
rect 39122 27411 43293 27460
rect 39061 27409 43293 27411
rect 39061 27406 39127 27409
rect 23584 27323 23650 27326
rect 35209 27323 35275 27326
rect 23584 27321 35275 27323
rect 23584 27265 23589 27321
rect 23645 27265 35214 27321
rect 35270 27265 35275 27321
rect 23584 27263 35275 27265
rect 23584 27260 23650 27263
rect 35209 27260 35275 27263
rect 33181 27154 33247 27157
rect 33181 27152 41186 27154
rect 33181 27096 33186 27152
rect 33242 27096 41186 27152
rect 33181 27094 41186 27096
rect 33181 27091 33247 27094
rect 25401 27025 25467 27028
rect 34469 27025 34535 27028
rect 25401 27023 34535 27025
rect 25401 26967 25406 27023
rect 25462 26967 34474 27023
rect 34530 26967 34535 27023
rect 25401 26965 34535 26967
rect 25401 26962 25467 26965
rect 34469 26962 34535 26965
rect 11845 26892 11921 26897
rect 27859 26893 27925 26896
rect 38335 26893 38401 26896
rect 11845 26826 11850 26892
rect 11916 26887 12321 26892
rect 11916 26831 12260 26887
rect 12316 26831 12321 26887
rect 11916 26826 12321 26831
rect 27859 26891 38401 26893
rect 27859 26835 27864 26891
rect 27920 26835 38340 26891
rect 38396 26835 38401 26891
rect 27859 26833 38401 26835
rect 27859 26830 27925 26833
rect 38335 26830 38401 26833
rect 11845 26821 11921 26826
rect 25559 26752 25625 26755
rect 37691 26752 37757 26755
rect 25559 26750 37757 26752
rect 25559 26694 25564 26750
rect 25620 26694 37696 26750
rect 37752 26694 37757 26750
rect 25559 26692 37757 26694
rect 25559 26689 25625 26692
rect 37691 26689 37757 26692
rect 41126 26734 41186 27094
rect 41367 27073 41433 27076
rect 42176 27073 42242 27076
rect 41367 27071 43293 27073
rect 41367 27015 41372 27071
rect 41428 27015 42181 27071
rect 42237 27015 43293 27071
rect 41367 27013 43293 27015
rect 41367 27010 41433 27013
rect 42176 27010 42242 27013
rect 42109 26734 42175 26737
rect 41126 26732 43293 26734
rect 41126 26676 42114 26732
rect 42170 26676 43293 26732
rect 41126 26674 43293 26676
rect 42109 26671 42175 26674
rect 27648 26590 27714 26593
rect 35761 26590 35827 26593
rect 27648 26588 35827 26590
rect 27648 26532 27653 26588
rect 27709 26532 35766 26588
rect 35822 26532 35827 26588
rect 27648 26530 35827 26532
rect 27648 26527 27714 26530
rect 35761 26527 35827 26530
rect 41901 26567 41971 26572
rect 42099 26567 42165 26570
rect 41901 26507 41906 26567
rect 41966 26565 42165 26567
rect 41966 26509 42104 26565
rect 42160 26509 42165 26565
rect 41966 26507 42165 26509
rect 41901 26502 41971 26507
rect 42099 26504 42165 26507
rect 23123 26451 23189 26454
rect 37049 26451 37115 26454
rect 23123 26449 37115 26451
rect 23123 26393 23128 26449
rect 23184 26393 37054 26449
rect 37110 26393 37115 26449
rect 23123 26391 37115 26393
rect 23123 26388 23189 26391
rect 37049 26388 37115 26391
rect 21142 26295 21208 26298
rect 36413 26295 36479 26298
rect 21142 26293 36479 26295
rect 21142 26237 21147 26293
rect 21203 26237 36418 26293
rect 36474 26237 36479 26293
rect 21142 26235 36479 26237
rect 21142 26232 21208 26235
rect 36413 26232 36479 26235
rect 19894 26133 19964 26138
rect 30478 26133 30544 26136
rect 19894 26073 19899 26133
rect 19959 26131 30544 26133
rect 19959 26075 30483 26131
rect 30539 26075 30544 26131
rect 19959 26073 30544 26075
rect 19894 26068 19964 26073
rect 30478 26070 30544 26073
rect 30659 26126 30725 26129
rect 38068 26126 38134 26129
rect 30659 26124 38134 26126
rect 30659 26068 30664 26124
rect 30720 26068 38073 26124
rect 38129 26068 38134 26124
rect 30659 26066 38134 26068
rect 30659 26063 30725 26066
rect 38068 26063 38134 26066
rect 32543 25968 32609 25971
rect 41365 25968 41435 25973
rect 32543 25966 41370 25968
rect 32543 25910 32548 25966
rect 32604 25910 41370 25966
rect 32543 25908 41370 25910
rect 41430 25908 41435 25968
rect 32543 25905 32609 25908
rect 41365 25903 41435 25908
rect 34821 25712 42435 25713
rect 34816 25394 34822 25712
rect 35140 25394 42435 25712
rect 34821 25393 42435 25394
rect 42755 25393 42761 25713
rect 41261 25137 41419 25142
rect 41261 24989 41266 25137
rect 41414 24989 42463 25137
rect 42611 24989 42617 25137
rect 41261 24984 41419 24989
rect 34161 24835 42939 24836
rect 34156 24517 34162 24835
rect 34480 24517 42939 24835
rect 34161 24516 42939 24517
rect 43259 24516 43265 24836
rect 41169 24425 41429 24430
rect 41169 24175 41174 24425
rect 41424 24175 42057 24425
rect 42307 24175 42313 24425
rect 41169 24170 41429 24175
rect 41153 24091 41261 24096
rect 41153 23993 41158 24091
rect 41256 23993 42933 24091
rect 43031 23993 43037 24091
rect 41153 23988 41261 23993
rect 38217 23859 38291 23864
rect 42092 23859 42158 23860
rect 38217 23795 38222 23859
rect 38286 23855 43293 23859
rect 38286 23799 42097 23855
rect 42153 23799 43293 23855
rect 38286 23795 43293 23799
rect 38217 23790 38291 23795
rect 42092 23794 42158 23795
rect 14073 23704 14147 23709
rect 14955 23704 15021 23705
rect 14073 23640 14078 23704
rect 14142 23700 15021 23704
rect 14142 23644 14960 23700
rect 15016 23644 15021 23700
rect 14142 23640 15021 23644
rect 14073 23635 14147 23640
rect 14955 23639 15021 23640
rect 41079 23611 41445 23616
rect 41079 23255 41084 23611
rect 41440 23255 42470 23611
rect 42826 23255 42832 23611
rect 41079 23250 41445 23255
rect 41219 22691 41479 22696
rect 41219 22441 41224 22691
rect 41474 22441 42015 22691
rect 42265 22441 42271 22691
rect 41219 22436 41479 22441
rect 41611 22357 41721 22362
rect 41611 22257 41616 22357
rect 41716 22257 42988 22357
rect 43088 22257 43094 22357
rect 41611 22252 41721 22257
rect 41040 21877 41360 21882
rect 41040 21567 41045 21877
rect 41355 21567 42503 21877
rect 42813 21567 42819 21877
rect 41040 21562 41360 21567
rect 41103 21372 41313 21377
rect 41103 21172 41108 21372
rect 41308 21172 42943 21372
rect 43143 21172 43149 21372
rect 41103 21167 41313 21172
rect 41073 21003 41283 21008
rect 41073 20803 41078 21003
rect 41278 20803 42063 21003
rect 42263 20803 42269 21003
rect 41073 20798 41283 20803
rect 34483 15019 34693 15024
rect 34483 14819 34488 15019
rect 34688 14819 42088 15019
rect 42288 14819 42294 15019
rect 34483 14814 34693 14819
rect 39201 14569 41613 14717
rect 41761 14569 41767 14717
rect 41887 4404 42041 4409
rect 41887 4260 41892 4404
rect 42036 4260 42538 4404
rect 42682 4260 42688 4404
rect 41887 4255 42041 4260
rect 15258 4251 15324 4254
rect 19896 4251 19962 4254
rect 15258 4249 19962 4251
rect 15258 4193 15263 4249
rect 15319 4193 19901 4249
rect 19957 4193 19962 4249
rect 15258 4191 19962 4193
rect 15258 4188 15324 4191
rect 19896 4188 19962 4191
rect 19645 3696 19715 3701
rect 18622 3636 19650 3696
rect 19710 3636 19715 3696
rect 19645 3631 19715 3636
rect 42949 132 43067 138
rect 42949 26 42955 132
rect 43061 26 43067 132
rect 42949 20 43067 26
rect 488 -110 898 -105
rect 488 -207 493 -110
rect -1604 -213 493 -207
rect -1604 -601 -218 -213
rect 170 -510 493 -213
rect 893 -207 898 -110
rect 893 -213 43293 -207
rect 893 -379 41519 -213
rect 893 -510 6850 -379
rect 170 -514 6850 -510
rect 6985 -514 41519 -379
rect 170 -601 41519 -514
rect 41907 -601 43293 -213
rect -1604 -607 43293 -601
rect -1604 -673 43293 -667
rect -1604 -1061 -678 -673
rect -290 -707 41979 -673
rect -290 -1039 28 -707
rect 383 -855 41979 -707
rect 383 -983 20321 -855
rect 20449 -983 41979 -855
rect 383 -1039 41979 -983
rect -290 -1061 41979 -1039
rect 42367 -1061 43293 -673
rect -1604 -1067 43293 -1061
rect -1604 -1133 43293 -1127
rect -1604 -1521 -1138 -1133
rect -750 -1286 42439 -1133
rect -750 -1414 20521 -1286
rect 20649 -1414 42439 -1286
rect -750 -1521 42439 -1414
rect 42827 -1521 43293 -1133
rect -1604 -1527 43293 -1521
rect -1604 -1593 43293 -1587
rect -1604 -1981 -1598 -1593
rect -1210 -1717 42899 -1593
rect -1210 -1845 20121 -1717
rect 20249 -1845 42899 -1717
rect -1210 -1981 42899 -1845
rect 43287 -1981 43293 -1593
rect -1604 -1987 43293 -1981
<< via3 >>
rect -1598 40888 -1210 41276
rect 34162 40930 34480 41248
rect 42899 40888 43287 41276
rect -1138 40428 -750 40816
rect 34822 40454 35140 40772
rect 42439 40428 42827 40816
rect -678 39968 -290 40356
rect 41979 39968 42367 40356
rect -218 39508 170 39896
rect 41519 39508 41907 39896
rect 34822 25394 35140 25712
rect 42435 25393 42755 25713
rect 42463 24989 42611 25137
rect 34162 24517 34480 24835
rect 42939 24516 43259 24836
rect 42057 24175 42307 24425
rect 42933 23993 43031 24091
rect 42470 23255 42826 23611
rect 42015 22441 42265 22691
rect 42988 22257 43088 22357
rect 42503 21567 42813 21877
rect 42943 21172 43143 21372
rect 42063 20803 42263 21003
rect 42088 14819 42288 15019
rect 41613 14569 41761 14717
rect 42538 4260 42682 4404
rect 42955 127 43061 132
rect 42955 31 42960 127
rect 42960 31 43056 127
rect 43056 31 43061 127
rect 42955 26 43061 31
rect -218 -601 170 -213
rect 41519 -601 41907 -213
rect -678 -1061 -290 -673
rect 41979 -1061 42367 -673
rect -1138 -1521 -750 -1133
rect 42439 -1521 42827 -1133
rect -1598 -1981 -1210 -1593
rect 42899 -1981 43287 -1593
<< metal4 >>
rect -1604 41276 -1204 41283
rect -1604 40888 -1598 41276
rect -1210 40888 -1204 41276
rect -1604 -1593 -1204 40888
rect -1604 -1981 -1598 -1593
rect -1210 -1981 -1204 -1593
rect -1604 -1987 -1204 -1981
rect -1144 40816 -744 41283
rect -1144 40428 -1138 40816
rect -750 40428 -744 40816
rect -1144 -1133 -744 40428
rect -1144 -1521 -1138 -1133
rect -750 -1521 -744 -1133
rect -1144 -1987 -744 -1521
rect -684 40356 -284 41283
rect -684 39968 -678 40356
rect -290 39968 -284 40356
rect -684 -673 -284 39968
rect -684 -1061 -678 -673
rect -290 -1061 -284 -673
rect -684 -1987 -284 -1061
rect -224 39896 176 41283
rect -224 39508 -218 39896
rect 170 39508 176 39896
rect -224 7639 176 39508
rect 34161 41248 34481 41249
rect 34161 40930 34162 41248
rect 34480 40930 34481 41248
rect 34161 36862 34481 40930
rect 34821 40772 35141 40773
rect 34821 40454 34822 40772
rect 35140 40454 35141 40772
rect 34821 36775 35141 40454
rect 41513 39896 41913 41283
rect 41513 39508 41519 39896
rect 41907 39508 41913 39896
rect 34161 24835 34481 28295
rect 34821 25712 35141 28344
rect 34821 25394 34822 25712
rect 35140 25394 35141 25712
rect 34821 25393 35141 25394
rect 34161 24517 34162 24835
rect 34480 24517 34481 24835
rect 34161 24516 34481 24517
rect 41513 14717 41913 39508
rect 41513 14569 41613 14717
rect 41761 14569 41913 14717
rect -224 7237 180 7639
rect -224 -213 176 7237
rect -224 -601 -218 -213
rect 170 -601 176 -213
rect -224 -1987 176 -601
rect 41513 -213 41913 14569
rect 41513 -601 41519 -213
rect 41907 -601 41913 -213
rect 41513 -1987 41913 -601
rect 41973 40356 42373 41283
rect 41973 39968 41979 40356
rect 42367 39968 42373 40356
rect 41973 24425 42373 39968
rect 41973 24175 42057 24425
rect 42307 24175 42373 24425
rect 41973 22691 42373 24175
rect 41973 22441 42015 22691
rect 42265 22441 42373 22691
rect 41973 21003 42373 22441
rect 41973 20803 42063 21003
rect 42263 20803 42373 21003
rect 41973 15019 42373 20803
rect 41973 14819 42088 15019
rect 42288 14819 42373 15019
rect 41973 -673 42373 14819
rect 41973 -1061 41979 -673
rect 42367 -1061 42373 -673
rect 41973 -1987 42373 -1061
rect 42433 40816 42833 41283
rect 42433 40428 42439 40816
rect 42827 40428 42833 40816
rect 42433 25713 42833 40428
rect 42433 25393 42435 25713
rect 42755 25393 42833 25713
rect 42433 25137 42833 25393
rect 42433 24989 42463 25137
rect 42611 24989 42833 25137
rect 42433 23611 42833 24989
rect 42433 23255 42470 23611
rect 42826 23255 42833 23611
rect 42433 21877 42833 23255
rect 42433 21567 42503 21877
rect 42813 21567 42833 21877
rect 42433 4404 42833 21567
rect 42433 4260 42538 4404
rect 42682 4260 42833 4404
rect 42433 -1133 42833 4260
rect 42433 -1521 42439 -1133
rect 42827 -1521 42833 -1133
rect 42433 -1987 42833 -1521
rect 42893 41276 43293 41283
rect 42893 40888 42899 41276
rect 43287 40888 43293 41276
rect 42893 24836 43293 40888
rect 42893 24516 42939 24836
rect 43259 24516 43293 24836
rect 42893 24091 43293 24516
rect 42893 23993 42933 24091
rect 43031 23993 43293 24091
rect 42893 22357 43293 23993
rect 42893 22257 42988 22357
rect 43088 22257 43293 22357
rect 42893 21372 43293 22257
rect 42893 21172 42943 21372
rect 43143 21172 43293 21372
rect 42893 132 43293 21172
rect 42893 26 42955 132
rect 43061 26 43293 132
rect 42893 -1593 43293 26
rect 42893 -1981 42899 -1593
rect 43287 -1981 43293 -1593
rect 42893 -1987 43293 -1981
use por_ana  por_ana_0
timestamp 1713454396
transform 1 0 29373 0 1 25849
box -29373 -25849 13304 13900
use por_dig  por_dig_0
timestamp 1713190415
transform 1 0 29953 0 1 25790
box 0 0 11593 13737
use sky130_fd_pr__nfet_g5v0d10v5_MUZ6AA  sky130_fd_pr__nfet_g5v0d10v5_MUZ6AA_0
timestamp 1713020960
transform 0 1 42184 -1 0 26851
box -989 -358 989 358
use sky130_fd_pr__nfet_g5v0d10v5_RBNV2H  sky130_fd_pr__nfet_g5v0d10v5_RBNV2H_0
timestamp 1713025662
transform 1 0 30369 0 1 38503
box -831 -358 831 358
use sky130_fd_pr__nfet_g5v0d10v5_X6E435  sky130_fd_pr__nfet_g5v0d10v5_X6E435_0
timestamp 1713026030
transform 1 0 -395 0 1 32520
box -357 -358 357 358
<< labels >>
flabel metal3 1723 -1527 1723 -1527 0 FreeSans 1600 0 0 0 dvss
port 4 nsew
flabel metal3 1723 -1987 1723 -1987 0 FreeSans 1600 0 0 0 dvdd
port 3 nsew
flabel metal3 1723 -607 1723 -607 0 FreeSans 1600 0 0 0 avss
port 2 nsew
flabel metal3 1723 -1067 1723 -1067 0 FreeSans 1600 0 0 0 avdd
port 1 nsew
flabel metal3 43093 27013 43293 27073 0 FreeSans 1600 0 0 0 otrip[1]
port 7 nsew
flabel metal3 43093 27409 43293 27469 0 FreeSans 1600 0 0 0 otrip[0]
port 8 nsew
flabel metal3 43093 26674 43293 26734 0 FreeSans 1600 0 0 0 otrip[2]
port 6 nsew
flabel metal2 s 30421 41082 30481 41282 0 FreeSans 1600 90 0 0 force_ena_rc_osc
port 10 nsew
flabel metal2 s 30879 41082 30939 41282 0 FreeSans 1600 90 0 0 force_pdn
port 9 nsew
flabel metal2 s 29921 41082 29981 41282 0 FreeSans 1600 90 0 0 force_dis_rc_osc
port 23 nsew
flabel metal2 s 29342 41082 29402 41282 0 FreeSans 1600 90 0 0 por_timed_out
port 22 nsew
flabel metal2 s 28854 41082 28914 41282 0 FreeSans 1600 90 0 0 osc_ck
port 18 nsew
flabel metal3 s 43093 33308 43293 33368 0 FreeSans 1600 0 0 0 startup_timed_out
port 21 nsew
flabel metal3 s 43093 31948 43293 32008 0 FreeSans 1600 0 0 0 force_short_oneshot
port 11 nsew
flabel metal2 s 26775 41082 26841 41282 0 FreeSans 1600 90 0 0 por
port 17 nsew
flabel metal2 s 26348 41082 26414 41282 0 FreeSans 1600 90 0 0 dcomp
port 24 nsew
flabel metal2 s 12255 41082 12321 41282 0 FreeSans 1600 90 0 0 itest
port 20 nsew
flabel metal2 s 10871 41082 10935 41282 0 FreeSans 1600 90 0 0 vbg_1v2
port 5 nsew
flabel metal3 s 43093 23795 43293 23859 0 FreeSans 1600 0 0 0 isrc_sel
port 12 nsew
flabel metal2 s 14956 41082 15020 41282 0 FreeSans 1600 90 0 0 ibg_200n
port 13 nsew
flabel metal2 s 21267 41082 21331 41282 0 FreeSans 1600 90 0 0 porb_h
port 15 nsew
flabel metal2 s 27432 41082 27496 41282 0 FreeSans 1600 90 0 0 porb
port 16 nsew
flabel metal3 s -1604 32510 -1404 32570 0 FreeSans 1600 0 0 0 vin
port 14 nsew
flabel metal3 s 43093 27737 43293 27797 0 FreeSans 1600 0 0 0 pwup_filt
port 19 nsew
<< end >>
