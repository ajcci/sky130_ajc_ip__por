** sch_path: /home/rtsang/chipalooza/sky130_ajc_ip__por/cace/trip_up_down.sch
**.subckt trip_up_down
Ibias vbp GND 200n
XM1 ibg_200n vbp avdd_bg avdd_bg sky130_fd_pr__pfet_g5v0d10v5 L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'  pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM0 vbp vbp avdd_bg avdd_bg sky130_fd_pr__pfet_g5v0d10v5 L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'  pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
R1 itest GND 1e6 m=1
C1 porb_h GND 20p m=1
Vavss avss GND DC 0
Vforce_pdn force_pdn GND DC 0.0
Vavdd avdd GND pwl (0 2 3m 3.6 6m 2) DC 3.3
.save i(vavdd)
Vbg1v2 vbg_1v2 GND DC 1.2
Vdvss dvss GND DC 0
Vdvdd dvdd GND DC 1.8
.save i(vdvdd)
Vvotrip0 otrip[0] GND DC 1.8
.save i(vvotrip0)
Vvotrip1 otrip[1] GND DC 1.8
.save i(vvotrip1)
Vvotrip2 otrip[2] GND DC 1.8
.save i(vvotrip2)
Vvotrip3 otrip[3] GND DC 1.8
.save i(vvotrip3)
Visrc_sel isrc_sel GND DC 0.0
Vforce_dis_rc_osc force_dis_rc_osc GND DC 1.8
Vforce_short_oneshot force_short_oneshot GND DC 0.0
Vavdd_bg avdd_bg GND DC 3.3
Vforce_ena_rc_osc force_ena_rc_osc GND DC 0.0
xIpor avdd porb_h porb avss dvdd por dvss osc_ck vbg_1v2 dcomp otrip[2] otrip[1] otrip[0] itest force_pdn pwup_filt vin  force_ena_rc_osc force_dis_rc_osc startup_timed_out por_timed_out force_short_oneshot isrc_sel ibg_200n sky130_ajc_ip__por
C2 porb GND 20p m=1
C3 por GND 20p m=1
**** begin user architecture code

* CACE gensim simulation file hysteresis_9
* Generated by CACE gensim, Efabless Corporation (c) 2023
* Find trip voltage by ramping Vavdd, both up and down.

.lib /usr/local/share/pdk/sky130A/libs.tech/combined/sky130.lib.spice tt
.include /usr/local/share/pdk/sky130A/libs.ref/sky130_fd_sc_hvl/spice/sky130_fd_sc_hvl.spice
.include /usr/local/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/spice/sky130_fd_sc_hd.spice

.option TEMP=85
* Flag unsafe operating conditions (exceeds models' specified limits)
.option warn=1

.option reltol=1e-3
.option abstol=1e-3

.save all



.csparam dvdd2=0.9
.control
tran 10u 6m
meas tran otrip_r find v(avdd) when v(dcomp)=$&dvdd2 td=300u rise=1
meas tran otrip_f find v(avdd) when v(dcomp)=$&dvdd2 td=3m fall=1
echo $&otrip_r > ngspice/hysteresis_9.data
echo $&otrip_f >> ngspice/hysteresis_9.data
quit
.endc


**** end user architecture code
**.ends

* expanding   symbol:  xschem/sky130_ajc_ip__por.sym # of pins=22
** sym_path: /home/rtsang/chipalooza/sky130_ajc_ip__por/xschem/sky130_ajc_ip__por.sym
** sch_path: /home/rtsang/chipalooza/sky130_ajc_ip__por/xschem/sky130_ajc_ip__por.sch
.subckt sky130_ajc_ip__por avdd porb_h porb avss dvdd por dvss osc_ck vbg_1v2 dcomp otrip[2] otrip[1] otrip[0] itest force_pdn pwup_filt vin force_ena_rc_osc force_dis_rc_osc startup_timed_out por_timed_out force_short_oneshot isrc_sel ibg_200n
*.ipin avdd
*.ipin avss
*.ipin dvdd
*.ipin dvss
*.ipin vbg_1v2
*.ipin otrip[2],otrip[1],otrip[0]
*.ipin force_pdn
*.ipin force_ena_rc_osc
*.ipin force_short_oneshot
*.ipin isrc_sel
*.ipin ibg_200n
*.opin vin
*.opin porb_h
*.opin porb
*.opin por
*.opin osc_ck
*.opin pwup_filt
*.opin itest
*.opin startup_timed_out
*.opin por_timed_out
*.ipin force_dis_rc_osc
*.opin dcomp
xIana vin otrip_decoded_7_ otrip_decoded_6_ otrip_decoded_5_ otrip_decoded_4_ otrip_decoded_3_ otrip_decoded_2_ otrip_decoded_1_ otrip_decoded_0_ vbg_1v2 avdd itest avss ibg_200n force_pdnb dvdd dvss dcomp isrc_sel pwup_filt osc_ck osc_ena porb_h por_unbuf por porb por_ana
**** begin user architecture code



r0 otrip[0] otrip0 1
r1 otrip[1] otrip1 1
r2 otrip[2] otrip2 1

*XSPICE CO-SIM netlist
.include por_dig.out.spice
xipor_dig dvss dvdd force_dis_rc_osc force_ena_rc_osc force_pdn force_pdnb force_short_oneshot osc_ck osc_ena otrip0 otrip1 otrip2 otrip_decoded_0_ otrip_decoded_1_ otrip_decoded_2_ otrip_decoded_3_ otrip_decoded_4_ otrip_decoded_5_ otrip_decoded_6_ otrip_decoded_7_ por_timed_out por_unbuf pwup_filt startup_timed_out por_dig


**** end user architecture code
.ends


* expanding   symbol:  xschem/por_ana.sym # of pins=19
** sym_path: /home/rtsang/chipalooza/sky130_ajc_ip__por/xschem/por_ana.sym
** sch_path: /home/rtsang/chipalooza/sky130_ajc_ip__por/xschem/por_ana.sch
.subckt por_ana vin otrip_decoded[7] otrip_decoded[6] otrip_decoded[5] otrip_decoded[4] otrip_decoded[3] otrip_decoded[2] otrip_decoded[1] otrip_decoded[0] vbg_1v2 avdd itest avss ibg_200n force_pdnb dvdd dvss dcomp isrc_sel pwup_filt osc_ck osc_ena porb_h por_unbuf por porb
*.ipin vbg_1v2
*.ipin avdd
*.ipin avss
*.ipin dvdd
*.ipin dvss
*.ipin force_pdnb
*.ipin isrc_sel
*.ipin ibg_200n
*.opin pwup_filt
*.opin itest
*.ipin osc_ena
*.opin osc_ck
*.ipin otrip_decoded[7],otrip_decoded[6],otrip_decoded[5],otrip_decoded[4],otrip_decoded[3],otrip_decoded[2],otrip_decoded[1],otrip_decoded[0]
*.opin vin
*.ipin por_unbuf
*.opin porb_h
*.opin por
*.opin porb
*.opin dcomp
xIlvls0 dcomp3v3 dvdd dvss dvss avdd avdd vl sky130_fd_sc_hvl__lsbufhv2lv_1
XC2 dcomp_filt dvss sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=6 m=6
xIlvls0[7] otrip_decoded[7] dvdd dvss dvss avdd avdd otrip_decoded_avdd[7] sky130_fd_sc_hvl__lsbuflv2hv_1
xIlvls0[6] otrip_decoded[6] dvdd dvss dvss avdd avdd otrip_decoded_avdd[6] sky130_fd_sc_hvl__lsbuflv2hv_1
xIlvls0[5] otrip_decoded[5] dvdd dvss dvss avdd avdd otrip_decoded_avdd[5] sky130_fd_sc_hvl__lsbuflv2hv_1
xIlvls0[4] otrip_decoded[4] dvdd dvss dvss avdd avdd otrip_decoded_avdd[4] sky130_fd_sc_hvl__lsbuflv2hv_1
xIlvls0[3] otrip_decoded[3] dvdd dvss dvss avdd avdd otrip_decoded_avdd[3] sky130_fd_sc_hvl__lsbuflv2hv_1
xIlvls0[2] otrip_decoded[2] dvdd dvss dvss avdd avdd otrip_decoded_avdd[2] sky130_fd_sc_hvl__lsbuflv2hv_1
xIlvls0[1] otrip_decoded[1] dvdd dvss dvss avdd avdd otrip_decoded_avdd[1] sky130_fd_sc_hvl__lsbuflv2hv_1
xIlvls0[0] otrip_decoded[0] dvdd dvss dvss avdd avdd otrip_decoded_avdd[0] sky130_fd_sc_hvl__lsbuflv2hv_1
xIlvls1 force_pdnb dvdd dvss dvss avdd avdd force_pdnb_avdd sky130_fd_sc_hvl__lsbuflv2hv_1
xIlvls2 isrc_sel dvdd dvss dvss avdd avdd isrc_sel_avdd sky130_fd_sc_hvl__lsbuflv2hv_1
xIrsmux avdd vin force_pdnb_avdd otrip_decoded_avdd[7] otrip_decoded_avdd[6] otrip_decoded_avdd[5] otrip_decoded_avdd[4] otrip_decoded_avdd[3] otrip_decoded_avdd[2] otrip_decoded_avdd[1] otrip_decoded_avdd[0] vtrip_decoded_avdd[7] vtrip_decoded_avdd[6] vtrip_decoded_avdd[5] vtrip_decoded_avdd[4] vtrip_decoded_avdd[3] vtrip_decoded_avdd[2] vtrip_decoded_avdd[1] vtrip_decoded_avdd[0] not_used avss rstring_mux
xIcomp avdd ibias0 dcomp3v3 force_pdnb_avdd vbg_1v2 vin avss comparator
xIbiasgen avdd ibias0 itest ibias1 ibg_200n vbg_1v2 isrc_sel_avdd force_pdnb_avdd net8 avss ibias_gen
xIosc dvdd osc_ck osc_ena dvss rc_osc
xIlvls3 por_unbuf dvdd dvss dvss avdd avdd net1 sky130_fd_sc_hvl__lsbuflv2hv_1
xIinv4 por_unbuf dvss dvss dvdd dvdd net4 sky130_fd_sc_hd__inv_4
xIinv5 net4 dvss dvss dvdd dvdd por sky130_fd_sc_hd__inv_16
xIinv7 net6 dvss dvss dvdd dvdd net5 sky130_fd_sc_hd__inv_4
xIinv88 net5 dvss dvss dvdd dvdd porb sky130_fd_sc_hd__inv_16
xIinv6 por_unbuf dvss dvss dvdd dvdd net6 sky130_fd_sc_hd__inv_4
xIinv8 net3 avss avss avdd avdd porb_h sky130_fd_sc_hvl__inv_16
xIinv2 net2 avss avss avdd avdd net3 sky130_fd_sc_hvl__inv_4
xIinv1 net1 avss avss avdd avdd net2 sky130_fd_sc_hvl__inv_1
xIschmitt dvdd dcomp_filt vsch dvss schmitt_trigger
xIinv3 net7 dvss dvss dvdd dvdd pwup_filt sky130_fd_sc_hd__inv_16
xIinv9 vsch dvss dvss dvdd dvdd net7 sky130_fd_sc_hd__inv_4
XR2 dcomp_filt vl avss sky130_fd_pr__res_xhigh_po_1p41 L=700 mult=1 m=1
xIlvls3[7] dvss dvdd dvss dvss avdd avdd vtrip_decoded_avdd[7] sky130_fd_sc_hvl__lsbuflv2hv_1
xIlvls3[6] dvss dvdd dvss dvss avdd avdd vtrip_decoded_avdd[6] sky130_fd_sc_hvl__lsbuflv2hv_1
xIlvls3[5] dvss dvdd dvss dvss avdd avdd vtrip_decoded_avdd[5] sky130_fd_sc_hvl__lsbuflv2hv_1
xIlvls3[4] dvss dvdd dvss dvss avdd avdd vtrip_decoded_avdd[4] sky130_fd_sc_hvl__lsbuflv2hv_1
xIlvls3[3] dvss dvdd dvss dvss avdd avdd vtrip_decoded_avdd[3] sky130_fd_sc_hvl__lsbuflv2hv_1
xIlvls3[2] dvss dvdd dvss dvss avdd avdd vtrip_decoded_avdd[2] sky130_fd_sc_hvl__lsbuflv2hv_1
xIlvls3[1] dvss dvdd dvss dvss avdd avdd vtrip_decoded_avdd[1] sky130_fd_sc_hvl__lsbuflv2hv_1
xIlvls3[0] dvss dvdd dvss dvss avdd avdd vtrip_decoded_avdd[0] sky130_fd_sc_hvl__lsbuflv2hv_1
xIcomp_vunder avdd ibias1 net9 avss not_used vbg_1v2 avss comparator
xIlvls5 net9 dvdd dvss dvss avdd avdd vlu sky130_fd_sc_hvl__lsbufhv2lv_1
* noconn vlu
xIinv10 vl dvss dvss dvdd dvdd net10 sky130_fd_sc_hd__inv_4
xIinv11 net10 dvss dvss dvdd dvdd dcomp sky130_fd_sc_hd__inv_16
XQ1 avss avss net8 avss sky130_fd_pr__pnp_05v5_W0p68L0p68 m=1 mult=1
.ends


* expanding   symbol:  rstring_mux.sym # of pins=7
** sym_path: /home/rtsang/chipalooza/sky130_ajc_ip__por/cace/rstring_mux.sym
** sch_path: /home/rtsang/chipalooza/sky130_ajc_ip__por/cace/rstring_mux.sch
.subckt rstring_mux avdd vout_brout ena otrip_decoded_avdd[7] otrip_decoded_avdd[6] otrip_decoded_avdd[5] otrip_decoded_avdd[4] otrip_decoded_avdd[3] otrip_decoded_avdd[2] otrip_decoded_avdd[1] otrip_decoded_avdd[0] vtrip_decoded_avdd[7] vtrip_decoded_avdd[6] vtrip_decoded_avdd[5] vtrip_decoded_avdd[4] vtrip_decoded_avdd[3] vtrip_decoded_avdd[2] vtrip_decoded_avdd[1] vtrip_decoded_avdd[0] vout_vunder avss
*.opin vout_brout
*.ipin otrip_decoded_avdd[7],otrip_decoded_avdd[6],otrip_decoded_avdd[5],otrip_decoded_avdd[4],otrip_decoded_avdd[3],otrip_decoded_avdd[2],otrip_decoded_avdd[1],otrip_decoded_avdd[0]
*.opin vout_vunder
*.ipin vtrip_decoded_avdd[7],vtrip_decoded_avdd[6],vtrip_decoded_avdd[5],vtrip_decoded_avdd[4],vtrip_decoded_avdd[3],vtrip_decoded_avdd[2],vtrip_decoded_avdd[1],vtrip_decoded_avdd[0]
*.ipin ena
*.ipin avdd
*.ipin avss
XR1 net2 net3 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR2 net3 net4 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR0 avss net2 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR3 net4 net5 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR4 net5 net6 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR5 net6 net7 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR6 net7 net8 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR7 net8 net9 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR8 net9 net10 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR9 net10 net11 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR10 net11 net12 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR11 net12 net13 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR12 net13 net14 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR13 net14 net15 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR14 net15 net16 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR15 net16 net17 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR16 net17 net18 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR17 net18 net19 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR18 net19 net20 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR19 net20 net21 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR20 net21 net22 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR21 net22 net23 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR22 net23 net24 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR23 net24 net25 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR24 net25 net26 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR25 net26 net27 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR26 net27 net28 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR27 net28 vtrip7 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR28 vtrip7 vtrip6 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR29 vtrip6 vtrip5 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR30 vtrip5 vtrip4 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR31 vtrip4 vtrip3 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR32 vtrip3 vtrip2 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR33 vtrip2 vtrip1 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR34 vtrip1 vtrip0 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR35 vtrip0 net29 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR36 net29 net30 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR37 net30 net31 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR38 net31 net32 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR39 net32 net33 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR40 net33 net34 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR41 net34 net35 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR42 net35 net36 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR43 net36 net37 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR44 net37 net38 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR45 net38 net39 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR46 net39 net40 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR47 net40 net41 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR48 net41 net42 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR49 net42 net43 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR50 net43 net44 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR51 net44 net45 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR52 net45 net46 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR53 net46 net47 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR54 net47 net48 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR55 net48 net49 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR56 net49 net50 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR57 net50 net51 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR58 net51 net52 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR59 net52 net53 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR60 net53 net54 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR61 net54 net55 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR62 net55 net56 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR63 net56 net57 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR64 net57 net58 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR65 net58 net59 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR66 net59 net60 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR67 net60 net61 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR68 net61 net62 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR69 net62 net1 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XMtp[7] vtrip7 otrip_decoded_b_avdd[7] vout_brout avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)  * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XMtp[6] vtrip6 otrip_decoded_b_avdd[6] vout_brout avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)  * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XMtp[5] vtrip5 otrip_decoded_b_avdd[5] vout_brout avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)  * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XMtp[4] vtrip4 otrip_decoded_b_avdd[4] vout_brout avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)  * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XMtp[3] vtrip3 otrip_decoded_b_avdd[3] vout_brout avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)  * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XMtp[2] vtrip2 otrip_decoded_b_avdd[2] vout_brout avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)  * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XMtp[1] vtrip1 otrip_decoded_b_avdd[1] vout_brout avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)  * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XMtp[0] vtrip0 otrip_decoded_b_avdd[0] vout_brout avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)  * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XMtn[7] vout_brout otrip_decoded_avdd[7] vtrip7 avss sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)  * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XMtn[6] vout_brout otrip_decoded_avdd[6] vtrip6 avss sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)  * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XMtn[5] vout_brout otrip_decoded_avdd[5] vtrip5 avss sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)  * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XMtn[4] vout_brout otrip_decoded_avdd[4] vtrip4 avss sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)  * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XMtn[3] vout_brout otrip_decoded_avdd[3] vtrip3 avss sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)  * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XMtn[2] vout_brout otrip_decoded_avdd[2] vtrip2 avss sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)  * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XMtn[1] vout_brout otrip_decoded_avdd[1] vtrip1 avss sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)  * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XMtn[0] vout_brout otrip_decoded_avdd[0] vtrip0 avss sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)  * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XMtp1[7] vtrip7 vtrip_decoded_b_avdd[7] vout_vunder avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)  * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XMtp1[6] vtrip6 vtrip_decoded_b_avdd[6] vout_vunder avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)  * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XMtp1[5] vtrip5 vtrip_decoded_b_avdd[5] vout_vunder avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)  * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XMtp1[4] vtrip4 vtrip_decoded_b_avdd[4] vout_vunder avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)  * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XMtp1[3] vtrip3 vtrip_decoded_b_avdd[3] vout_vunder avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)  * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XMtp1[2] vtrip2 vtrip_decoded_b_avdd[2] vout_vunder avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)  * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XMtp1[1] vtrip1 vtrip_decoded_b_avdd[1] vout_vunder avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)  * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XMtp1[0] vtrip0 vtrip_decoded_b_avdd[0] vout_vunder avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)  * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XMtn1[7] vout_vunder vtrip_decoded_avdd[7] vtrip7 avss sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)  * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XMtn1[6] vout_vunder vtrip_decoded_avdd[6] vtrip6 avss sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)  * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XMtn1[5] vout_vunder vtrip_decoded_avdd[5] vtrip5 avss sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)  * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XMtn1[4] vout_vunder vtrip_decoded_avdd[4] vtrip4 avss sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)  * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XMtn1[3] vout_vunder vtrip_decoded_avdd[3] vtrip3 avss sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)  * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XMtn1[2] vout_vunder vtrip_decoded_avdd[2] vtrip2 avss sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)  * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XMtn1[1] vout_vunder vtrip_decoded_avdd[1] vtrip1 avss sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)  * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XMtn1[0] vout_vunder vtrip_decoded_avdd[0] vtrip0 avss sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)  * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
xIinv0[7] otrip_decoded_avdd[7] avss avss avdd avdd otrip_decoded_b_avdd[7] sky130_fd_sc_hvl__inv_1
xIinv0[6] otrip_decoded_avdd[6] avss avss avdd avdd otrip_decoded_b_avdd[6] sky130_fd_sc_hvl__inv_1
xIinv0[5] otrip_decoded_avdd[5] avss avss avdd avdd otrip_decoded_b_avdd[5] sky130_fd_sc_hvl__inv_1
xIinv0[4] otrip_decoded_avdd[4] avss avss avdd avdd otrip_decoded_b_avdd[4] sky130_fd_sc_hvl__inv_1
xIinv0[3] otrip_decoded_avdd[3] avss avss avdd avdd otrip_decoded_b_avdd[3] sky130_fd_sc_hvl__inv_1
xIinv0[2] otrip_decoded_avdd[2] avss avss avdd avdd otrip_decoded_b_avdd[2] sky130_fd_sc_hvl__inv_1
xIinv0[1] otrip_decoded_avdd[1] avss avss avdd avdd otrip_decoded_b_avdd[1] sky130_fd_sc_hvl__inv_1
xIinv0[0] otrip_decoded_avdd[0] avss avss avdd avdd otrip_decoded_b_avdd[0] sky130_fd_sc_hvl__inv_1
xIinv1[7] vtrip_decoded_avdd[7] avss avss avdd avdd vtrip_decoded_b_avdd[7] sky130_fd_sc_hvl__inv_1
xIinv1[6] vtrip_decoded_avdd[6] avss avss avdd avdd vtrip_decoded_b_avdd[6] sky130_fd_sc_hvl__inv_1
xIinv1[5] vtrip_decoded_avdd[5] avss avss avdd avdd vtrip_decoded_b_avdd[5] sky130_fd_sc_hvl__inv_1
xIinv1[4] vtrip_decoded_avdd[4] avss avss avdd avdd vtrip_decoded_b_avdd[4] sky130_fd_sc_hvl__inv_1
xIinv1[3] vtrip_decoded_avdd[3] avss avss avdd avdd vtrip_decoded_b_avdd[3] sky130_fd_sc_hvl__inv_1
xIinv1[2] vtrip_decoded_avdd[2] avss avss avdd avdd vtrip_decoded_b_avdd[2] sky130_fd_sc_hvl__inv_1
xIinv1[1] vtrip_decoded_avdd[1] avss avss avdd avdd vtrip_decoded_b_avdd[1] sky130_fd_sc_hvl__inv_1
xIinv1[0] vtrip_decoded_avdd[0] avss avss avdd avdd vtrip_decoded_b_avdd[0] sky130_fd_sc_hvl__inv_1
xIinv2 ena avss avss avdd avdd ena_b sky130_fd_sc_hvl__inv_1
XMpdn net1 ena_b avss avss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2)  * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMpdp avdd ena_b net1 avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf *  0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=16 m=16
XMdum0 vout_brout avdd vout_brout avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)  * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=7 m=7
XMdum1 vout_brout avss vout_brout avss sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)  * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=7 m=7
XMdum2 vout_brout avdd vout_vunder avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)  * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMdum3 vout_vunder avss vout_brout avss sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)  * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMdum4 vout_vunder avdd vout_vunder avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)  * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=7 m=7
XMdum5 vout_vunder avss vout_vunder avss sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2)  * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=7 m=7
.ends


* expanding   symbol:  comparator.sym # of pins=7
** sym_path: /home/rtsang/chipalooza/sky130_ajc_ip__por/cace/comparator.sym
** sch_path: /home/rtsang/chipalooza/sky130_ajc_ip__por/cace/comparator.sch
.subckt comparator avdd ibias out ena vinn vinp avss
*.ipin ena
*.ipin avdd
*.ipin avss
*.ipin ibias
*.ipin vinn
*.ipin vinp
*.opin out
XMb vn vn avss avss sky130_fd_pr__nfet_g5v0d10v5 L=8 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2)  * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XMta vt vn avss avss sky130_fd_pr__nfet_g5v0d10v5 L=8 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2)  * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XMl0 vn ena_b avss avss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2)  * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMinv0 ena_b ena avss avss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2)  * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMinv1 ena_b ena avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2)  * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMi0 vnn vinn vt vt sky130_fd_pr__nfet_g5v0d10v5 L=8 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2)  * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=16 m=16
XMi1 vpp vinp vt vt sky130_fd_pr__nfet_g5v0d10v5 L=8 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2)  * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=16 m=16
XMld1 vpp vpp avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=8 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2)  * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=8 m=8
XMh1 vnn vpp avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=8 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2)  * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=14 m=14
XMh0 vpp vnn avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=8 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2)  * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=14 m=14
XMld0 vnn vnn avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=8 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2)  * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=8 m=8
XMpp1 n0 vpp avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=8 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2)  * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XMnn1 n0 vm avss avss sky130_fd_pr__nfet_g5v0d10v5 L=8 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2)  * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XMpp0 vm vnn avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=8 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2)  * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XMnn0 vm vm avss avss sky130_fd_pr__nfet_g5v0d10v5 L=8 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2)  * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XMinv3 n1 n0 avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2)  * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XMinv2 n1 n0 avss avss sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2)  * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XMinv5 out n1 avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2)  * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=8 m=8
XMinv4 out n1 avss avss sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2)  * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=8 m=8
XMl1 vm ena_b avss avss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2)  * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMl3 vnn ena avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2)  * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMl4 vpp ena avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2)  * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMt1 ibias ena vn avss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2)  * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMt0 vn ena_b ibias avdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2)  * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMl2 n0 ena_b avss avss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2)  * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMdum0 vnn avss vt vt sky130_fd_pr__nfet_g5v0d10v5 L=8 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2)  * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=16 m=16
XMdum1 avss avss avss avss sky130_fd_pr__nfet_g5v0d10v5 L=8 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2)  * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=4 m=4
XMdum2 avdd avdd avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=8 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2)  * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XMdum3 avdd avdd avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=8 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2)  * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=22 m=22
.ends


* expanding   symbol:  ibias_gen.sym # of pins=10
** sym_path: /home/rtsang/chipalooza/sky130_ajc_ip__por/cace/ibias_gen.sym
** sch_path: /home/rtsang/chipalooza/sky130_ajc_ip__por/cace/ibias_gen.sch
.subckt ibias_gen avdd ibias0 itest ibias1 ibg_200n vbg_1v2 isrc_sel ena ve avss
*.ipin vbg_1v2
*.ipin ena
*.opin ibias0
*.ipin ibg_200n
*.ipin isrc_sel
*.ipin avdd
*.ipin avss
*.opin itest
*.ipin ve
*.opin ibias1
XM17 vstart vbg_1v2 vn0 avss sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf  * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=10 m=10
XMt9 vstart ena_b vstartena avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf  * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMn0 vn0 vn0 ve avss sky130_fd_pr__nfet_g5v0d10v5 L=4 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2)  * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XMp0 vn0 vp0 avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=4 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2)  * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XMn1 vp0 vn0 vr avss sky130_fd_pr__nfet_g5v0d10v5 L=4 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2)  * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XMp1 vp0 vp0 avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=4 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2)  * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XMpb0 ibias0 vp avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=4 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2)  * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XMt0 vp0 isrc_sel vp avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2)  * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMt1 vp isrc_sel_b vp0 avss sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf *  0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMl6 vp ena avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=2 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2)  * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMl3 vp0 ena avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=2 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2)  * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMl1 vn0 ena_b avss avss sky130_fd_pr__nfet_g5v0d10v5 L=2 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2)  * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMnn1 vp1 vn1 avss avss sky130_fd_pr__nfet_g5v0d10v5 L=8 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2)  * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=8 m=8
XMnn0 vn1 vn1 avss avss sky130_fd_pr__nfet_g5v0d10v5 L=8 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2)  * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XMl9 vn1 isrc_sel_b avss avss sky130_fd_pr__nfet_g5v0d10v5 L=2 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf *  0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMt6 net1 isrc_sel vn1 avss sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf *  0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMt7 vn1 isrc_sel_b net2 avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf  * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMpp1 vp1 vp1 avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=4 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2)  * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XMt2 vp isrc_sel_b vp1 avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf *  0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMt3 vp1 isrc_sel vp avss sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2)  * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMt4 ibg_200n ena net1 avss sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf *  0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMt5 net2 ena_b ibg_200n avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf  * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMl7 vp1 isrc_sel avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=2 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2)  * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMl8 vp1 ena avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=2 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2)  * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMl10 vn1 ena_b avss avss sky130_fd_pr__nfet_g5v0d10v5 L=2 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2)  * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMl2 vp0 isrc_sel_b avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=2 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf *  0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMl0 vn0 isrc_sel avss avss sky130_fd_pr__nfet_g5v0d10v5 L=2 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2)  * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMt8 vstartena isrc_sel avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) *  W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMn2 ena_b ena avss avss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2)  * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMp2 ena_b ena avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2)  * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMn3 isrc_sel_b isrc_sel avss avss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf  * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMp3 isrc_sel_b isrc_sel avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf  * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMtst itest vp avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=4 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2)  * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XR1 avss vr avss sky130_fd_pr__res_xhigh_po_1p41 L=700 mult=1 m=1
XMdum0 avss avss avss avss sky130_fd_pr__nfet_g5v0d10v5 L=8 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2)  * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=10 m=10
XMdum1 vp0 avss vn0 avss sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2)  * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMdum2 vp avss vp avss sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2)  * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMdum3 vp1 avss vn1 avss sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2)  * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMdum4 ena_b avss isrc_sel_b avss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf  * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMdum5 isrc_sel_b avdd ena_b avdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf  * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMdum6 vp0 avdd avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2)  * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMdum7 vp avdd vp avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2)  * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMdum8 vn1 avdd vp1 avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2)  * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMdum9 avdd avdd avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=4 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2)  * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=4 m=4
XMdum10 avss avss ve avss sky130_fd_pr__nfet_g5v0d10v5 L=4 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2)  * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMdum11 vr avss ve avss sky130_fd_pr__nfet_g5v0d10v5 L=4 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2)  * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMdum12 vr avss avss avss sky130_fd_pr__nfet_g5v0d10v5 L=4 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2)  * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMpb1 ibias1 vp avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=4 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2)  * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
.ends


* expanding   symbol:  rc_osc.sym # of pins=4
** sym_path: /home/rtsang/chipalooza/sky130_ajc_ip__por/cace/rc_osc.sym
** sch_path: /home/rtsang/chipalooza/sky130_ajc_ip__por/cace/rc_osc.sch
.subckt rc_osc dvdd out ena dvss
*.ipin dvdd
*.ipin dvss
*.opin out
*.ipin ena
XM1 m in dvss dvss sky130_fd_pr__nfet_01v8 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2)  * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XM3 m in dvdd dvdd sky130_fd_pr__pfet_01v8 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2)  * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=6 m=6
XM2 m n dvss dvss sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2)  * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM4 m n dvdd dvdd sky130_fd_pr__pfet_01v8 L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2)  * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=3 m=3
XM5 n m dvss dvss sky130_fd_pr__nfet_01v8 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2)  * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM6 n m dvdd dvdd sky130_fd_pr__pfet_01v8 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2)  * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=3 m=3
XM7 out n dvss dvss sky130_fd_pr__nfet_01v8 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2)  * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM8 out n dvdd dvdd sky130_fd_pr__pfet_01v8 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2)  * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=3 m=3
XC1 in dvss sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=6 m=6
XR1 net1 in dvss sky130_fd_pr__res_xhigh_po_1p41 L=111 mult=1 m=1
XM12 in ena dvdd dvdd sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2)  * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM9 out ena vr dvss sky130_fd_pr__nfet_01v8 L=0.18 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2)  * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM10 out ena_b vr dvdd sky130_fd_pr__pfet_01v8 L=0.18 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2)  * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM11 ena_b ena dvss dvss sky130_fd_pr__nfet_01v8 L=0.6 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2)  * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM13 ena_b ena dvdd dvdd sky130_fd_pr__pfet_01v8 L=0.6 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2)  * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XR2 net2 net1 dvss sky130_fd_pr__res_xhigh_po_1p41 L=111 mult=1 m=1
XR3 net3 net2 dvss sky130_fd_pr__res_xhigh_po_1p41 L=111 mult=1 m=1
XR4 net4 net3 dvss sky130_fd_pr__res_xhigh_po_1p41 L=111 mult=1 m=1
XR5 net5 net4 dvss sky130_fd_pr__res_xhigh_po_1p41 L=111 mult=1 m=1
XR6 net6 net5 dvss sky130_fd_pr__res_xhigh_po_1p41 L=111 mult=1 m=1
XR7 net7 net6 dvss sky130_fd_pr__res_xhigh_po_1p41 L=111 mult=1 m=1
XR8 net8 net7 dvss sky130_fd_pr__res_xhigh_po_1p41 L=111 mult=1 m=1
XR9 net9 net8 dvss sky130_fd_pr__res_xhigh_po_1p41 L=111 mult=1 m=1
XR10 vr net9 dvss sky130_fd_pr__res_xhigh_po_1p41 L=111 mult=1 m=1
XMdum0 vr dvss dvss dvss sky130_fd_pr__nfet_01v8 L=0.6 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2)  * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMdum1 out dvss dvss dvss sky130_fd_pr__nfet_01v8 L=0.18 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2)  * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMdum2 m dvss dvss dvss sky130_fd_pr__nfet_01v8 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2)  * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMdum3 n dvss dvss dvss sky130_fd_pr__nfet_01v8 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2)  * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMdum4 m dvdd n dvdd sky130_fd_pr__pfet_01v8 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2)  * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMdum5 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8 L=0.18 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2)  * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMdum6 ena_b dvdd vr dvdd sky130_fd_pr__pfet_01v8 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2)  * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMdum7 dvdd dvdd out dvdd sky130_fd_pr__pfet_01v8 L=0.18 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2)  * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  xschem/schmitt_trigger.sym # of pins=4
** sym_path: /home/rtsang/chipalooza/sky130_ajc_ip__por/xschem/schmitt_trigger.sym
** sch_path: /home/rtsang/chipalooza/sky130_ajc_ip__por/xschem/schmitt_trigger.sch
.subckt schmitt_trigger dvdd in out dvss
*.ipin dvdd
*.ipin dvss
*.opin out
*.ipin in
XM1 m in dvss dvss sky130_fd_pr__nfet_01v8 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2)  * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XM3 m in dvdd dvdd sky130_fd_pr__pfet_01v8 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2)  * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=6 m=6
XM2 m out dvss dvss sky130_fd_pr__nfet_01v8 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2)  * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM4 m out dvdd dvdd sky130_fd_pr__pfet_01v8 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2)  * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=3 m=3
XM5 out m dvss dvss sky130_fd_pr__nfet_01v8 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2)  * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM6 out m dvdd dvdd sky130_fd_pr__pfet_01v8 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2)  * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=3 m=3
XMdum0 m dvss dvss dvss sky130_fd_pr__nfet_01v8 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2)  * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMdum1 dvdd dvdd m dvdd sky130_fd_pr__pfet_01v8 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2)  * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends

.GLOBAL GND
.end
