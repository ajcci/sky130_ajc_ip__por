* NGSPICE file created from por_dig.ext - technology: sky130A

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

.subckt por_dig VGND VPWR force_pdn force_pdnb force_rc_osc force_short_oneshot osc_ck
+ osc_ck_256 osc_ena otrip[0] otrip[1] otrip[2] otrip_decoded[0] otrip_decoded[1]
+ otrip_decoded[2] otrip_decoded[3] otrip_decoded[4] otrip_decoded[5] otrip_decoded[6]
+ otrip_decoded[7] por_timed_out por_unbuf pwup_filt startup_timed_out
XFILLER_0_18_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_200_ _087_ _088_ _068_ VGND VGND VPWR VPWR _027_ sky130_fd_sc_hd__o21ai_1
X_131_ cnt_ck_256\[1\] cnt_ck_256\[0\] cnt_ck_256\[2\] VGND VGND VPWR VPWR _045_ sky130_fd_sc_hd__and3_1
XFILLER_0_0_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_5_56 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_114_ cnt_por\[5\] cnt_por\[7\] cnt_por\[6\] VGND VGND VPWR VPWR _033_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_20_87 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_15_76 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput20 net20 VGND VGND VPWR VPWR por_unbuf sky130_fd_sc_hd__buf_2
XFILLER_0_2_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_21_Right_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_12_Right_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_130_ net40 net37 VGND VGND VPWR VPWR _001_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_5_57 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_113_ _094_ _097_ VGND VGND VPWR VPWR _032_ sky130_fd_sc_hd__nor2_1
Xclkbuf_2_3__f_osc_ck clknet_0_osc_ck VGND VGND VPWR VPWR clknet_2_3__leaf_osc_ck
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_21_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold20 cnt_st\[2\] VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_16_Left_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_15_77 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput8 net8 VGND VGND VPWR VPWR force_pdnb sky130_fd_sc_hd__buf_2
Xoutput21 net21 VGND VGND VPWR VPWR startup_timed_out sky130_fd_sc_hd__buf_2
Xoutput10 net10 VGND VGND VPWR VPWR osc_ena sky130_fd_sc_hd__buf_2
XFILLER_0_5_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_19_Left_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_4_Left_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_189_ cnt_por\[5\] cnt_por\[6\] _032_ net20 net52 VGND VGND VPWR VPWR _081_ sky130_fd_sc_hd__a41o_1
X_112_ cnt_por\[1\] cnt_por\[0\] cnt_por\[3\] cnt_por\[2\] VGND VGND VPWR VPWR _097_
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_21_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold10 cnt_ck_256\[1\] VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__dlygate4sd3_1
Xhold21 cnt_st\[4\] VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_16_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput11 net11 VGND VGND VPWR VPWR otrip_decoded[0] sky130_fd_sc_hd__clkbuf_4
Xoutput9 net9 VGND VGND VPWR VPWR osc_ck_256 sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_20_Left_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_188_ _079_ _080_ net22 VGND VGND VPWR VPWR _023_ sky130_fd_sc_hd__a21o_1
X_111_ cnt_por\[1\] cnt_por\[0\] cnt_por\[3\] cnt_por\[2\] VGND VGND VPWR VPWR _096_
+ sky130_fd_sc_hd__and4_1
Xhold22 cnt_por\[7\] VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__dlygate4sd3_1
Xhold11 cnt_por\[14\] VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_16_98 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput12 net12 VGND VGND VPWR VPWR otrip_decoded[1] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_13_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_187_ cnt_por\[5\] cnt_por\[6\] _032_ net20 VGND VGND VPWR VPWR _080_ sky130_fd_sc_hd__nand4_1
XFILLER_0_19_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_110_ cnt_por\[9\] cnt_por\[8\] VGND VGND VPWR VPWR _095_ sky130_fd_sc_hd__nand2_1
X_239_ clknet_2_2__leaf_osc_ck _030_ net27 VGND VGND VPWR VPWR cnt_por\[13\] sky130_fd_sc_hd__dfrtp_1
Xhold23 cnt_por\[9\] VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_15_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold12 cnt_ck_256\[3\] VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput13 net13 VGND VGND VPWR VPWR otrip_decoded[2] sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_21_90 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_19_Right_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_110 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_98 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_186_ cnt_por\[5\] _032_ net20 cnt_por\[6\] VGND VGND VPWR VPWR _079_ sky130_fd_sc_hd__a31o_1
XFILLER_0_19_77 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_169_ _036_ _038_ net21 net3 VGND VGND VPWR VPWR _067_ sky130_fd_sc_hd__o211a_1
X_238_ clknet_2_2__leaf_osc_ck _029_ net27 VGND VGND VPWR VPWR cnt_por\[12\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_77 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold24 cnt_por\[10\] VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__dlygate4sd3_1
Xhold13 cnt_ck_256\[2\] VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_16_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_91 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput14 net14 VGND VGND VPWR VPWR otrip_decoded[3] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_4_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_185_ _077_ _078_ _068_ VGND VGND VPWR VPWR _022_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_19_89 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_237_ clknet_2_1__leaf_osc_ck _028_ net26 VGND VGND VPWR VPWR cnt_por\[11\] sky130_fd_sc_hd__dfrtp_1
X_099_ net7 VGND VGND VPWR VPWR _093_ sky130_fd_sc_hd__inv_2
X_168_ net23 _066_ cnt_por\[0\] VGND VGND VPWR VPWR _017_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_89 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold14 _046_ VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_16_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_11_Left_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput15 net15 VGND VGND VPWR VPWR otrip_decoded[4] sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_13 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_184_ cnt_por\[5\] _032_ net24 VGND VGND VPWR VPWR _078_ sky130_fd_sc_hd__and3_1
XFILLER_0_21_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_098_ net1 VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__inv_2
X_236_ clknet_2_1__leaf_osc_ck _027_ net26 VGND VGND VPWR VPWR cnt_por\[10\] sky130_fd_sc_hd__dfrtp_1
X_167_ net3 net23 VGND VGND VPWR VPWR _066_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_11_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold15 cnt_ck_256\[4\] VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_16_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_219_ clknet_2_3__leaf_osc_ck _001_ net28 VGND VGND VPWR VPWR cnt_ck_256\[1\] sky130_fd_sc_hd__dfrtp_1
Xoutput16 net16 VGND VGND VPWR VPWR otrip_decoded[5] sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_15_Right_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_3_52 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_13_72 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_25 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_183_ _032_ net24 cnt_por\[5\] VGND VGND VPWR VPWR _077_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_21_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_235_ clknet_2_1__leaf_osc_ck _026_ net28 VGND VGND VPWR VPWR cnt_por\[9\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_166_ net35 _051_ VGND VGND VPWR VPWR _016_ sky130_fd_sc_hd__xnor2_1
Xhold16 cnt_por\[12\] VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__dlygate4sd3_1
X_218_ clknet_2_3__leaf_osc_ck _000_ net27 VGND VGND VPWR VPWR cnt_ck_256\[0\] sky130_fd_sc_hd__dfrtp_1
X_149_ _040_ _055_ _053_ VGND VGND VPWR VPWR _009_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_12_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput17 net17 VGND VGND VPWR VPWR otrip_decoded[6] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_7_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_3_53 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_73 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_182_ _075_ _076_ net22 VGND VGND VPWR VPWR _021_ sky130_fd_sc_hd__a21o_1
XFILLER_0_21_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_234_ clknet_2_1__leaf_osc_ck _025_ net28 VGND VGND VPWR VPWR cnt_por\[8\] sky130_fd_sc_hd__dfrtp_1
X_165_ _044_ _065_ VGND VGND VPWR VPWR _015_ sky130_fd_sc_hd__nand2_1
XFILLER_0_1_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold17 cnt_st\[8\] VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_217_ clknet_2_1__leaf_osc_ck _015_ net26 VGND VGND VPWR VPWR cnt_st\[8\] sky130_fd_sc_hd__dfrtp_1
X_148_ cnt_st\[1\] cnt_st\[0\] net50 VGND VGND VPWR VPWR _055_ sky130_fd_sc_hd__a21oi_1
Xoutput18 net18 VGND VGND VPWR VPWR otrip_decoded[7] sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_15_Left_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_2_2__f_osc_ck clknet_0_osc_ck VGND VGND VPWR VPWR clknet_2_2__leaf_osc_ck
+ sky130_fd_sc_hd__clkbuf_16
XPHY_EDGE_ROW_18_Left_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_44 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_181_ _096_ net24 cnt_por\[4\] VGND VGND VPWR VPWR _076_ sky130_fd_sc_hd__a21o_1
XFILLER_0_19_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_9_64 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_3_Left_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_164_ net47 _064_ VGND VGND VPWR VPWR _065_ sky130_fd_sc_hd__xor2_1
X_233_ clknet_2_1__leaf_osc_ck _024_ net28 VGND VGND VPWR VPWR cnt_por\[7\] sky130_fd_sc_hd__dfrtp_1
Xhold18 cnt_st\[0\] VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_84 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_216_ clknet_2_0__leaf_osc_ck _014_ net26 VGND VGND VPWR VPWR cnt_st\[7\] sky130_fd_sc_hd__dfrtp_1
X_147_ _039_ _054_ net21 net3 VGND VGND VPWR VPWR _008_ sky130_fd_sc_hd__a211o_1
XFILLER_0_7_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_108 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput19 net19 VGND VGND VPWR VPWR por_timed_out sky130_fd_sc_hd__buf_2
XFILLER_0_7_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_20_Right_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_180_ _032_ net24 VGND VGND VPWR VPWR _075_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_0_45 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_65 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_163_ _044_ _063_ _064_ net21 VGND VGND VPWR VPWR _014_ sky130_fd_sc_hd__a31o_1
X_232_ clknet_2_1__leaf_osc_ck _023_ net28 VGND VGND VPWR VPWR cnt_por\[6\] sky130_fd_sc_hd__dfrtp_1
Xhold19 cnt_st\[3\] VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_19_85 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_215_ clknet_2_1__leaf_osc_ck _013_ net28 VGND VGND VPWR VPWR cnt_st\[6\] sky130_fd_sc_hd__dfrtp_1
X_146_ cnt_st\[1\] cnt_st\[0\] VGND VGND VPWR VPWR _054_ sky130_fd_sc_hd__or2_1
X_129_ _036_ _038_ net21 VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__o21a_1
XFILLER_0_1_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout22 _067_ VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__buf_2
XFILLER_0_14_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_0_46 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_162_ net3 _043_ VGND VGND VPWR VPWR _064_ sky130_fd_sc_hd__nand2_1
X_231_ clknet_2_1__leaf_osc_ck _022_ net28 VGND VGND VPWR VPWR cnt_por\[5\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput1 force_pdn VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_10_66 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_214_ clknet_2_1__leaf_osc_ck _012_ net28 VGND VGND VPWR VPWR cnt_st\[5\] sky130_fd_sc_hd__dfrtp_1
X_145_ net48 _053_ VGND VGND VPWR VPWR _007_ sky130_fd_sc_hd__nand2_1
XFILLER_0_7_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_128_ cnt_st\[4\] cnt_st\[8\] _041_ _043_ VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__and4_2
XFILLER_0_7_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_0_47 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout23 net24 VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__buf_2
X_161_ cnt_st\[6\] _058_ cnt_st\[7\] VGND VGND VPWR VPWR _063_ sky130_fd_sc_hd__a21o_1
X_230_ clknet_2_3__leaf_osc_ck _021_ net29 VGND VGND VPWR VPWR cnt_por\[4\] sky130_fd_sc_hd__dfrtp_1
Xinput2 force_rc_osc VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_7_Left_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_67 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_213_ clknet_2_0__leaf_osc_ck _011_ net26 VGND VGND VPWR VPWR cnt_st\[4\] sky130_fd_sc_hd__dfrtp_1
X_144_ net3 net21 VGND VGND VPWR VPWR _053_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_21_88 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_127_ _042_ _043_ VGND VGND VPWR VPWR _044_ sky130_fd_sc_hd__nand2_1
Xfanout24 net20 VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__buf_2
XFILLER_0_18_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_160_ _061_ _062_ net21 VGND VGND VPWR VPWR _013_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_18_Right_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput3 force_short_oneshot VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__clkbuf_2
X_212_ clknet_2_0__leaf_osc_ck _010_ net26 VGND VGND VPWR VPWR cnt_st\[3\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_6_58 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_143_ _051_ _052_ VGND VGND VPWR VPWR _006_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_21_89 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_126_ cnt_st\[5\] cnt_st\[7\] cnt_st\[6\] VGND VGND VPWR VPWR _043_ sky130_fd_sc_hd__and3_1
XFILLER_0_17_20 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_10_Left_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_16_78 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_109_ net6 net5 net4 VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__and3_1
XFILLER_0_8_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput4 otrip[0] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_11_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_211_ clknet_2_0__leaf_osc_ck _009_ net26 VGND VGND VPWR VPWR cnt_st\[2\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_6_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_142_ cnt_ck_256\[6\] _049_ VGND VGND VPWR VPWR _052_ sky130_fd_sc_hd__or2_1
XFILLER_0_2_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_125_ cnt_st\[4\] _041_ VGND VGND VPWR VPWR _042_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_16_79 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_108_ net4 net5 net6 VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__and3b_1
XFILLER_0_0_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout26 net29 VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_3_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput5 otrip[1] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__dlymetal6s2s_1
X_210_ clknet_2_0__leaf_osc_ck _008_ net26 VGND VGND VPWR VPWR cnt_st\[1\] sky130_fd_sc_hd__dfrtp_1
X_141_ cnt_ck_256\[6\] _049_ VGND VGND VPWR VPWR _051_ sky130_fd_sc_hd__nand2_1
XFILLER_0_11_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_124_ cnt_st\[1\] cnt_st\[0\] cnt_st\[3\] cnt_st\[2\] VGND VGND VPWR VPWR _041_ sky130_fd_sc_hd__and4_1
XFILLER_0_17_77 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_107_ net5 net4 net6 VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__and3b_1
XFILLER_0_0_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout27 net29 VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__buf_2
XFILLER_0_18_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput6 otrip[2] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_20_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_140_ _049_ net39 VGND VGND VPWR VPWR _005_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_14_Right_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_123_ cnt_st\[1\] cnt_st\[0\] cnt_st\[2\] VGND VGND VPWR VPWR _040_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_7_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_89 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_106_ net5 net4 net6 VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__nor3b_1
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_14_Left_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_17_80 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout28 net29 VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_17_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput7 pwup_filt VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__dlymetal6s2s_1
XPHY_EDGE_ROW_2_Left_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_199_ net25 net23 net54 VGND VGND VPWR VPWR _088_ sky130_fd_sc_hd__a21oi_1
Xmax_cap25 _035_ VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__clkbuf_1
X_122_ cnt_st\[1\] cnt_st\[0\] VGND VGND VPWR VPWR _039_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_7_61 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_2_1__f_osc_ck clknet_0_osc_ck VGND VGND VPWR VPWR clknet_2_1__leaf_osc_ck
+ sky130_fd_sc_hd__clkbuf_16
X_105_ net6 net5 net4 VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__and3b_1
XFILLER_0_8_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_81 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout29 net31 VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_14_114 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_198_ cnt_por\[10\] net25 _038_ net21 VGND VGND VPWR VPWR _087_ sky130_fd_sc_hd__and4_1
X_121_ _093_ net19 net2 VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__o21bai_1
XFILLER_0_3_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_104_ net6 net4 net5 VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__nor3b_1
XFILLER_0_8_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_241__30 VGND VGND VPWR VPWR net30 _241__30/LO sky130_fd_sc_hd__conb_1
XFILLER_0_5_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_197_ _085_ _086_ _067_ VGND VGND VPWR VPWR _026_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_120_ _036_ _038_ VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__nor2_1
XFILLER_0_3_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_103_ net6 net5 net4 VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__nor3b_1
XFILLER_0_0_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1 cnt_rsb VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_17_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_196_ _035_ net23 VGND VGND VPWR VPWR _086_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_6_Left_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_179_ _073_ _074_ net22 VGND VGND VPWR VPWR _020_ sky130_fd_sc_hd__a21o_1
X_102_ net6 net5 net4 VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__nor3_1
Xclkbuf_0_osc_ck osc_ck VGND VGND VPWR VPWR clknet_0_osc_ck sky130_fd_sc_hd__clkbuf_16
XPHY_EDGE_ROW_9_Left_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_4_54 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2 cnt_rsb_stg1 VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_14_74 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_195_ cnt_por\[8\] _034_ net23 net53 VGND VGND VPWR VPWR _085_ sky130_fd_sc_hd__a31o_1
X_178_ _096_ net24 VGND VGND VPWR VPWR _074_ sky130_fd_sc_hd__nand2_1
XFILLER_0_3_92 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_101_ cnt_por\[4\] VGND VGND VPWR VPWR _094_ sky130_fd_sc_hd__inv_2
XFILLER_0_18_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_4_55 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3 cnt_rsb_stg2 VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_75 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_194_ _083_ _084_ _068_ VGND VGND VPWR VPWR _025_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_3_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_177_ cnt_por\[1\] cnt_por\[0\] cnt_por\[2\] net24 cnt_por\[3\] VGND VGND VPWR VPWR
+ _073_ sky130_fd_sc_hd__a41o_1
X_100_ net37 VGND VGND VPWR VPWR _000_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_229_ clknet_2_3__leaf_osc_ck _020_ net29 VGND VGND VPWR VPWR cnt_por\[3\] sky130_fd_sc_hd__dfrtp_1
Xhold4 cnt_por\[13\] VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_17_Right_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_72 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_193_ cnt_por\[8\] _034_ net23 VGND VGND VPWR VPWR _084_ sky130_fd_sc_hd__and3_1
XFILLER_0_6_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_176_ _071_ _072_ net22 VGND VGND VPWR VPWR _019_ sky130_fd_sc_hd__a21o_1
XFILLER_0_19_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_159_ cnt_st\[6\] _058_ VGND VGND VPWR VPWR _062_ sky130_fd_sc_hd__or2_1
X_228_ clknet_2_3__leaf_osc_ck _019_ net28 VGND VGND VPWR VPWR cnt_por\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold5 net9 VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_192_ _034_ net23 cnt_por\[8\] VGND VGND VPWR VPWR _083_ sky130_fd_sc_hd__a21oi_1
X_175_ cnt_por\[1\] cnt_por\[0\] cnt_por\[2\] net24 VGND VGND VPWR VPWR _072_ sky130_fd_sc_hd__nand4_1
XFILLER_0_18_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_158_ cnt_st\[6\] _058_ VGND VGND VPWR VPWR _061_ sky130_fd_sc_hd__nand2_1
X_227_ clknet_2_3__leaf_osc_ck _018_ net28 VGND VGND VPWR VPWR cnt_por\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_20_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold6 _016_ VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_13_Left_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_1_48 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_191_ _081_ _082_ net22 VGND VGND VPWR VPWR _024_ sky130_fd_sc_hd__a21o_1
XFILLER_0_6_107 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_1_Left_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_243_ clknet_2_2__leaf_osc_ck net33 net7 VGND VGND VPWR VPWR cnt_rsb sky130_fd_sc_hd__dfrtp_1
X_174_ cnt_por\[1\] cnt_por\[0\] net23 cnt_por\[2\] VGND VGND VPWR VPWR _071_ sky130_fd_sc_hd__a31o_1
XFILLER_0_2_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_157_ _059_ _060_ net21 VGND VGND VPWR VPWR _012_ sky130_fd_sc_hd__a21o_1
X_226_ clknet_2_3__leaf_osc_ck _017_ net29 VGND VGND VPWR VPWR cnt_por\[0\] sky130_fd_sc_hd__dfrtp_4
Xhold7 cnt_ck_256\[0\] VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_209_ clknet_2_0__leaf_osc_ck _007_ net26 VGND VGND VPWR VPWR cnt_st\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_13_Right_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_1_49 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_2_0__f_osc_ck clknet_0_osc_ck VGND VGND VPWR VPWR clknet_2_0__leaf_osc_ck
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_13_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_190_ _034_ net23 VGND VGND VPWR VPWR _082_ sky130_fd_sc_hd__nand2_1
XFILLER_0_6_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_11_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_242_ clknet_2_0__leaf_osc_ck net32 net7 VGND VGND VPWR VPWR cnt_rsb_stg2 sky130_fd_sc_hd__dfrtp_1
X_173_ _069_ _070_ net22 VGND VGND VPWR VPWR _018_ sky130_fd_sc_hd__a21o_1
X_156_ net3 cnt_st\[5\] _042_ VGND VGND VPWR VPWR _060_ sky130_fd_sc_hd__or3_1
X_225_ clknet_2_2__leaf_osc_ck net36 net27 VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__dfrtp_1
Xhold8 cnt_ck_256\[5\] VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_208_ net41 _092_ VGND VGND VPWR VPWR _031_ sky130_fd_sc_hd__xor2_1
X_139_ cnt_ck_256\[4\] _047_ net38 VGND VGND VPWR VPWR _050_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_17_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_241_ clknet_2_0__leaf_osc_ck net30 net7 VGND VGND VPWR VPWR cnt_rsb_stg1 sky130_fd_sc_hd__dfrtp_1
X_172_ cnt_por\[1\] cnt_por\[0\] net24 VGND VGND VPWR VPWR _070_ sky130_fd_sc_hd__nand3_1
XFILLER_0_3_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_155_ _058_ VGND VGND VPWR VPWR _059_ sky130_fd_sc_hd__inv_2
X_224_ clknet_2_2__leaf_osc_ck _006_ net27 VGND VGND VPWR VPWR cnt_ck_256\[6\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold9 _050_ VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__dlygate4sd3_1
X_207_ net34 _091_ VGND VGND VPWR VPWR _030_ sky130_fd_sc_hd__xor2_1
X_138_ cnt_ck_256\[4\] cnt_ck_256\[5\] _047_ VGND VGND VPWR VPWR _049_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_17_Left_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_110 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_50 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_240_ clknet_2_3__leaf_osc_ck _031_ net29 VGND VGND VPWR VPWR cnt_por\[14\] sky130_fd_sc_hd__dfrtp_1
X_171_ cnt_por\[0\] net24 cnt_por\[1\] VGND VGND VPWR VPWR _069_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_5_Left_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_12_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_223_ clknet_2_2__leaf_osc_ck _005_ net27 VGND VGND VPWR VPWR cnt_ck_256\[5\] sky130_fd_sc_hd__dfrtp_1
X_154_ net3 _042_ cnt_st\[5\] VGND VGND VPWR VPWR _058_ sky130_fd_sc_hd__o21a_1
X_206_ net22 _087_ cnt_por\[11\] _037_ VGND VGND VPWR VPWR _092_ sky130_fd_sc_hd__o211a_1
X_137_ net45 _047_ VGND VGND VPWR VPWR _004_ sky130_fd_sc_hd__xor2_1
XFILLER_0_0_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_8_Left_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_2_51 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_170_ net3 net23 VGND VGND VPWR VPWR _068_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_21_Left_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_12_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_153_ _042_ _057_ _053_ VGND VGND VPWR VPWR _011_ sky130_fd_sc_hd__o21ai_1
X_222_ clknet_2_2__leaf_osc_ck _004_ net27 VGND VGND VPWR VPWR cnt_ck_256\[4\] sky130_fd_sc_hd__dfrtp_1
X_205_ net46 _089_ VGND VGND VPWR VPWR _029_ sky130_fd_sc_hd__xnor2_1
X_136_ _047_ _048_ VGND VGND VPWR VPWR _003_ sky130_fd_sc_hd__nor2_1
X_119_ cnt_por\[11\] cnt_por\[14\] cnt_por\[10\] _037_ VGND VGND VPWR VPWR _038_ sky130_fd_sc_hd__nand4_2
XFILLER_0_12_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_152_ net51 _041_ VGND VGND VPWR VPWR _057_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_8_62 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_221_ clknet_2_2__leaf_osc_ck _003_ net26 VGND VGND VPWR VPWR cnt_ck_256\[3\] sky130_fd_sc_hd__dfrtp_1
X_204_ net22 _087_ cnt_por\[12\] cnt_por\[11\] VGND VGND VPWR VPWR _091_ sky130_fd_sc_hd__o211a_1
X_135_ net42 _045_ VGND VGND VPWR VPWR _048_ sky130_fd_sc_hd__nor2_1
XFILLER_0_9_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_18_82 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_118_ cnt_por\[12\] cnt_por\[13\] VGND VGND VPWR VPWR _037_ sky130_fd_sc_hd__and2_1
XFILLER_0_16_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_151_ _041_ _056_ _053_ VGND VGND VPWR VPWR _010_ sky130_fd_sc_hd__o21ai_1
X_220_ clknet_2_3__leaf_osc_ck _002_ net27 VGND VGND VPWR VPWR cnt_ck_256\[2\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_8_63 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_203_ _089_ _090_ VGND VGND VPWR VPWR _028_ sky130_fd_sc_hd__and2_1
X_134_ cnt_ck_256\[3\] _045_ VGND VGND VPWR VPWR _047_ sky130_fd_sc_hd__and2_1
XFILLER_0_19_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_83 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_117_ _094_ _095_ _097_ _033_ VGND VGND VPWR VPWR _036_ sky130_fd_sc_hd__or4_1
XFILLER_0_6_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_150_ net49 _040_ VGND VGND VPWR VPWR _056_ sky130_fd_sc_hd__nor2_1
XFILLER_0_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_16_Right_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_202_ cnt_por\[11\] net22 _087_ VGND VGND VPWR VPWR _090_ sky130_fd_sc_hd__or3_1
X_133_ _045_ net44 VGND VGND VPWR VPWR _002_ sky130_fd_sc_hd__nor2_1
XFILLER_0_19_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_116_ _094_ _095_ _097_ _033_ VGND VGND VPWR VPWR _035_ sky130_fd_sc_hd__nor4_1
XPHY_EDGE_ROW_12_Left_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_0_Left_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_201_ net22 _087_ cnt_por\[11\] VGND VGND VPWR VPWR _089_ sky130_fd_sc_hd__o21ai_1
X_132_ net40 cnt_ck_256\[0\] net43 VGND VGND VPWR VPWR _046_ sky130_fd_sc_hd__a21oi_1
X_115_ _094_ _097_ _033_ VGND VGND VPWR VPWR _034_ sky130_fd_sc_hd__nor3_1
XFILLER_0_21_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_86 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
.ends

