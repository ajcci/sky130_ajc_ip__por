magic
tech sky130A
magscale 1 2
timestamp 1712986583
<< error_s >>
rect 39865 24944 39991 24960
rect 39827 23173 39828 23227
rect 39865 23210 39990 23226
rect 39887 23123 39888 23173
rect 39887 22853 39888 22937
rect 392 14217 426 14753
<< pwell >>
rect -1182 40391 42901 40527
rect -1182 -559 -1046 40391
rect 42765 -559 42901 40391
rect -1182 -695 42901 -559
<< psubdiff >>
rect -1146 40457 -1086 40491
rect 42805 40457 42865 40491
rect -1146 40431 -1112 40457
rect -1146 -625 -1112 -599
rect 42831 40431 42865 40457
rect 42831 -625 42865 -599
rect -1146 -659 -1086 -625
rect 42805 -659 42865 -625
<< psubdiffcont >>
rect -1086 40457 42805 40491
rect -1146 -599 -1112 40431
rect 42831 -599 42865 40431
rect -1086 -659 42805 -625
<< locali >>
rect -1146 40457 -1086 40491
rect 42805 40457 42865 40491
rect -1146 40431 -1112 40457
rect -1146 -625 -1112 -599
rect 42831 40431 42865 40457
rect 42831 -625 42865 -599
rect -1146 -659 -1086 -625
rect 42805 -659 42865 -625
<< viali >>
rect -1086 40457 42805 40491
rect -1146 -556 -1112 40404
rect 42831 -567 42865 40393
rect -1086 -659 42805 -625
<< metal1 >>
rect 41177 40601 41325 40612
rect 41177 40531 41188 40601
rect -1186 40491 41188 40531
rect 41314 40531 41325 40601
rect 41314 40491 42905 40531
rect -1186 40457 -1086 40491
rect 42805 40457 42905 40491
rect -1186 40404 42905 40457
rect -1186 -556 -1146 40404
rect -1112 40393 42905 40404
rect -1112 40391 42831 40393
rect -1112 -556 -1046 40391
rect 42765 25388 42831 40391
rect 42764 25281 42831 25388
rect 41034 24175 41174 24425
rect 41424 24175 41430 24425
rect 41158 24106 41256 24147
rect 41158 24091 41475 24106
rect 41256 24049 41475 24091
rect 41158 23987 41256 23993
rect 41078 23255 41084 23611
rect 41440 23255 41446 23611
rect 41020 22441 41224 22691
rect 41474 22441 41480 22691
rect 41193 22357 41716 22413
rect 41193 22313 41616 22357
rect 41616 22251 41716 22257
rect 41039 21567 41045 21877
rect 41355 21567 41361 21877
rect -1186 -559 -1046 -556
rect 42765 -559 42831 25281
rect -1186 -567 42831 -559
rect 42865 -567 42905 40393
rect -1186 -625 42905 -567
rect -1186 -659 -1086 -625
rect 42805 -659 42905 -625
rect -1186 -699 42905 -659
<< via1 >>
rect 41188 40491 41314 40601
rect 41188 40475 41314 40491
rect 41266 24989 41414 25137
rect 41174 24175 41424 24425
rect 41158 23993 41256 24091
rect 41084 23255 41440 23611
rect 41224 22441 41474 22691
rect 41616 22257 41716 22357
rect 41045 21567 41355 21877
<< metal2 >>
rect 1111 40272 1507 40292
rect 1111 39982 1131 40272
rect 1471 39982 1507 40272
rect 1111 39265 1507 39982
rect 1577 39865 1962 39896
rect 1577 39606 1599 39865
rect 1934 39606 1962 39865
rect 1577 39251 1962 39606
rect 10871 32731 10935 41282
rect 10871 32667 11144 32731
rect 11080 32217 11144 32667
rect 11841 26826 11850 26892
rect 11916 26826 11925 26892
rect 12255 26887 12321 41282
rect 12255 26831 12260 26887
rect 12316 26831 12321 26887
rect 12255 26826 12321 26831
rect 11850 26541 11916 26826
rect 12260 26822 12316 26826
rect 14078 23704 14142 23713
rect 14956 23700 15020 41282
rect 21267 37305 21331 41282
rect 25575 37439 25631 37446
rect 25573 37437 25633 37439
rect 25573 37381 25575 37437
rect 25631 37381 25633 37437
rect 19650 35406 19710 35408
rect 19643 35350 19652 35406
rect 19708 35350 19717 35406
rect 14956 23644 14960 23700
rect 15016 23644 15020 23700
rect 14956 23640 15020 23644
rect 14078 23631 14142 23640
rect 14960 23635 15016 23640
rect 15162 4251 15222 4260
rect 15162 3329 15222 4191
rect 19650 3696 19710 35350
rect 25573 32795 25633 37381
rect 26348 30339 26414 41282
rect 26775 30842 26841 41282
rect 27432 33447 27496 41282
rect 28854 35411 28914 41282
rect 28847 35406 28921 35411
rect 28847 35350 28856 35406
rect 28912 35350 28921 35406
rect 28847 35341 28921 35350
rect 27235 33383 27496 33447
rect 26348 30283 26353 30339
rect 26409 30283 26414 30339
rect 26348 30278 26414 30283
rect 26766 30278 26775 30344
rect 26841 30278 26850 30344
rect 26353 30274 26409 30278
rect 26775 29996 26841 30278
rect 26795 27891 26851 27900
rect 26795 27826 26851 27835
rect 21332 27605 21388 27612
rect 21330 27603 21390 27605
rect 21330 27547 21332 27603
rect 21388 27547 21390 27603
rect 21147 26295 21203 26302
rect 21145 26293 21205 26295
rect 21145 26237 21147 26293
rect 21203 26237 21205 26293
rect 19899 26133 19959 26142
rect 19899 4249 19959 26073
rect 21145 22193 21205 26237
rect 21330 23778 21390 27547
rect 23589 27323 23645 27330
rect 23587 27321 23647 27323
rect 23587 27265 23589 27321
rect 23645 27265 23647 27321
rect 23128 26451 23184 26458
rect 23126 26449 23186 26451
rect 23126 26393 23128 26449
rect 23184 26393 23186 26449
rect 23126 23796 23186 26393
rect 23126 23736 23490 23796
rect 23587 22311 23647 27265
rect 27235 27077 27299 33383
rect 29342 32686 29402 41282
rect 29921 39211 29981 41282
rect 30421 39463 30481 41282
rect 30421 39403 30724 39463
rect 29921 39155 29923 39211
rect 29979 39155 29981 39211
rect 29921 39153 29981 39155
rect 30471 39153 30480 39213
rect 30540 39153 30549 39213
rect 29923 39146 29979 39153
rect 29342 32630 29344 32686
rect 29400 32630 29402 32686
rect 29342 32628 29402 32630
rect 29344 32621 29400 32628
rect 30480 32006 30540 39153
rect 30480 31950 30482 32006
rect 30538 31950 30540 32006
rect 30480 31948 30540 31950
rect 30482 31941 30538 31948
rect 30338 31328 30394 31335
rect 30336 31326 30396 31328
rect 30336 31270 30338 31326
rect 30394 31270 30396 31326
rect 30336 27893 30396 31270
rect 30336 27824 30396 27833
rect 30481 30627 30541 30636
rect 25406 27025 25462 27032
rect 25404 27023 25464 27025
rect 25404 26967 25406 27023
rect 25462 26967 25464 27023
rect 25404 23416 25464 26967
rect 27864 26893 27920 26900
rect 27862 26891 27922 26893
rect 27862 26835 27864 26891
rect 27920 26835 27922 26891
rect 25564 26752 25620 26759
rect 25562 26750 25622 26752
rect 25562 26694 25564 26750
rect 25620 26694 25622 26750
rect 25562 23807 25622 26694
rect 27653 26590 27709 26597
rect 27651 26588 27711 26590
rect 27651 26532 27653 26588
rect 27709 26532 27711 26588
rect 27651 23763 27711 26532
rect 25404 23356 25603 23416
rect 23436 22251 23647 22311
rect 21145 22133 21389 22193
rect 23436 22068 23496 22251
rect 25543 22062 25603 23356
rect 27862 22350 27922 26835
rect 30481 26131 30541 30567
rect 30664 29966 30724 39403
rect 30664 29910 30666 29966
rect 30722 29910 30724 29966
rect 30664 29908 30724 29910
rect 30666 29901 30722 29908
rect 30879 28611 30939 41282
rect 41177 40603 41325 40612
rect 41177 40473 41186 40603
rect 41316 40473 41325 40603
rect 41177 40464 41325 40473
rect 35756 37439 35834 37448
rect 35756 37379 35765 37439
rect 35825 37379 35834 37439
rect 35756 37370 35834 37379
rect 31041 29424 31097 29431
rect 31039 29422 31099 29424
rect 31039 29366 31041 29422
rect 31097 29366 31099 29422
rect 30872 28606 30946 28611
rect 30872 28550 30881 28606
rect 30937 28550 30946 28606
rect 30872 28540 30946 28550
rect 30481 26075 30483 26131
rect 30539 26075 30541 26131
rect 30481 26073 30541 26075
rect 31039 26126 31099 29366
rect 32536 27605 32614 27614
rect 32536 27545 32545 27605
rect 32605 27545 32614 27605
rect 32536 27536 32614 27545
rect 31984 27469 32062 27478
rect 31984 27409 31993 27469
rect 32053 27409 32062 27469
rect 31984 27400 32062 27409
rect 33180 27323 33258 27332
rect 33180 27263 33189 27323
rect 33249 27263 33258 27323
rect 33877 27321 33902 27340
rect 33180 27254 33258 27263
rect 33824 27312 33902 27321
rect 33824 27252 33833 27312
rect 33893 27252 33902 27312
rect 33824 27243 33902 27252
rect 34468 27154 34546 27163
rect 34468 27094 34477 27154
rect 34537 27094 34546 27154
rect 34468 27085 34546 27094
rect 34744 27025 34822 27034
rect 34744 26965 34753 27025
rect 34813 26965 34822 27025
rect 34744 26956 34822 26965
rect 35756 26893 35834 26902
rect 35756 26833 35765 26893
rect 35825 26833 35834 26893
rect 35756 26824 35834 26833
rect 36400 26752 36478 26761
rect 36400 26692 36409 26752
rect 36469 26692 36478 26752
rect 36400 26683 36478 26692
rect 37069 26599 37097 26632
rect 37053 26590 37113 26599
rect 37053 26521 37113 26530
rect 37713 26460 37741 26674
rect 37697 26451 37757 26460
rect 37697 26382 37757 26391
rect 38357 26304 38385 26677
rect 38341 26295 38401 26304
rect 38341 26226 38401 26235
rect 38073 26126 38129 26133
rect 30483 26066 30539 26073
rect 31039 26057 31099 26066
rect 38071 26124 38131 26126
rect 38071 26068 38073 26124
rect 38129 26068 38131 26124
rect 27666 22290 27922 22350
rect 27666 22067 27726 22290
rect 38071 22163 38131 26068
rect 41257 25137 41423 25146
rect 41257 24989 41266 25137
rect 41414 24989 41423 25137
rect 41257 24980 41423 24989
rect 41165 24425 41433 24434
rect 41165 24175 41174 24425
rect 41424 24175 41433 24425
rect 41165 24166 41433 24175
rect 41149 24091 41265 24100
rect 41149 23993 41158 24091
rect 41256 23993 41265 24091
rect 41149 23984 41265 23993
rect 38223 23859 38286 23861
rect 38223 23732 38286 23795
rect 41075 23611 41449 23620
rect 41075 23255 41084 23611
rect 41440 23255 41449 23611
rect 41075 23246 41449 23255
rect 41215 22691 41483 22700
rect 41215 22441 41224 22691
rect 41474 22441 41483 22691
rect 41215 22432 41483 22441
rect 41606 22357 41725 22366
rect 41606 22257 41616 22357
rect 41716 22257 41725 22357
rect 41606 22248 41725 22257
rect 38071 22103 38286 22163
rect 41036 21877 41364 21886
rect 41036 21567 41045 21877
rect 41355 21567 41364 21877
rect 41036 21558 41364 21567
rect 19899 4193 19901 4249
rect 19957 4193 19959 4249
rect 19899 4191 19959 4193
rect 19901 4184 19957 4191
rect 19650 3627 19710 3636
rect 10 -707 396 1690
rect 493 -110 893 1899
rect 493 -519 893 -510
rect 10 -1039 28 -707
rect 383 -1039 396 -707
rect 10 -1056 396 -1039
<< via2 >>
rect 1131 39982 1471 40272
rect 1599 39606 1934 39865
rect 11850 26826 11916 26892
rect 12260 26831 12316 26887
rect 14078 23640 14142 23704
rect 25575 37381 25631 37437
rect 19652 35350 19708 35406
rect 14960 23644 15016 23700
rect 15162 4191 15222 4251
rect 28856 35350 28912 35406
rect 26353 30283 26409 30339
rect 26775 30278 26841 30344
rect 26795 27835 26851 27891
rect 21332 27547 21388 27603
rect 21147 26237 21203 26293
rect 19899 26073 19959 26133
rect 23589 27265 23645 27321
rect 23128 26393 23184 26449
rect 29923 39155 29979 39211
rect 30480 39153 30540 39213
rect 29344 32630 29400 32686
rect 30482 31950 30538 32006
rect 30338 31270 30394 31326
rect 30336 27833 30396 27893
rect 30481 30567 30541 30627
rect 25406 26967 25462 27023
rect 27864 26835 27920 26891
rect 25564 26694 25620 26750
rect 27653 26532 27709 26588
rect 30666 29910 30722 29966
rect 41186 40601 41316 40603
rect 41186 40475 41188 40601
rect 41188 40475 41314 40601
rect 41314 40475 41316 40601
rect 41186 40473 41316 40475
rect 35765 37379 35825 37439
rect 31041 29366 31097 29422
rect 30881 28550 30937 28606
rect 30483 26075 30539 26131
rect 32545 27545 32605 27605
rect 31993 27409 32053 27469
rect 33189 27263 33249 27323
rect 33833 27252 33893 27312
rect 34477 27094 34537 27154
rect 34753 26965 34813 27025
rect 35765 26833 35825 26893
rect 36409 26692 36469 26752
rect 37053 26530 37113 26590
rect 37697 26391 37757 26451
rect 38341 26235 38401 26295
rect 31039 26066 31099 26126
rect 38073 26068 38129 26124
rect 41266 24989 41414 25137
rect 41174 24175 41424 24425
rect 41158 23993 41256 24091
rect 38222 23795 38286 23859
rect 41084 23255 41440 23611
rect 41224 22441 41474 22691
rect 41616 22257 41716 22357
rect 41045 21567 41355 21877
rect 19901 4193 19957 4249
rect 19650 3636 19710 3696
rect 493 -510 893 -110
rect 28 -1039 383 -707
<< metal3 >>
rect -1604 41276 43293 41282
rect -1604 40888 -1598 41276
rect -1210 41248 42899 41276
rect -1210 40930 34162 41248
rect 34480 40930 42899 41248
rect -1210 40888 42899 40930
rect 43287 40888 43293 41276
rect -1604 40882 43293 40888
rect -1604 40816 43293 40822
rect -1604 40428 -1138 40816
rect -750 40772 42439 40816
rect -750 40454 34822 40772
rect 35140 40603 42439 40772
rect 35140 40473 41186 40603
rect 41316 40473 42439 40603
rect 35140 40454 42439 40473
rect -750 40428 42439 40454
rect 42827 40428 43293 40816
rect -1604 40422 43293 40428
rect -1604 40356 43293 40362
rect -1604 39968 -678 40356
rect -290 40272 41979 40356
rect -290 39982 1131 40272
rect 1471 39982 41979 40272
rect -290 39968 41979 39982
rect 42367 39968 43293 40356
rect -1604 39962 43293 39968
rect -1604 39896 43293 39902
rect -1604 39508 -218 39896
rect 170 39865 41519 39896
rect 170 39606 1599 39865
rect 1934 39606 41519 39865
rect 170 39508 41519 39606
rect 41907 39508 43293 39896
rect -1604 39502 43293 39508
rect 947 39492 1357 39502
rect 29918 39213 29984 39216
rect 30475 39213 30545 39218
rect 29918 39211 30480 39213
rect 29918 39155 29923 39211
rect 29979 39155 30480 39211
rect 29918 39153 30480 39155
rect 30540 39153 30545 39213
rect 29918 39150 29984 39153
rect 30475 39148 30545 39153
rect 25570 37439 25636 37442
rect 35760 37439 35830 37444
rect 25570 37437 35765 37439
rect 25570 37381 25575 37437
rect 25631 37381 35765 37437
rect 25570 37379 35765 37381
rect 35825 37379 35830 37439
rect 25570 37376 25636 37379
rect 35760 37374 35830 37379
rect 19647 35408 19713 35411
rect 28851 35408 28917 35411
rect 19647 35406 30837 35408
rect 19647 35350 19652 35406
rect 19708 35350 28856 35406
rect 28912 35350 30837 35406
rect 19647 35348 30837 35350
rect 19647 35345 19713 35348
rect 28851 35345 28917 35348
rect 40579 33308 43293 33368
rect 29339 32688 29405 32691
rect 29339 32686 30842 32688
rect 29339 32630 29344 32686
rect 29400 32630 30842 32686
rect 29339 32628 30842 32630
rect 29339 32625 29405 32628
rect -1604 32510 4716 32570
rect 30477 32008 30543 32011
rect 30477 32006 30829 32008
rect 30477 31950 30482 32006
rect 30538 31950 30829 32006
rect 30477 31948 30829 31950
rect 40619 31948 43293 32008
rect 30477 31945 30543 31948
rect 30333 31328 30399 31331
rect 30333 31326 30828 31328
rect 30333 31270 30338 31326
rect 30394 31270 30828 31326
rect 30333 31268 30828 31270
rect 30333 31265 30399 31268
rect 30476 30627 30546 30632
rect 30476 30567 30481 30627
rect 30541 30567 30546 30627
rect 30476 30562 30546 30567
rect 26770 30344 26846 30349
rect 26348 30339 26775 30344
rect 26348 30283 26353 30339
rect 26409 30283 26775 30339
rect 26348 30278 26775 30283
rect 26841 30278 26846 30344
rect 26770 30273 26846 30278
rect 30661 29968 30727 29971
rect 30661 29966 30851 29968
rect 30661 29910 30666 29966
rect 30722 29910 30851 29966
rect 30661 29908 30851 29910
rect 30661 29905 30727 29908
rect 31036 29424 31102 29427
rect 31036 29422 31140 29424
rect 31036 29366 31041 29422
rect 31097 29366 31140 29422
rect 31036 29364 31140 29366
rect 31036 29361 31120 29364
rect 30876 28606 30942 28611
rect 30876 28550 30881 28606
rect 30937 28550 30942 28606
rect 30876 28545 30942 28550
rect 26790 27893 26856 27896
rect 30331 27893 30401 27898
rect 26790 27891 30336 27893
rect 26790 27835 26795 27891
rect 26851 27835 30336 27891
rect 26790 27833 30336 27835
rect 30396 27833 34089 27893
rect 26790 27830 26856 27833
rect 30331 27828 30401 27833
rect 34029 27797 34089 27833
rect 34029 27737 43293 27797
rect 21327 27605 21393 27608
rect 32540 27605 32610 27610
rect 21327 27603 32545 27605
rect 21327 27547 21332 27603
rect 21388 27547 32545 27603
rect 21327 27545 32545 27547
rect 32605 27545 32610 27605
rect 21327 27542 21393 27545
rect 32540 27540 32610 27545
rect 31988 27469 32058 27474
rect 31988 27409 31993 27469
rect 32053 27409 43293 27469
rect 31988 27404 32058 27409
rect 23584 27323 23650 27326
rect 33184 27323 33254 27328
rect 23584 27321 33189 27323
rect 23584 27265 23589 27321
rect 23645 27265 33189 27321
rect 23584 27263 33189 27265
rect 33249 27263 33254 27323
rect 23584 27260 23650 27263
rect 33184 27258 33254 27263
rect 33828 27312 33898 27317
rect 33828 27252 33833 27312
rect 33893 27252 41440 27312
rect 33828 27247 33898 27252
rect 34472 27154 34542 27159
rect 34472 27094 34477 27154
rect 34537 27094 41186 27154
rect 34472 27089 34542 27094
rect 25401 27025 25467 27028
rect 34748 27025 34818 27030
rect 25401 27023 34753 27025
rect 25401 26967 25406 27023
rect 25462 26967 34753 27023
rect 25401 26965 34753 26967
rect 34813 26965 34818 27025
rect 25401 26962 25467 26965
rect 34748 26960 34818 26965
rect 11845 26892 11921 26897
rect 27859 26893 27925 26896
rect 35760 26893 35830 26898
rect 11845 26826 11850 26892
rect 11916 26887 12321 26892
rect 11916 26831 12260 26887
rect 12316 26831 12321 26887
rect 11916 26826 12321 26831
rect 27859 26891 35765 26893
rect 27859 26835 27864 26891
rect 27920 26835 35765 26891
rect 27859 26833 35765 26835
rect 35825 26833 35830 26893
rect 27859 26830 27925 26833
rect 35760 26828 35830 26833
rect 11845 26821 11921 26826
rect 25559 26752 25625 26755
rect 36404 26752 36474 26757
rect 25559 26750 36409 26752
rect 25559 26694 25564 26750
rect 25620 26694 36409 26750
rect 25559 26692 36409 26694
rect 36469 26692 36474 26752
rect 25559 26689 25625 26692
rect 36404 26687 36474 26692
rect 41126 26734 41186 27094
rect 41380 27073 41440 27252
rect 41380 27013 43293 27073
rect 41126 26674 43293 26734
rect 27648 26590 27714 26593
rect 37048 26590 37118 26595
rect 27648 26588 37053 26590
rect 27648 26532 27653 26588
rect 27709 26532 37053 26588
rect 27648 26530 37053 26532
rect 37113 26530 37118 26590
rect 27648 26527 27714 26530
rect 37048 26525 37118 26530
rect 23123 26451 23189 26454
rect 37692 26451 37762 26456
rect 23123 26449 37697 26451
rect 23123 26393 23128 26449
rect 23184 26393 37697 26449
rect 23123 26391 37697 26393
rect 37757 26391 37762 26451
rect 23123 26388 23189 26391
rect 37692 26386 37762 26391
rect 21142 26295 21208 26298
rect 38336 26295 38406 26300
rect 21142 26293 38341 26295
rect 21142 26237 21147 26293
rect 21203 26237 38341 26293
rect 21142 26235 38341 26237
rect 38401 26235 38406 26295
rect 21142 26232 21208 26235
rect 38336 26230 38406 26235
rect 19894 26133 19964 26138
rect 30478 26133 30544 26136
rect 19894 26073 19899 26133
rect 19959 26131 30544 26133
rect 19959 26075 30483 26131
rect 30539 26075 30544 26131
rect 19959 26073 30544 26075
rect 19894 26068 19964 26073
rect 30478 26070 30544 26073
rect 31034 26126 31104 26131
rect 38068 26126 38134 26129
rect 31034 26066 31039 26126
rect 31099 26124 38134 26126
rect 31099 26068 38073 26124
rect 38129 26068 38134 26124
rect 31099 26066 38134 26068
rect 31034 26061 31104 26066
rect 38068 26063 38134 26066
rect 41261 25137 41419 25142
rect 41261 24989 41266 25137
rect 41414 24989 42463 25137
rect 42611 24989 42617 25137
rect 41261 24984 41419 24989
rect 41169 24425 41429 24430
rect 41169 24175 41174 24425
rect 41424 24175 42057 24425
rect 42307 24175 42313 24425
rect 41169 24170 41429 24175
rect 41153 24091 41261 24096
rect 41153 23993 41158 24091
rect 41256 23993 42933 24091
rect 43031 23993 43037 24091
rect 41153 23988 41261 23993
rect 38217 23859 38291 23864
rect 38217 23795 38222 23859
rect 38286 23795 43293 23859
rect 38217 23790 38291 23795
rect 14073 23704 14147 23709
rect 14955 23704 15021 23705
rect 14073 23640 14078 23704
rect 14142 23700 15021 23704
rect 14142 23644 14960 23700
rect 15016 23644 15021 23700
rect 14142 23640 15021 23644
rect 14073 23635 14147 23640
rect 14955 23639 15021 23640
rect 41079 23611 41445 23616
rect 41079 23255 41084 23611
rect 41440 23255 42470 23611
rect 42826 23255 42832 23611
rect 41079 23250 41445 23255
rect 41219 22691 41479 22696
rect 41219 22441 41224 22691
rect 41474 22441 42015 22691
rect 42265 22441 42271 22691
rect 41219 22436 41479 22441
rect 41611 22357 41721 22362
rect 41611 22257 41616 22357
rect 41716 22257 42988 22357
rect 43088 22257 43094 22357
rect 41611 22252 41721 22257
rect 41040 21877 41360 21882
rect 41040 21567 41045 21877
rect 41355 21567 42503 21877
rect 42813 21567 42819 21877
rect 41040 21562 41360 21567
rect 15157 4251 15227 4256
rect 19896 4251 19962 4254
rect 15157 4191 15162 4251
rect 15222 4249 19962 4251
rect 15222 4193 19901 4249
rect 19957 4193 19962 4249
rect 15222 4191 19962 4193
rect 15157 4186 15227 4191
rect 19896 4188 19962 4191
rect 19645 3696 19715 3701
rect 18622 3636 19650 3696
rect 19710 3636 19715 3696
rect 19645 3631 19715 3636
rect 488 -110 898 -105
rect 488 -207 493 -110
rect -1604 -213 493 -207
rect -1604 -601 -218 -213
rect 170 -510 493 -213
rect 893 -207 898 -110
rect 893 -213 43293 -207
rect 893 -510 41519 -213
rect 170 -601 41519 -510
rect 41907 -601 43293 -213
rect -1604 -607 43293 -601
rect -1604 -673 43293 -667
rect -1604 -1061 -678 -673
rect -290 -707 41979 -673
rect -290 -1039 28 -707
rect 383 -1039 41979 -707
rect -290 -1061 41979 -1039
rect 42367 -1061 43293 -673
rect -1604 -1067 43293 -1061
rect -1604 -1133 43293 -1127
rect -1604 -1521 -1138 -1133
rect -750 -1521 42439 -1133
rect 42827 -1521 43293 -1133
rect -1604 -1527 43293 -1521
rect -1604 -1593 43293 -1587
rect -1604 -1981 -1598 -1593
rect -1210 -1981 42899 -1593
rect 43287 -1981 43293 -1593
rect -1604 -1987 43293 -1981
<< via3 >>
rect -1598 40888 -1210 41276
rect 34162 40930 34480 41248
rect 42899 40888 43287 41276
rect -1138 40428 -750 40816
rect 34822 40454 35140 40772
rect 42439 40428 42827 40816
rect -678 39968 -290 40356
rect 41979 39968 42367 40356
rect -218 39508 170 39896
rect 41519 39508 41907 39896
rect 42463 24989 42611 25137
rect 42057 24175 42307 24425
rect 42933 23993 43031 24091
rect 42470 23255 42826 23611
rect 42015 22441 42265 22691
rect 42988 22257 43088 22357
rect 42503 21567 42813 21877
rect -218 -601 170 -213
rect 41519 -601 41907 -213
rect -678 -1061 -290 -673
rect 41979 -1061 42367 -673
rect -1138 -1521 -750 -1133
rect 42439 -1521 42827 -1133
rect -1598 -1981 -1210 -1593
rect 42899 -1981 43287 -1593
<< metal4 >>
rect -1604 41276 -1204 41283
rect -1604 40888 -1598 41276
rect -1210 40888 -1204 41276
rect -1604 -1593 -1204 40888
rect -1604 -1981 -1598 -1593
rect -1210 -1981 -1204 -1593
rect -1604 -1987 -1204 -1981
rect -1144 40816 -744 41283
rect -1144 40428 -1138 40816
rect -750 40428 -744 40816
rect -1144 -1133 -744 40428
rect -1144 -1521 -1138 -1133
rect -750 -1521 -744 -1133
rect -1144 -1987 -744 -1521
rect -684 40356 -284 41283
rect -684 39968 -678 40356
rect -290 39968 -284 40356
rect -684 -673 -284 39968
rect -684 -1061 -678 -673
rect -290 -1061 -284 -673
rect -684 -1987 -284 -1061
rect -224 39896 176 41283
rect -224 39508 -218 39896
rect 170 39508 176 39896
rect -224 7639 176 39508
rect 34161 41248 34481 41249
rect 34161 40930 34162 41248
rect 34480 40930 34481 41248
rect 34161 36862 34481 40930
rect 34821 40772 35141 40773
rect 34821 40454 34822 40772
rect 35140 40454 35141 40772
rect 34821 36775 35141 40454
rect 41513 39896 41913 41283
rect 41513 39508 41519 39896
rect 41907 39508 41913 39896
rect -224 7237 180 7639
rect -224 -213 176 7237
rect -224 -601 -218 -213
rect 170 -601 176 -213
rect -224 -1987 176 -601
rect 41513 -213 41913 39508
rect 41513 -601 41519 -213
rect 41907 -601 41913 -213
rect 41513 -1987 41913 -601
rect 41973 40356 42373 41283
rect 41973 39968 41979 40356
rect 42367 39968 42373 40356
rect 41973 24425 42373 39968
rect 41973 24175 42057 24425
rect 42307 24175 42373 24425
rect 41973 22691 42373 24175
rect 41973 22441 42015 22691
rect 42265 22441 42373 22691
rect 41973 -673 42373 22441
rect 41973 -1061 41979 -673
rect 42367 -1061 42373 -673
rect 41973 -1987 42373 -1061
rect 42433 40816 42833 41283
rect 42433 40428 42439 40816
rect 42827 40428 42833 40816
rect 42433 25137 42833 40428
rect 42433 24989 42463 25137
rect 42611 24989 42833 25137
rect 42433 23611 42833 24989
rect 42433 23255 42470 23611
rect 42826 23255 42833 23611
rect 42433 21877 42833 23255
rect 42433 21567 42503 21877
rect 42813 21567 42833 21877
rect 42433 -1133 42833 21567
rect 42433 -1521 42439 -1133
rect 42827 -1521 42833 -1133
rect 42433 -1987 42833 -1521
rect 42893 41276 43293 41283
rect 42893 40888 42899 41276
rect 43287 40888 43293 41276
rect 42893 24091 43293 40888
rect 42893 23993 42933 24091
rect 43031 23993 43293 24091
rect 42893 22357 43293 23993
rect 42893 22257 42988 22357
rect 43088 22257 43293 22357
rect 42893 -1593 43293 22257
rect 42893 -1981 42899 -1593
rect 43287 -1981 43293 -1593
rect 42893 -1987 43293 -1981
use por_ana  por_ana_0
timestamp 1712980491
transform 1 0 29373 0 1 25849
box -29373 -25849 13304 13900
use por_dig  por_dig_0
timestamp 1712980491
transform 1 0 29953 0 1 25790
box 0 0 11540 13684
<< labels >>
flabel metal3 1723 -1527 1723 -1527 0 FreeSans 1600 0 0 0 dvss
port 6 nsew
flabel metal3 1723 -1987 1723 -1987 0 FreeSans 1600 0 0 0 dvdd
port 4 nsew
flabel metal3 1723 -607 1723 -607 0 FreeSans 1600 0 0 0 avss
port 2 nsew
flabel metal3 1723 -1067 1723 -1067 0 FreeSans 1600 0 0 0 avdd
port 1 nsew
flabel metal3 43093 27013 43293 27073 0 FreeSans 1600 0 0 0 otrip[1]
port 7 nsew
flabel metal3 43093 27409 43293 27469 0 FreeSans 1600 0 0 0 otrip[0]
port 8 nsew
flabel metal3 43093 26674 43293 26734 0 FreeSans 1600 0 0 0 otrip[2]
port 9 nsew
flabel metal2 s 30421 41082 30481 41282 0 FreeSans 1600 90 0 0 force_ena_rc_osc
port 11 nsew
flabel metal2 s 30879 41082 30939 41282 0 FreeSans 1600 90 0 0 force_pdn
port 12 nsew
flabel metal2 s 29921 41082 29981 41282 0 FreeSans 1600 90 0 0 force_dis_rc_osc
port 13 nsew
flabel metal2 s 29342 41082 29402 41282 0 FreeSans 1600 90 0 0 por_timed_out
port 14 nsew
flabel metal2 s 28854 41082 28914 41282 0 FreeSans 1600 90 0 0 osc_ck
port 15 nsew
flabel metal3 s 43093 33308 43293 33368 0 FreeSans 1600 0 0 0 startup_timed_out
port 17 nsew
flabel metal3 s 43093 31948 43293 32008 0 FreeSans 1600 0 0 0 force_short_oneshot
port 18 nsew
flabel metal2 s 26775 41082 26841 41282 0 FreeSans 1600 90 0 0 por
port 19 nsew
flabel metal2 s 26348 41082 26414 41282 0 FreeSans 1600 90 0 0 dcomp
port 20 nsew
flabel metal2 s 12255 41082 12321 41282 0 FreeSans 1600 90 0 0 itest
port 21 nsew
flabel metal2 s 10871 41082 10935 41282 0 FreeSans 1600 90 0 0 vbg_1v2
port 22 nsew
flabel metal3 s 43093 23795 43293 23859 0 FreeSans 1600 0 0 0 isrc_sel
port 23 nsew
flabel metal2 s 14956 41082 15020 41282 0 FreeSans 1600 90 0 0 ibg_200n
port 24 nsew
flabel metal2 s 21267 41082 21331 41282 0 FreeSans 1600 90 0 0 porb_h
port 25 nsew
flabel metal2 s 27432 41082 27496 41282 0 FreeSans 1600 90 0 0 porb
port 26 nsew
flabel metal3 s -1604 32510 -1404 32570 0 FreeSans 1600 0 0 0 vin
port 27 nsew
flabel metal3 s 43093 27737 43293 27797 0 FreeSans 1600 0 0 0 pwup_filt
port 28 nsew
<< end >>
