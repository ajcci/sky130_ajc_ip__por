* XSpice netlist created from SPICE and liberty sources by spi2xspice.py
* NGSPICE file created from por_dig.ext - technology: sky130A
* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt por_dig a_VGND a_VPWR a_force_dis_rc_osc a_force_ena_rc_osc a_force_pdn a_force_pdnb a_force_short_oneshot a_osc_ck a_osc_ena a_otrip_0_ a_otrip_1_ a_otrip_2_ a_otrip_decoded_0_ a_otrip_decoded_1_ a_otrip_decoded_2_ a_otrip_decoded_3_ a_otrip_decoded_4_ a_otrip_decoded_5_ a_otrip_decoded_6_ a_otrip_decoded_7_ a_por_timed_out a_por_unbuf a_pwup_filt a_startup_timed_out
A_131_ _010_ clknet_1_0__leaf_osc_ck NULL ~net24 cnt_por\_5\_ NULL ddflop
A_062_ [cnt_por\_5\_ cnt_por\_4\_ cnt_por\_7\_ cnt_por\_6\_] _035_ d_lut_sky130_fd_sc_hd__nand4_1
A_114_ [_024_ _025_ _047_] _012_ d_lut_sky130_fd_sc_hd__a21o_1
Aoutput20 [net20] por_unbuf d_lut_sky130_fd_sc_hd__buf_2
A_130_ _009_ clknet_1_1__leaf_osc_ck NULL ~net24 cnt_por\_4\_ NULL ddflop
A_061_ [cnt_por\_1\_ cnt_por\_0\_ cnt_por\_3\_ cnt_por\_2\_] _034_ d_lut_sky130_fd_sc_hd__nand4_2
A_113_ [cnt_por\_7\_ cnt_por\_6\_ net22 _019_] _025_ d_lut_sky130_fd_sc_hd__nand4_1
Aoutput21 [net21] startup_timed_out d_lut_sky130_fd_sc_hd__buf_2
Aoutput10 [net10] osc_ena d_lut_sky130_fd_sc_hd__buf_2
A_060_ [cnt_por\_1\_ cnt_por\_0\_ cnt_por\_3\_ cnt_por\_2\_] _033_ d_lut_sky130_fd_sc_hd__and4_1
A_112_ [cnt_por\_6\_ net22 _019_ cnt_por\_7\_] _024_ d_lut_sky130_fd_sc_hd__a31o_1
Aoutput11 [net11] otrip_decoded_0_ d_lut_sky130_fd_sc_hd__buf_2
Aoutput9 [net9] force_pdnb d_lut_sky130_fd_sc_hd__buf_2
A_111_ [_022_ _023_ _048_] _011_ d_lut_sky130_fd_sc_hd__o21ai_1
Aoutput12 [net12] otrip_decoded_1_ d_lut_sky130_fd_sc_hd__buf_2
A_110_ [cnt_por\_6\_ net22 _019_] _023_ d_lut_sky130_fd_sc_hd__and3_1
Aoutput13 [net13] otrip_decoded_2_ d_lut_sky130_fd_sc_hd__buf_2
Aoutput14 [net14] otrip_decoded_3_ d_lut_sky130_fd_sc_hd__buf_2
A_099_ [cnt_por\_1\_ cnt_por\_0\_ cnt_por\_2\_ net20 cnt_por\_3\_] _053_ d_lut_sky130_fd_sc_hd__a41o_1
Aoutput15 [net15] otrip_decoded_4_ d_lut_sky130_fd_sc_hd__buf_2
A_098_ [_051_ _052_ _047_] _007_ d_lut_sky130_fd_sc_hd__a21o_1
Aoutput16 [net16] otrip_decoded_5_ d_lut_sky130_fd_sc_hd__buf_2
A_097_ [cnt_por\_1\_ cnt_por\_0\_ net23 cnt_por\_2\_] _052_ d_lut_sky130_fd_sc_hd__a31o_1
Aoutput17 [net17] otrip_decoded_6_ d_lut_sky130_fd_sc_hd__buf_2
A_137__260 net26 done
A_137__261 _137__26/LO dzero
A_096_ [cnt_por\_1\_ cnt_por\_0\_ cnt_por\_2\_ net23] _051_ d_lut_sky130_fd_sc_hd__nand4_1
A_079_ [cnt_st\_1\_ cnt_st\_0\_] _040_ d_lut_sky130_fd_sc_hd__or2_1
Aoutput18 [net18] otrip_decoded_7_ d_lut_sky130_fd_sc_hd__buf_2
A_095_ [_049_ _050_ _048_] _006_ d_lut_sky130_fd_sc_hd__o21ai_1
A_078_ [net31 _039_] _000_ d_lut_sky130_fd_sc_hd__nand2_1
Aoutput19 [net19] por_timed_out d_lut_sky130_fd_sc_hd__buf_2
A_094_ [cnt_por\_1\_ cnt_por\_0\_ net23] _050_ d_lut_sky130_fd_sc_hd__and3_1
A_129_ _008_ clknet_1_1__leaf_osc_ck NULL ~net24 cnt_por\_3\_ NULL ddflop
A_077_ [net4 net21] _039_ d_lut_sky130_fd_sc_hd__nor2_1
A_093_ [cnt_por\_0\_ net23 cnt_por\_1\_] _049_ d_lut_sky130_fd_sc_hd__a21oi_1
Afanout22 [net23] net22 d_lut_sky130_fd_sc_hd__clkbuf_2
Ainput1 [force_dis_rc_osc] net1 d_lut_sky130_fd_sc_hd__clkbuf_1
A_076_ [_034_ _035_ _037_ _031_ cnt_st\_4\_] net20 d_lut_sky130_fd_sc_hd__o311a_1
A_128_ _007_ clknet_1_1__leaf_osc_ck NULL ~net24 cnt_por\_2\_ NULL ddflop
A_059_ [cnt_st\_4\_ _031_] net21 d_lut_sky130_fd_sc_hd__and2_1
Afanout23 [net20] net23 d_lut_sky130_fd_sc_hd__clkbuf_2
A_092_ [net4 net22] _048_ d_lut_sky130_fd_sc_hd__nand2_1
Ainput2 [force_ena_rc_osc] net2 d_lut_sky130_fd_sc_hd__clkbuf_1
A_127_ _006_ clknet_1_1__leaf_osc_ck NULL ~net24 cnt_por\_1\_ NULL ddflop
A_058_ [_031_] _032_ d_lut_sky130_fd_sc_hd__inv_2
A_075_ [net2 _038_] net10 d_lut_sky130_fd_sc_hd__nand2b_1
Afanout24 [net27] net24 d_lut_sky130_fd_sc_hd__clkbuf_4
A_091_ [net4 net22] _047_ d_lut_sky130_fd_sc_hd__and2_1
A_074_ [net1 net19 net8] _038_ d_lut_sky130_fd_sc_hd__or3b_1
Ainput3 [force_pdn] net3 d_lut_sky130_fd_sc_hd__clkbuf_1
A_126_ _005_ clknet_1_1__leaf_osc_ck NULL ~net24 cnt_por\_0\_ NULL ddflop
A_057_ [cnt_st\_1\_ cnt_st\_0\_ cnt_st\_3\_ cnt_st\_2\_] _031_ d_lut_sky130_fd_sc_hd__and4_1
A_109_ [net22 _019_ cnt_por\_6\_] _022_ d_lut_sky130_fd_sc_hd__a21oi_1
Afanout25 [net27] net25 d_lut_sky130_fd_sc_hd__clkbuf_2
A_090_ [net23 _046_ cnt_por\_0\_] _005_ d_lut_sky130_fd_sc_hd__mux2_1
Ainput4 [force_short_oneshot] net4 d_lut_sky130_fd_sc_hd__buf_2
A_056_ [cnt_st\_1\_ cnt_st\_0\_ cnt_st\_2\_] _030_ d_lut_sky130_fd_sc_hd__and3_1
A_125_ _004_ clknet_1_0__leaf_osc_ck NULL ~net25 cnt_st\_4\_ NULL ddflop
A_073_ [net7 net6 net5] net18 d_lut_sky130_fd_sc_hd__and3_1
A_108_ [_020_ _021_ _047_] _010_ d_lut_sky130_fd_sc_hd__a21o_1
Ainput5 [otrip_0_] net5 d_lut_sky130_fd_sc_hd__dlymetal6s2s_1
A_072_ [net5 net6 net7] net17 d_lut_sky130_fd_sc_hd__and3b_1
A_055_ [cnt_st\_1\_ cnt_st\_0\_] _029_ d_lut_sky130_fd_sc_hd__nand2_1
A_124_ _003_ clknet_1_0__leaf_osc_ck NULL ~net25 cnt_st\_3\_ NULL ddflop
A_107_ [cnt_por\_4\_ _033_ net22 cnt_por\_5\_] _021_ d_lut_sky130_fd_sc_hd__a31o_1
Ainput6 [otrip_1_] net6 d_lut_sky130_fd_sc_hd__dlymetal6s2s_1
A_071_ [net6 net5 net7] net16 d_lut_sky130_fd_sc_hd__and3b_1
A_106_ [net22 _019_] _020_ d_lut_sky130_fd_sc_hd__nand2_1
A_123_ _002_ clknet_1_1__leaf_osc_ck NULL ~net24 cnt_st\_2\_ NULL ddflop
A_054_ [net3] net9 d_lut_sky130_fd_sc_hd__inv_2
Ainput7 [otrip_2_] net7 d_lut_sky130_fd_sc_hd__dlymetal6s2s_1
A_070_ [net6 net5 net7] net15 d_lut_sky130_fd_sc_hd__nor3b_1
A_122_ _001_ clknet_1_1__leaf_osc_ck NULL ~net25 cnt_st\_1\_ NULL ddflop
A_105_ [cnt_por\_5\_ cnt_por\_4\_ _033_] _019_ d_lut_sky130_fd_sc_hd__and3_1
Aclkbuf_1_1__f_osc_ck [clknet_0_osc_ck] clknet_1_1__leaf_osc_ck d_lut_sky130_fd_sc_hd__clkbuf_16
Ainput8 [pwup_filt] net8 d_lut_sky130_fd_sc_hd__buf_1
A_121_ _000_ clknet_1_1__leaf_osc_ck NULL ~net25 cnt_st\_0\_ NULL ddflop
A_104_ [_017_ _018_ _048_] _009_ d_lut_sky130_fd_sc_hd__o21ai_1
A_120_ [net29 _028_] _015_ d_lut_sky130_fd_sc_hd__xor2_1
A_103_ [_033_ net23 cnt_por\_4\_] _018_ d_lut_sky130_fd_sc_hd__a21oi_1
Ahold1 [cnt_rsb] net27 d_lut_sky130_fd_sc_hd__dlygate4sd3_1
Aclkbuf_0_osc_ck [osc_ck] clknet_0_osc_ck d_lut_sky130_fd_sc_hd__clkbuf_16
A_102_ [cnt_por\_4\_ _033_ net23] _017_ d_lut_sky130_fd_sc_hd__and3_1
Ahold2 [cnt_rsb_stg1] net28 d_lut_sky130_fd_sc_hd__dlygate4sd3_1
A_101_ [_053_ _016_ _047_] _008_ d_lut_sky130_fd_sc_hd__a21o_1
Ahold3 [cnt_por\_10\_] net29 d_lut_sky130_fd_sc_hd__dlygate4sd3_1
A_100_ [_033_ net20] _016_ d_lut_sky130_fd_sc_hd__nand2_1
Ahold4 [cnt_por\_9\_] net30 d_lut_sky130_fd_sc_hd__dlygate4sd3_1
Ahold5 [cnt_st\_0\_] net31 d_lut_sky130_fd_sc_hd__dlygate4sd3_1
A_089_ [net4 net23] _046_ d_lut_sky130_fd_sc_hd__nand2b_1
Ahold6 [cnt_por\_8\_] net32 d_lut_sky130_fd_sc_hd__dlygate4sd3_1
A_088_ [net34 _042_ _045_] _004_ d_lut_sky130_fd_sc_hd__a21bo_1
Ahold7 [cnt_st\_2\_] net33 d_lut_sky130_fd_sc_hd__dlygate4sd3_1
Ahold8 [cnt_st\_4\_] net34 d_lut_sky130_fd_sc_hd__dlygate4sd3_1
A_087_ [cnt_st\_4\_ _042_ _032_] _045_ d_lut_sky130_fd_sc_hd__o21a_1
Aclkbuf_1_0__f_osc_ck [clknet_0_osc_ck] clknet_1_0__leaf_osc_ck d_lut_sky130_fd_sc_hd__clkbuf_16
A_086_ [net34 _032_ _044_] _003_ d_lut_sky130_fd_sc_hd__o21a_1
A_138_ net28 clknet_1_0__leaf_osc_ck NULL ~net8 cnt_rsb NULL ddflop
A_069_ [net7 net6 net5] net14 d_lut_sky130_fd_sc_hd__and3b_1
A_085_ [_042_ _043_ _030_] _044_ d_lut_sky130_fd_sc_hd__a21o_1
A_137_ net26 clknet_1_0__leaf_osc_ck NULL ~net8 cnt_rsb_stg1 NULL ddflop
A_068_ [net7 net5 net6] net13 d_lut_sky130_fd_sc_hd__nor3b_1
A_136_ _015_ clknet_1_0__leaf_osc_ck NULL ~net25 cnt_por\_10\_ NULL ddflop
A_084_ [cnt_st\_3\_ net4] _043_ d_lut_sky130_fd_sc_hd__or2_1
A_067_ [net7 net6 net5] net12 d_lut_sky130_fd_sc_hd__nor3b_1
A_119_ [net30 _027_] _014_ d_lut_sky130_fd_sc_hd__xor2_1
A_083_ [cnt_st\_3\_ net4] _042_ d_lut_sky130_fd_sc_hd__nand2_1
A_118_ [net4 _036_ net23 cnt_por\_8\_ cnt_por\_9\_] _028_ d_lut_sky130_fd_sc_hd__o2111a_1
A_066_ [net7 net6 net5] net11 d_lut_sky130_fd_sc_hd__nor3_1
A_135_ _014_ clknet_1_0__leaf_osc_ck NULL ~net25 cnt_por\_9\_ NULL ddflop
A_082_ [_030_ _041_ _039_] _002_ d_lut_sky130_fd_sc_hd__o21ai_1
A_065_ [_034_ _035_ _037_] net19 d_lut_sky130_fd_sc_hd__nor3_1
A_134_ _013_ clknet_1_0__leaf_osc_ck NULL ~net24 cnt_por\_8\_ NULL ddflop
A_117_ [net32 _026_] _013_ d_lut_sky130_fd_sc_hd__xnor2_1
A_081_ [cnt_st\_1\_ cnt_st\_0\_ net33] _041_ d_lut_sky130_fd_sc_hd__a21oi_1
A_133_ _012_ clknet_1_0__leaf_osc_ck NULL ~net24 cnt_por\_7\_ NULL ddflop
A_064_ [cnt_por\_9\_ cnt_por\_8\_ cnt_por\_10\_] _037_ d_lut_sky130_fd_sc_hd__nand3_1
A_116_ [net4 _036_ net22 cnt_por\_8\_] _027_ d_lut_sky130_fd_sc_hd__o211a_1
A_132_ _011_ clknet_1_1__leaf_osc_ck NULL ~net24 cnt_por\_6\_ NULL ddflop
A_080_ [_029_ _040_ net21 net4] _001_ d_lut_sky130_fd_sc_hd__a211o_1
A_063_ [_034_ _035_] _036_ d_lut_sky130_fd_sc_hd__nor2_1
A_115_ [net4 _036_ net22] _026_ d_lut_sky130_fd_sc_hd__o21ai_1

.model todig_1v8 adc_bridge(in_high=1.2 in_low=0.6 rise_delay=10n fall_delay=10n)
.model toana_1v8 dac_bridge(out_high=1.8 out_low=0)

.model ddflop d_dff(ic=0 rise_delay=1n fall_delay=1n)
.model dlatch d_dlatch(ic=0 rise_delay=1n fall_delay=1n)
.model dzero d_pulldown(load=1p)
.model done d_pullup(load=1p)

AA2D1 [a_VGND] [VGND] todig_1v8
AA2D2 [a_VPWR] [VPWR] todig_1v8
AA2D3 [a_force_dis_rc_osc] [force_dis_rc_osc] todig_1v8
AA2D4 [a_force_ena_rc_osc] [force_ena_rc_osc] todig_1v8
AA2D5 [a_force_pdn] [force_pdn] todig_1v8
AD2A1 [force_pdnb] [a_force_pdnb] toana_1v8
AA2D6 [a_force_short_oneshot] [force_short_oneshot] todig_1v8
AA2D7 [a_osc_ck] [osc_ck] todig_1v8
AD2A2 [osc_ena] [a_osc_ena] toana_1v8
AA2D8 [a_otrip_0_] [otrip_0_] todig_1v8
AA2D9 [a_otrip_1_] [otrip_1_] todig_1v8
AA2D10 [a_otrip_2_] [otrip_2_] todig_1v8
AD2A3 [otrip_decoded_0_] [a_otrip_decoded_0_] toana_1v8
AD2A4 [otrip_decoded_1_] [a_otrip_decoded_1_] toana_1v8
AD2A5 [otrip_decoded_2_] [a_otrip_decoded_2_] toana_1v8
AD2A6 [otrip_decoded_3_] [a_otrip_decoded_3_] toana_1v8
AD2A7 [otrip_decoded_4_] [a_otrip_decoded_4_] toana_1v8
AD2A8 [otrip_decoded_5_] [a_otrip_decoded_5_] toana_1v8
AD2A9 [otrip_decoded_6_] [a_otrip_decoded_6_] toana_1v8
AD2A10 [otrip_decoded_7_] [a_otrip_decoded_7_] toana_1v8
AD2A11 [por_timed_out] [a_por_timed_out] toana_1v8
AD2A12 [por_unbuf] [a_por_unbuf] toana_1v8
AA2D11 [a_pwup_filt] [pwup_filt] todig_1v8
AD2A13 [startup_timed_out] [a_startup_timed_out] toana_1v8

.ends


* sky130_fd_sc_hd__tapvpwrvgnd_1 (no function)
* sky130_ef_sc_hd__decap_12 (no function)
* sky130_fd_sc_hd__dfrtp_1 IQ
* sky130_fd_sc_hd__decap_3 (no function)
* sky130_fd_sc_hd__nand4_1 (!A) | (!B) | (!C) | (!D)
.model d_lut_sky130_fd_sc_hd__nand4_1 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "1111111111111110")
* sky130_fd_sc_hd__decap_8 (no function)
* sky130_fd_sc_hd__a21o_1 (A1&A2) | (B1)
.model d_lut_sky130_fd_sc_hd__a21o_1 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "00011111")
* sky130_fd_sc_hd__buf_2 (A)
.model d_lut_sky130_fd_sc_hd__buf_2 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "01")
* sky130_fd_sc_hd__nand4_2 (!A) | (!B) | (!C) | (!D)
.model d_lut_sky130_fd_sc_hd__nand4_2 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "1111111111111110")
* sky130_fd_sc_hd__fill_1 (no function)
* sky130_fd_sc_hd__and4_1 (A&B&C&D)
.model d_lut_sky130_fd_sc_hd__and4_1 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "0000000000000001")
* sky130_fd_sc_hd__fill_2 (no function)
* sky130_fd_sc_hd__a31o_1 (A1&A2&A3) | (B1)
.model d_lut_sky130_fd_sc_hd__a31o_1 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "0000000111111111")
* sky130_fd_sc_hd__o21ai_1 (!A1&!A2) | (!B1)
.model d_lut_sky130_fd_sc_hd__o21ai_1 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "11111000")
* sky130_fd_sc_hd__and3_1 (A&B&C)
.model d_lut_sky130_fd_sc_hd__and3_1 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "00000001")
* sky130_fd_sc_hd__decap_6 (no function)
* sky130_fd_sc_hd__a41o_1 (A1&A2&A3&A4) | (B1)
.model d_lut_sky130_fd_sc_hd__a41o_1 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "00000000000000011111111111111111")
* sky130_fd_sc_hd__conb_1 1
* sky130_fd_sc_hd__or2_1 (A) | (B)
.model d_lut_sky130_fd_sc_hd__or2_1 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "0111")
* sky130_fd_sc_hd__nand2_1 (!A) | (!B)
.model d_lut_sky130_fd_sc_hd__nand2_1 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "1110")
* sky130_fd_sc_hd__decap_4 (no function)
* sky130_fd_sc_hd__nor2_1 (!A&!B)
.model d_lut_sky130_fd_sc_hd__nor2_1 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "1000")
* sky130_fd_sc_hd__a21oi_1 (!A1&!B1) | (!A2&!B1)
.model d_lut_sky130_fd_sc_hd__a21oi_1 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "11100000")
* sky130_fd_sc_hd__clkbuf_2 (A)
.model d_lut_sky130_fd_sc_hd__clkbuf_2 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "01")
* sky130_fd_sc_hd__clkbuf_1 (A)
.model d_lut_sky130_fd_sc_hd__clkbuf_1 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "01")
* sky130_fd_sc_hd__o311a_1 (A1&B1&C1) | (A2&B1&C1) | (A3&B1&C1)
.model d_lut_sky130_fd_sc_hd__o311a_1 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "00000000000000000000000001111111")
* sky130_fd_sc_hd__and2_1 (A&B)
.model d_lut_sky130_fd_sc_hd__and2_1 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "0001")
* sky130_fd_sc_hd__dfrtp_2 IQ
* sky130_fd_sc_hd__inv_2 (!A)
.model d_lut_sky130_fd_sc_hd__inv_2 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "10")
* sky130_fd_sc_hd__nand2b_1 (A_N) | (!B)
.model d_lut_sky130_fd_sc_hd__nand2b_1 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "1101")
* sky130_fd_sc_hd__clkbuf_4 (A)
.model d_lut_sky130_fd_sc_hd__clkbuf_4 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "01")
* sky130_fd_sc_hd__or3b_1 (A) | (B) | (!C_N)
.model d_lut_sky130_fd_sc_hd__or3b_1 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "11110111")
* sky130_fd_sc_hd__dfrtp_4 IQ
* sky130_fd_sc_hd__mux2_1 (A0&!S) | (A1&S)
.model d_lut_sky130_fd_sc_hd__mux2_1 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "01010011")
* sky130_fd_sc_hd__dlymetal6s2s_1 (A)
.model d_lut_sky130_fd_sc_hd__dlymetal6s2s_1 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "01")
* sky130_fd_sc_hd__and3b_1 (!A_N&B&C)
.model d_lut_sky130_fd_sc_hd__and3b_1 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "00000010")
* sky130_fd_sc_hd__nor3b_1 (!A&!B&C_N)
.model d_lut_sky130_fd_sc_hd__nor3b_1 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "00001000")
* sky130_fd_sc_hd__clkbuf_16 (A)
.model d_lut_sky130_fd_sc_hd__clkbuf_16 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "01")
* sky130_fd_sc_hd__buf_1 (A)
.model d_lut_sky130_fd_sc_hd__buf_1 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "01")
* sky130_fd_sc_hd__xor2_1 (A&!B) | (!A&B)
.model d_lut_sky130_fd_sc_hd__xor2_1 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "0110")
* sky130_fd_sc_hd__dlygate4sd3_1 (A)
.model d_lut_sky130_fd_sc_hd__dlygate4sd3_1 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "01")
* sky130_fd_sc_hd__a21bo_1 (A1&A2) | (!B1_N)
.model d_lut_sky130_fd_sc_hd__a21bo_1 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "11110001")
* sky130_fd_sc_hd__o21a_1 (A1&B1) | (A2&B1)
.model d_lut_sky130_fd_sc_hd__o21a_1 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "00000111")
* sky130_fd_sc_hd__o2111a_1 (A1&B1&C1&D1) | (A2&B1&C1&D1)
.model d_lut_sky130_fd_sc_hd__o2111a_1 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "00000000000000000000000000000111")
* sky130_fd_sc_hd__nor3_1 (!A&!B&!C)
.model d_lut_sky130_fd_sc_hd__nor3_1 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "10000000")
* sky130_fd_sc_hd__xnor2_1 (!A&!B) | (A&B)
.model d_lut_sky130_fd_sc_hd__xnor2_1 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "1001")
* sky130_fd_sc_hd__nand3_1 (!A) | (!B) | (!C)
.model d_lut_sky130_fd_sc_hd__nand3_1 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "11111110")
* sky130_fd_sc_hd__o211a_1 (A1&B1&C1) | (A2&B1&C1)
.model d_lut_sky130_fd_sc_hd__o211a_1 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "0000000000000111")
* sky130_fd_sc_hd__a211o_1 (A1&A2) | (B1) | (C1)
.model d_lut_sky130_fd_sc_hd__a211o_1 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "0001111111111111")
.end
