* XSpice netlist created from SPICE and liberty sources by spi2xspice.py
* NGSPICE file created from por_dig.ext - technology: sky130A
* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt por_dig a_VGND a_VPWR a_force_dis_rc_osc a_force_ena_rc_osc a_force_pdn a_force_pdnb a_force_short_oneshot a_osc_ck a_osc_ena a_otrip_0_ a_otrip_1_ a_otrip_2_ a_otrip_decoded_0_ a_otrip_decoded_1_ a_otrip_decoded_2_ a_otrip_decoded_3_ a_otrip_decoded_4_ a_otrip_decoded_5_ a_otrip_decoded_6_ a_otrip_decoded_7_ a_por_timed_out a_por_unbuf a_pwup_filt a_startup_timed_out
A_131_ net29 clknet_1_0__leaf_osc_ck NULL ~net8 cnt_rsb NULL ddflop
A_062_ [net7 net6 net5] net12 d_lut_sky130_fd_sc_hd__nor3b_1
A_114_ net36 clknet_1_0__leaf_osc_ck NULL ~net24 cnt_st\_1\_ NULL ddflop
Aoutput20 [net20] por_unbuf d_lut_sky130_fd_sc_hd__buf_2
A_130_ net27 clknet_1_0__leaf_osc_ck NULL ~net8 cnt_rsb_stg1 NULL ddflop
A_113_ _000_ clknet_1_0__leaf_osc_ck NULL ~net24 cnt_st\_0\_ NULL ddflop
A_061_ [net7 net6 net5] net11 d_lut_sky130_fd_sc_hd__nor3_1
Aoutput21 [net23] startup_timed_out d_lut_sky130_fd_sc_hd__buf_2
Aoutput10 [net10] osc_ena d_lut_sky130_fd_sc_hd__buf_2
A_060_ [net22] net19 d_lut_sky130_fd_sc_hd__inv_2
Ahold10 [cnt_por\_5\_] net37 d_lut_sky130_fd_sc_hd__dlygate4sd3_1
A_112_ [net31 _026_] _016_ d_lut_sky130_fd_sc_hd__xor2_1
Aoutput11 [net11] otrip_decoded_0_ d_lut_sky130_fd_sc_hd__buf_2
Aoutput9 [net9] force_pdnb d_lut_sky130_fd_sc_hd__buf_2
A_111_ [_026_ _027_] _015_ d_lut_sky130_fd_sc_hd__and2b_1
Ahold11 [cnt_por\_1\_] net38 d_lut_sky130_fd_sc_hd__dlygate4sd3_1
Aoutput12 [net12] otrip_decoded_1_ d_lut_sky130_fd_sc_hd__buf_2
A_110_ [cnt_por\_8\_ net23 net22 _024_ net42] _027_ d_lut_sky130_fd_sc_hd__a41o_1
Ahold12 [cnt_por\_7\_] net39 d_lut_sky130_fd_sc_hd__dlygate4sd3_1
Aoutput13 [net13] otrip_decoded_2_ d_lut_sky130_fd_sc_hd__buf_2
Ahold13 [cnt_por\_2\_] net40 d_lut_sky130_fd_sc_hd__dlygate4sd3_1
Aoutput14 [net14] otrip_decoded_3_ d_lut_sky130_fd_sc_hd__buf_2
A_099_ [_034_ _049_] _020_ d_lut_sky130_fd_sc_hd__and2_1
Ahold14 [cnt_st\_2\_] net41 d_lut_sky130_fd_sc_hd__dlygate4sd3_1
Aoutput15 [net15] otrip_decoded_4_ d_lut_sky130_fd_sc_hd__buf_2
A_098_ [cnt_por\_4\_ _049_ cnt_por\_5\_] _019_ d_lut_sky130_fd_sc_hd__a21oi_1
Ahold15 [cnt_por\_9\_] net42 d_lut_sky130_fd_sc_hd__dlygate4sd3_1
Aoutput16 [net16] otrip_decoded_5_ d_lut_sky130_fd_sc_hd__buf_2
A_097_ [net26 _036_ _018_ _017_ net34] _010_ d_lut_sky130_fd_sc_hd__o32a_1
Aoutput17 [net17] otrip_decoded_6_ d_lut_sky130_fd_sc_hd__buf_2
A_096_ [cnt_por\_4\_ _049_] _018_ d_lut_sky130_fd_sc_hd__nand2_1
A_079_ [cnt_st\_3\_ net26 _039_ _040_ _030_] _003_ d_lut_sky130_fd_sc_hd__o311a_1
Aoutput18 [net18] otrip_decoded_7_ d_lut_sky130_fd_sc_hd__buf_2
A_095_ [net33 _048_ _017_] _009_ d_lut_sky130_fd_sc_hd__o21ba_1
Aoutput19 [net19] por_timed_out d_lut_sky130_fd_sc_hd__buf_2
A_078_ [net26 _039_ cnt_st\_3\_] _040_ d_lut_sky130_fd_sc_hd__o21ai_1
A_094_ [net4 _049_ _035_ net21] _017_ d_lut_sky130_fd_sc_hd__o211a_1
A_129_ _016_ clknet_1_0__leaf_osc_ck NULL ~net24 cnt_por\_10\_ NULL ddflop
A_077_ [_038_ _039_ net26] _002_ d_lut_sky130_fd_sc_hd__o21bai_1
A_093_ [cnt_por\_1\_ cnt_por\_0\_ cnt_por\_3\_ cnt_por\_2\_] _049_ d_lut_sky130_fd_sc_hd__and4_1
Afanout22 [_035_] net22 d_lut_sky130_fd_sc_hd__buf_2
A_076_ [cnt_st\_0\_ cnt_st\_1\_ cnt_st\_2\_] _039_ d_lut_sky130_fd_sc_hd__and3_1
Ainput1 [force_dis_rc_osc] net1 d_lut_sky130_fd_sc_hd__clkbuf_1
A_128_ _015_ clknet_1_0__leaf_osc_ck NULL ~net24 cnt_por\_9\_ NULL ddflop
A_059_ [_031_ _032_ _033_ _034_] _035_ d_lut_sky130_fd_sc_hd__or4bb_1
Afanout23 [net21] net23 d_lut_sky130_fd_sc_hd__buf_2
Ainput2 [force_ena_rc_osc] net2 d_lut_sky130_fd_sc_hd__clkbuf_1
A_092_ [cnt_por\_2\_ net21 net22 _045_] _048_ d_lut_sky130_fd_sc_hd__and4_1
A_058_ [cnt_por\_5\_ cnt_por\_4\_] _034_ d_lut_sky130_fd_sc_hd__and2_1
A_127_ _014_ clknet_1_0__leaf_osc_ck NULL ~net24 cnt_por\_8\_ NULL ddflop
A_075_ [cnt_st\_0\_ cnt_st\_1\_ net41] _038_ d_lut_sky130_fd_sc_hd__a21oi_1
Afanout24 [net28] net24 d_lut_sky130_fd_sc_hd__clkbuf_4
A_091_ [_043_ _046_ _047_ _036_ net40] _008_ d_lut_sky130_fd_sc_hd__a32o_1
A_074_ [cnt_st\_0\_ net35 net23 _037_] _001_ d_lut_sky130_fd_sc_hd__a211oi_1
Ainput3 [force_pdn] net3 d_lut_sky130_fd_sc_hd__clkbuf_1
A_057_ [cnt_por\_9\_ cnt_por\_8\_] _033_ d_lut_sky130_fd_sc_hd__and2_1
A_126_ _013_ clknet_1_0__leaf_osc_ck NULL ~net24 cnt_por\_7\_ NULL ddflop
A_109_ [net23 _033_ net22 _024_] _026_ d_lut_sky130_fd_sc_hd__and4_1
Afanout25 [net28] net25 d_lut_sky130_fd_sc_hd__buf_2
A_090_ [cnt_por\_2\_ _045_] _047_ d_lut_sky130_fd_sc_hd__nand2_1
Ainput4 [force_short_oneshot] net4 d_lut_sky130_fd_sc_hd__buf_1
A_125_ _012_ clknet_1_0__leaf_osc_ck NULL ~net24 cnt_por\_6\_ NULL ddflop
A_073_ [cnt_st\_0\_ cnt_st\_1\_ net26] _037_ d_lut_sky130_fd_sc_hd__o21bai_1
A_056_ [cnt_por\_0\_ cnt_por\_3\_ cnt_por\_2\_ cnt_por\_1\_] _032_ d_lut_sky130_fd_sc_hd__or4b_1
A_130__270 net27 done
A_130__271 _130__27/LO dzero
A_108_ [net32 _025_] _014_ d_lut_sky130_fd_sc_hd__xor2_1
Afanout26 [net4] net26 d_lut_sky130_fd_sc_hd__clkbuf_2
Ainput5 [otrip_0_] net5 d_lut_sky130_fd_sc_hd__dlymetal6s2s_1
A_072_ [net26 net23 cnt_st\_0\_] _000_ d_lut_sky130_fd_sc_hd__or3b_1
A_124_ _011_ clknet_1_0__leaf_osc_ck NULL ~net24 cnt_por\_5\_ NULL ddflop
A_055_ [cnt_por\_7\_ cnt_por\_6\_ cnt_por\_10\_] _031_ d_lut_sky130_fd_sc_hd__or3b_1
A_107_ [net39 _023_ _025_] _013_ d_lut_sky130_fd_sc_hd__o21ba_1
A_071_ [_036_] net20 d_lut_sky130_fd_sc_hd__inv_2
Ainput6 [otrip_1_] net6 d_lut_sky130_fd_sc_hd__dlymetal6s2s_1
A_054_ [net23] _030_ d_lut_sky130_fd_sc_hd__inv_2
A_123_ _010_ clknet_1_0__leaf_osc_ck NULL ~net24 cnt_por\_4\_ NULL ddflop
A_106_ [net23 net22 _024_] _025_ d_lut_sky130_fd_sc_hd__and3_1
A_070_ [net23 net22] _036_ d_lut_sky130_fd_sc_hd__nand2_2
Ainput7 [otrip_2_] net7 d_lut_sky130_fd_sc_hd__dlymetal6s2s_1
A_122_ _009_ clknet_1_1__leaf_osc_ck NULL ~net25 cnt_por\_3\_ NULL ddflop
A_053_ [cnt_st\_1\_ _029_ cnt_st\_0\_] net21 d_lut_sky130_fd_sc_hd__and3b_1
A_105_ [cnt_por\_7\_ cnt_por\_6\_ _034_ _049_ net26] _024_ d_lut_sky130_fd_sc_hd__a41o_1
Aclkbuf_1_1__f_osc_ck [clknet_0_osc_ck] clknet_1_1__leaf_osc_ck d_lut_sky130_fd_sc_hd__clkbuf_16
Ainput8 [pwup_filt] net8 d_lut_sky130_fd_sc_hd__buf_1
A_121_ _008_ clknet_1_1__leaf_osc_ck NULL ~net25 cnt_por\_2\_ NULL ddflop
A_104_ [cnt_por\_6\_ net23 net22 _020_] _023_ d_lut_sky130_fd_sc_hd__and4_1
A_052_ [cnt_st\_3\_ cnt_st\_4\_ cnt_st\_5\_ cnt_st\_2\_] _029_ d_lut_sky130_fd_sc_hd__and4bb_1
A_120_ _007_ clknet_1_1__leaf_osc_ck NULL ~net25 cnt_por\_1\_ NULL ddflop
A_051_ [net1] _028_ d_lut_sky130_fd_sc_hd__inv_2
A_103_ [cnt_por\_6\_ _036_ _043_ _022_] _012_ d_lut_sky130_fd_sc_hd__a22o_1
Ahold1 [cnt_rsb] net28 d_lut_sky130_fd_sc_hd__dlygate4sd3_1
A_102_ [cnt_por\_6\_ _020_] _022_ d_lut_sky130_fd_sc_hd__xor2_1
Aclkbuf_0_osc_ck [osc_ck] clknet_0_osc_ck d_lut_sky130_fd_sc_hd__clkbuf_16
A_050_ [net3] net9 d_lut_sky130_fd_sc_hd__inv_2
Ahold2 [cnt_rsb_stg1] net29 d_lut_sky130_fd_sc_hd__dlygate4sd3_1
A_101_ [_043_ _021_ net37 net20] _011_ d_lut_sky130_fd_sc_hd__o2bb2a_1
Ahold3 [cnt_st\_5\_] net30 d_lut_sky130_fd_sc_hd__dlygate4sd3_1
A_100_ [_019_ _020_] _021_ d_lut_sky130_fd_sc_hd__or2_1
Ahold4 [cnt_por\_10\_] net31 d_lut_sky130_fd_sc_hd__dlygate4sd3_1
Ahold5 [cnt_por\_8\_] net32 d_lut_sky130_fd_sc_hd__dlygate4sd3_1
A_089_ [cnt_por\_2\_ _045_] _046_ d_lut_sky130_fd_sc_hd__or2_1
Ahold6 [cnt_por\_3\_] net33 d_lut_sky130_fd_sc_hd__dlygate4sd3_1
A_088_ [_043_ _045_ _044_ net38] _007_ d_lut_sky130_fd_sc_hd__o2bb2a_1
Ahold7 [cnt_por\_4\_] net34 d_lut_sky130_fd_sc_hd__dlygate4sd3_1
A_087_ [cnt_por\_1\_ cnt_por\_0\_] _045_ d_lut_sky130_fd_sc_hd__and2_1
Ahold8 [cnt_st\_1\_] net35 d_lut_sky130_fd_sc_hd__dlygate4sd3_1
Aclkbuf_1_0__f_osc_ck [clknet_0_osc_ck] clknet_1_0__leaf_osc_ck d_lut_sky130_fd_sc_hd__clkbuf_16
A_086_ [cnt_por\_0\_ net26 net21 net22] _044_ d_lut_sky130_fd_sc_hd__o211a_1
Ahold9 [_001_] net36 d_lut_sky130_fd_sc_hd__dlygate4sd3_1
A_069_ [net8 _028_ net22 net2] net10 d_lut_sky130_fd_sc_hd__a31o_1
A_085_ [_043_ _036_ cnt_por\_0\_] _006_ d_lut_sky130_fd_sc_hd__mux2_1
A_068_ [net7 net6 net5] net18 d_lut_sky130_fd_sc_hd__and3_1
A_084_ [net26 net23 net22] _043_ d_lut_sky130_fd_sc_hd__and3b_1
A_067_ [net5 net6 net7] net17 d_lut_sky130_fd_sc_hd__and3b_1
A_119_ _006_ clknet_1_1__leaf_osc_ck NULL ~net24 cnt_por\_0\_ NULL ddflop
A_083_ [net30 _041_] _005_ d_lut_sky130_fd_sc_hd__xor2_1
A_118_ _005_ clknet_1_1__leaf_osc_ck NULL ~net25 cnt_st\_5\_ NULL ddflop
A_066_ [net6 net5 net7] net16 d_lut_sky130_fd_sc_hd__and3b_1
A_082_ [_041_ _042_] _004_ d_lut_sky130_fd_sc_hd__nor2_1
A_065_ [net6 net5 net7] net15 d_lut_sky130_fd_sc_hd__nor3b_1
A_117_ _004_ clknet_1_1__leaf_osc_ck NULL ~net25 cnt_st\_4\_ NULL ddflop
A_081_ [cnt_st\_4\_ _040_] _042_ d_lut_sky130_fd_sc_hd__and2b_1
A_064_ [net7 net6 net5] net14 d_lut_sky130_fd_sc_hd__and3b_1
A_116_ _003_ clknet_1_1__leaf_osc_ck NULL ~net25 cnt_st\_3\_ NULL ddflop
A_080_ [net26 _039_ cnt_st\_3\_ cnt_st\_4\_] _041_ d_lut_sky130_fd_sc_hd__o211a_1
A_063_ [net7 net5 net6] net13 d_lut_sky130_fd_sc_hd__nor3b_1
A_115_ _002_ clknet_1_0__leaf_osc_ck NULL ~net25 cnt_st\_2\_ NULL ddflop

.model todig_1v8 adc_bridge(in_high=1.2 in_low=0.6 rise_delay=10n fall_delay=10n)
.model toana_1v8 dac_bridge(out_high=1.8 out_low=0)

.model ddflop d_dff(ic=0 rise_delay=1n fall_delay=1n)
.model dlatch d_dlatch(ic=0 rise_delay=1n fall_delay=1n)
.model dzero d_pulldown(load=1p)
.model done d_pullup(load=1p)

AA2D1 [a_VGND] [VGND] todig_1v8
AA2D2 [a_VPWR] [VPWR] todig_1v8
AA2D3 [a_force_dis_rc_osc] [force_dis_rc_osc] todig_1v8
AA2D4 [a_force_ena_rc_osc] [force_ena_rc_osc] todig_1v8
AA2D5 [a_force_pdn] [force_pdn] todig_1v8
AD2A1 [force_pdnb] [a_force_pdnb] toana_1v8
AA2D6 [a_force_short_oneshot] [force_short_oneshot] todig_1v8
AA2D7 [a_osc_ck] [osc_ck] todig_1v8
AD2A2 [osc_ena] [a_osc_ena] toana_1v8
AA2D8 [a_otrip_0_] [otrip_0_] todig_1v8
AA2D9 [a_otrip_1_] [otrip_1_] todig_1v8
AA2D10 [a_otrip_2_] [otrip_2_] todig_1v8
AD2A3 [otrip_decoded_0_] [a_otrip_decoded_0_] toana_1v8
AD2A4 [otrip_decoded_1_] [a_otrip_decoded_1_] toana_1v8
AD2A5 [otrip_decoded_2_] [a_otrip_decoded_2_] toana_1v8
AD2A6 [otrip_decoded_3_] [a_otrip_decoded_3_] toana_1v8
AD2A7 [otrip_decoded_4_] [a_otrip_decoded_4_] toana_1v8
AD2A8 [otrip_decoded_5_] [a_otrip_decoded_5_] toana_1v8
AD2A9 [otrip_decoded_6_] [a_otrip_decoded_6_] toana_1v8
AD2A10 [otrip_decoded_7_] [a_otrip_decoded_7_] toana_1v8
AD2A11 [por_timed_out] [a_por_timed_out] toana_1v8
AD2A12 [por_unbuf] [a_por_unbuf] toana_1v8
AA2D11 [a_pwup_filt] [pwup_filt] todig_1v8
AD2A13 [startup_timed_out] [a_startup_timed_out] toana_1v8

.ends


* sky130_fd_sc_hd__decap_4 (no function)
* sky130_fd_sc_hd__tapvpwrvgnd_1 (no function)
* sky130_fd_sc_hd__decap_3 (no function)
* sky130_fd_sc_hd__dfrtp_1 IQ
* sky130_fd_sc_hd__nor3b_1 (!A&!B&C_N)
.model d_lut_sky130_fd_sc_hd__nor3b_1 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "00001000")
* sky130_fd_sc_hd__buf_2 (A)
.model d_lut_sky130_fd_sc_hd__buf_2 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "01")
* sky130_fd_sc_hd__fill_1 (no function)
* sky130_fd_sc_hd__fill_2 (no function)
* sky130_fd_sc_hd__nor3_1 (!A&!B&!C)
.model d_lut_sky130_fd_sc_hd__nor3_1 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "10000000")
* sky130_ef_sc_hd__decap_12 (no function)
* sky130_fd_sc_hd__inv_2 (!A)
.model d_lut_sky130_fd_sc_hd__inv_2 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "10")
* sky130_fd_sc_hd__dlygate4sd3_1 (A)
.model d_lut_sky130_fd_sc_hd__dlygate4sd3_1 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "01")
* sky130_fd_sc_hd__xor2_1 (A&!B) | (!A&B)
.model d_lut_sky130_fd_sc_hd__xor2_1 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "0110")
* sky130_fd_sc_hd__and2b_1 (!A_N&B)
.model d_lut_sky130_fd_sc_hd__and2b_1 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "0010")
* sky130_fd_sc_hd__a41o_1 (A1&A2&A3&A4) | (B1)
.model d_lut_sky130_fd_sc_hd__a41o_1 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "00000000000000011111111111111111")
* sky130_fd_sc_hd__decap_6 (no function)
* sky130_fd_sc_hd__decap_8 (no function)
* sky130_fd_sc_hd__and2_1 (A&B)
.model d_lut_sky130_fd_sc_hd__and2_1 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "0001")
* sky130_fd_sc_hd__a21oi_1 (!A1&!B1) | (!A2&!B1)
.model d_lut_sky130_fd_sc_hd__a21oi_1 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "11100000")
* sky130_fd_sc_hd__o32a_1 (A1&B1) | (A1&B2) | (A2&B1) | (A3&B1) | (A2&B2) | (A3&B2)
.model d_lut_sky130_fd_sc_hd__o32a_1 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "00000000011111110111111101111111")
* sky130_fd_sc_hd__nand2_1 (!A) | (!B)
.model d_lut_sky130_fd_sc_hd__nand2_1 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "1110")
* sky130_fd_sc_hd__o311a_1 (A1&B1&C1) | (A2&B1&C1) | (A3&B1&C1)
.model d_lut_sky130_fd_sc_hd__o311a_1 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "00000000000000000000000001111111")
* sky130_fd_sc_hd__o21ba_1 (A1&!B1_N) | (A2&!B1_N)
.model d_lut_sky130_fd_sc_hd__o21ba_1 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "01110000")
* sky130_fd_sc_hd__o21ai_1 (!A1&!A2) | (!B1)
.model d_lut_sky130_fd_sc_hd__o21ai_1 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "11111000")
* sky130_fd_sc_hd__o211a_1 (A1&B1&C1) | (A2&B1&C1)
.model d_lut_sky130_fd_sc_hd__o211a_1 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "0000000000000111")
* sky130_fd_sc_hd__o21bai_1 (!A1&!A2) | (B1_N)
.model d_lut_sky130_fd_sc_hd__o21bai_1 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "10001111")
* sky130_fd_sc_hd__and4_1 (A&B&C&D)
.model d_lut_sky130_fd_sc_hd__and4_1 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "0000000000000001")
* sky130_fd_sc_hd__and3_1 (A&B&C)
.model d_lut_sky130_fd_sc_hd__and3_1 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "00000001")
* sky130_fd_sc_hd__clkbuf_1 (A)
.model d_lut_sky130_fd_sc_hd__clkbuf_1 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "01")
* sky130_fd_sc_hd__or4bb_1 (A) | (B) | (!C_N) | (!D_N)
.model d_lut_sky130_fd_sc_hd__or4bb_1 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "1111111111110111")
* sky130_fd_sc_hd__clkbuf_4 (A)
.model d_lut_sky130_fd_sc_hd__clkbuf_4 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "01")
* sky130_fd_sc_hd__a32o_1 (A1&A2&A3) | (B1&B2)
.model d_lut_sky130_fd_sc_hd__a32o_1 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "00000001000000010000000111111111")
* sky130_fd_sc_hd__a211oi_1 (!A1&!B1&!C1) | (!A2&!B1&!C1)
.model d_lut_sky130_fd_sc_hd__a211oi_1 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "1110000000000000")
* sky130_fd_sc_hd__buf_1 (A)
.model d_lut_sky130_fd_sc_hd__buf_1 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "01")
* sky130_fd_sc_hd__or4b_1 (A) | (B) | (C) | (!D_N)
.model d_lut_sky130_fd_sc_hd__or4b_1 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "1111111101111111")
* sky130_fd_sc_hd__conb_1 1
* sky130_fd_sc_hd__clkbuf_2 (A)
.model d_lut_sky130_fd_sc_hd__clkbuf_2 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "01")
* sky130_fd_sc_hd__dlymetal6s2s_1 (A)
.model d_lut_sky130_fd_sc_hd__dlymetal6s2s_1 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "01")
* sky130_fd_sc_hd__or3b_1 (A) | (B) | (!C_N)
.model d_lut_sky130_fd_sc_hd__or3b_1 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "11110111")
* sky130_fd_sc_hd__nand2_2 (!A) | (!B)
.model d_lut_sky130_fd_sc_hd__nand2_2 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "1110")
* sky130_fd_sc_hd__and3b_1 (!A_N&B&C)
.model d_lut_sky130_fd_sc_hd__and3b_1 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "00000010")
* sky130_fd_sc_hd__clkbuf_16 (A)
.model d_lut_sky130_fd_sc_hd__clkbuf_16 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "01")
* sky130_fd_sc_hd__and4bb_1 (!A_N&!B_N&C&D)
.model d_lut_sky130_fd_sc_hd__and4bb_1 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "0000000000001000")
* sky130_fd_sc_hd__a22o_1 (B1&B2) | (A1&A2)
.model d_lut_sky130_fd_sc_hd__a22o_1 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "0001000100011111")
* sky130_fd_sc_hd__o2bb2a_1 (!A1_N&B1) | (!A2_N&B1) | (!A1_N&B2) | (!A2_N&B2)
.model d_lut_sky130_fd_sc_hd__o2bb2a_1 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "0000111011101110")
* sky130_fd_sc_hd__or2_1 (A) | (B)
.model d_lut_sky130_fd_sc_hd__or2_1 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "0111")
* sky130_fd_sc_hd__a31o_1 (A1&A2&A3) | (B1)
.model d_lut_sky130_fd_sc_hd__a31o_1 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "0000000111111111")
* sky130_fd_sc_hd__mux2_1 (A0&!S) | (A1&S)
.model d_lut_sky130_fd_sc_hd__mux2_1 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "01010011")
* sky130_fd_sc_hd__nor2_1 (!A&!B)
.model d_lut_sky130_fd_sc_hd__nor2_1 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "1000")
.end
