magic
tech sky130A
magscale 1 2
timestamp 1712974290
<< nwell >>
rect 12433 8662 20863 9182
<< locali >>
rect 12546 8650 12610 8665
rect 12546 8616 12561 8650
rect 12595 8616 12610 8650
rect 12546 8601 12610 8616
rect 12701 8644 12765 8659
rect 12701 8546 12716 8644
rect 12750 8546 12765 8644
rect 13080 8650 13144 8665
rect 13080 8616 13095 8650
rect 13129 8616 13144 8650
rect 13080 8601 13144 8616
rect 13235 8644 13299 8659
rect 12701 8531 12765 8546
rect 13235 8546 13250 8644
rect 13284 8546 13299 8644
rect 13614 8650 13678 8665
rect 13614 8616 13629 8650
rect 13663 8616 13678 8650
rect 13614 8601 13678 8616
rect 13769 8644 13833 8659
rect 13235 8531 13299 8546
rect 13769 8546 13784 8644
rect 13818 8546 13833 8644
rect 14148 8650 14212 8665
rect 14148 8616 14163 8650
rect 14197 8616 14212 8650
rect 14148 8601 14212 8616
rect 14303 8644 14367 8659
rect 13769 8531 13833 8546
rect 14303 8546 14318 8644
rect 14352 8546 14367 8644
rect 14682 8650 14746 8665
rect 14682 8616 14697 8650
rect 14731 8616 14746 8650
rect 14682 8601 14746 8616
rect 14837 8644 14901 8659
rect 14303 8531 14367 8546
rect 14837 8546 14852 8644
rect 14886 8546 14901 8644
rect 15216 8650 15280 8665
rect 15216 8616 15231 8650
rect 15265 8616 15280 8650
rect 15216 8601 15280 8616
rect 15371 8644 15435 8659
rect 14837 8531 14901 8546
rect 15371 8546 15386 8644
rect 15420 8546 15435 8644
rect 15750 8650 15814 8665
rect 15750 8616 15765 8650
rect 15799 8616 15814 8650
rect 15750 8601 15814 8616
rect 15905 8644 15969 8659
rect 15371 8531 15435 8546
rect 15905 8546 15920 8644
rect 15954 8546 15969 8644
rect 16284 8650 16348 8665
rect 16284 8616 16299 8650
rect 16333 8616 16348 8650
rect 16284 8601 16348 8616
rect 16439 8644 16503 8659
rect 15905 8531 15969 8546
rect 16439 8546 16454 8644
rect 16488 8546 16503 8644
rect 16818 8650 16882 8665
rect 16818 8616 16833 8650
rect 16867 8616 16882 8650
rect 16818 8601 16882 8616
rect 16973 8644 17037 8659
rect 16439 8531 16503 8546
rect 16973 8546 16988 8644
rect 17022 8546 17037 8644
rect 17352 8650 17416 8665
rect 17352 8616 17367 8650
rect 17401 8616 17416 8650
rect 17352 8601 17416 8616
rect 17507 8644 17571 8659
rect 16973 8531 17037 8546
rect 17507 8546 17522 8644
rect 17556 8546 17571 8644
rect 17886 8650 17950 8665
rect 17886 8616 17901 8650
rect 17935 8616 17950 8650
rect 17886 8601 17950 8616
rect 18041 8644 18105 8659
rect 17507 8531 17571 8546
rect 18041 8546 18056 8644
rect 18090 8546 18105 8644
rect 18420 8650 18484 8665
rect 18420 8616 18435 8650
rect 18469 8616 18484 8650
rect 18420 8601 18484 8616
rect 18575 8644 18639 8659
rect 18041 8531 18105 8546
rect 18575 8546 18590 8644
rect 18624 8546 18639 8644
rect 18954 8650 19018 8665
rect 18954 8616 18969 8650
rect 19003 8616 19018 8650
rect 18954 8601 19018 8616
rect 19109 8644 19173 8659
rect 18575 8531 18639 8546
rect 19109 8546 19124 8644
rect 19158 8546 19173 8644
rect 19488 8650 19552 8665
rect 19488 8616 19503 8650
rect 19537 8616 19552 8650
rect 19488 8601 19552 8616
rect 19643 8644 19707 8659
rect 19109 8531 19173 8546
rect 19643 8546 19658 8644
rect 19692 8546 19707 8644
rect 20022 8650 20086 8665
rect 20022 8616 20037 8650
rect 20071 8616 20086 8650
rect 20022 8601 20086 8616
rect 20177 8644 20241 8659
rect 19643 8531 19707 8546
rect 20177 8546 20192 8644
rect 20226 8546 20241 8644
rect 20556 8650 20620 8665
rect 20556 8616 20571 8650
rect 20605 8616 20620 8650
rect 20556 8601 20620 8616
rect 20711 8644 20775 8659
rect 20177 8531 20241 8546
rect 20711 8546 20726 8644
rect 20760 8546 20775 8644
rect 20711 8531 20775 8546
rect 12426 8066 12490 8081
rect 21040 8066 21104 8081
rect 12426 8032 12441 8066
rect 12475 8032 12490 8066
rect 21040 8032 21055 8066
rect 21089 8032 21104 8066
rect 12426 8017 12490 8032
rect 21040 8017 21104 8032
rect 11466 7349 11530 7364
rect 11466 7251 11481 7349
rect 11515 7251 11530 7349
rect 11466 7236 11530 7251
rect 11119 7187 11183 7202
rect 11119 7089 11134 7187
rect 11168 7089 11183 7187
rect 11119 7074 11183 7089
rect 12422 6732 12486 6747
rect 21040 6732 21104 6747
rect 12422 6698 12437 6732
rect 12471 6698 12486 6732
rect 21040 6698 21055 6732
rect 21089 6698 21104 6732
rect 12422 6683 12486 6698
rect 21040 6683 21104 6698
rect 12417 6505 12475 6517
rect 15657 6505 15715 6517
rect 17446 6505 17504 6517
rect 19402 6505 19460 6517
rect 21051 6505 21109 6517
rect 12417 6471 12429 6505
rect 21051 6471 21063 6505
rect 21097 6471 21109 6505
rect 12417 6459 12475 6471
rect 15657 6459 15715 6471
rect 17446 6459 17504 6471
rect 19402 6459 19460 6471
rect 21051 6459 21109 6471
rect 8623 6383 8687 6398
rect 8623 6285 8638 6383
rect 8672 6285 8687 6383
rect 8623 6270 8687 6285
rect 11739 6383 11803 6398
rect 11739 6285 11754 6383
rect 11788 6285 11803 6383
rect 11739 6270 11803 6285
rect 12512 5179 12570 5191
rect 12512 5145 12524 5179
rect 12558 5145 12570 5179
rect 12512 5133 12570 5145
rect 14554 5179 14612 5191
rect 14554 5145 14566 5179
rect 14600 5145 14612 5179
rect 14554 5133 14612 5145
rect 16169 5188 16227 5200
rect 16169 5154 16181 5188
rect 16215 5154 16227 5188
rect 16169 5142 16227 5154
rect 18825 5185 18883 5197
rect 18825 5151 18837 5185
rect 18871 5151 18883 5185
rect 18825 5139 18883 5151
rect 20965 5183 21023 5195
rect 20965 5149 20977 5183
rect 21011 5149 21023 5183
rect 20965 5137 21023 5149
rect 500 4582 596 4616
rect 27028 4582 27124 4616
rect 500 4520 534 4582
rect 500 -3442 534 -3380
rect 27090 4520 27124 4582
rect 27090 -3442 27124 -3380
rect 500 -3476 596 -3442
rect 27028 -3476 27124 -3442
<< viali >>
rect 12561 8616 12595 8650
rect 12716 8546 12750 8644
rect 13095 8616 13129 8650
rect 13250 8546 13284 8644
rect 13629 8616 13663 8650
rect 13784 8546 13818 8644
rect 14163 8616 14197 8650
rect 14318 8546 14352 8644
rect 14697 8616 14731 8650
rect 14852 8546 14886 8644
rect 15231 8616 15265 8650
rect 15386 8546 15420 8644
rect 15765 8616 15799 8650
rect 15920 8546 15954 8644
rect 16299 8616 16333 8650
rect 16454 8546 16488 8644
rect 16833 8616 16867 8650
rect 16988 8546 17022 8644
rect 17367 8616 17401 8650
rect 17522 8546 17556 8644
rect 17901 8616 17935 8650
rect 18056 8546 18090 8644
rect 18435 8616 18469 8650
rect 18590 8546 18624 8644
rect 18969 8616 19003 8650
rect 19124 8546 19158 8644
rect 19503 8616 19537 8650
rect 19658 8546 19692 8644
rect 20037 8616 20071 8650
rect 20192 8546 20226 8644
rect 20571 8616 20605 8650
rect 20726 8546 20760 8644
rect 12441 8032 12475 8066
rect 12525 8032 21001 8066
rect 21055 8032 21089 8066
rect 11481 7251 11515 7349
rect 11134 7089 11168 7187
rect 11675 7168 11714 7204
rect 12437 6698 12471 6732
rect 12525 6698 21001 6732
rect 21055 6698 21089 6732
rect 8734 6620 11692 6654
rect 12429 6471 20905 6505
rect 21063 6471 21097 6505
rect 8638 6285 8672 6383
rect 11754 6285 11788 6383
rect 8734 5286 11692 5320
rect 12524 5145 12558 5179
rect 14566 5145 14600 5179
rect 16181 5154 16215 5188
rect 18837 5151 18871 5185
rect 20977 5149 21011 5183
rect 596 4582 27028 4616
rect 500 -3380 534 4520
rect 27090 -3380 27124 4520
rect 596 -3476 27028 -3442
<< metal1 >>
rect 11916 8974 21594 9122
rect 11916 8075 12116 8974
rect 12546 8659 12610 8665
rect 13080 8659 13144 8665
rect 13614 8659 13678 8665
rect 14148 8659 14212 8665
rect 14682 8659 14746 8665
rect 15216 8659 15280 8665
rect 15750 8659 15814 8665
rect 16284 8659 16348 8665
rect 16818 8659 16882 8665
rect 17352 8659 17416 8665
rect 17886 8659 17950 8665
rect 18420 8659 18484 8665
rect 18954 8659 19018 8665
rect 19488 8659 19552 8665
rect 20022 8659 20086 8665
rect 20556 8659 20620 8665
rect 12546 8607 12552 8659
rect 12604 8607 12610 8659
rect 12546 8601 12610 8607
rect 12701 8653 12765 8659
rect 12701 8537 12707 8653
rect 12759 8537 12765 8653
rect 13080 8607 13086 8659
rect 13138 8607 13144 8659
rect 13080 8601 13144 8607
rect 13235 8653 13299 8659
rect 12701 8531 12765 8537
rect 13235 8537 13241 8653
rect 13293 8537 13299 8653
rect 13614 8607 13620 8659
rect 13672 8607 13678 8659
rect 13614 8601 13678 8607
rect 13769 8653 13833 8659
rect 13235 8531 13299 8537
rect 13769 8537 13775 8653
rect 13827 8537 13833 8653
rect 14148 8607 14154 8659
rect 14206 8607 14212 8659
rect 14148 8601 14212 8607
rect 14303 8653 14367 8659
rect 13769 8531 13833 8537
rect 14303 8537 14309 8653
rect 14361 8537 14367 8653
rect 14682 8607 14688 8659
rect 14740 8607 14746 8659
rect 14682 8601 14746 8607
rect 14837 8653 14901 8659
rect 14303 8531 14367 8537
rect 14837 8537 14843 8653
rect 14895 8537 14901 8653
rect 15216 8607 15222 8659
rect 15274 8607 15280 8659
rect 15216 8601 15280 8607
rect 15371 8653 15435 8659
rect 14837 8531 14901 8537
rect 15371 8537 15377 8653
rect 15429 8537 15435 8653
rect 15750 8607 15756 8659
rect 15808 8607 15814 8659
rect 15750 8601 15814 8607
rect 15905 8653 15969 8659
rect 15371 8531 15435 8537
rect 15905 8537 15911 8653
rect 15963 8537 15969 8653
rect 16284 8607 16290 8659
rect 16342 8607 16348 8659
rect 16284 8601 16348 8607
rect 16439 8653 16503 8659
rect 15905 8531 15969 8537
rect 16439 8537 16445 8653
rect 16497 8537 16503 8653
rect 16818 8607 16824 8659
rect 16876 8607 16882 8659
rect 16818 8601 16882 8607
rect 16973 8653 17037 8659
rect 16439 8531 16503 8537
rect 16973 8537 16979 8653
rect 17031 8537 17037 8653
rect 17352 8607 17358 8659
rect 17410 8607 17416 8659
rect 17352 8601 17416 8607
rect 17507 8653 17571 8659
rect 16973 8531 17037 8537
rect 17507 8537 17513 8653
rect 17565 8537 17571 8653
rect 17886 8607 17892 8659
rect 17944 8607 17950 8659
rect 17886 8601 17950 8607
rect 18041 8653 18105 8659
rect 17507 8531 17571 8537
rect 18041 8537 18047 8653
rect 18099 8537 18105 8653
rect 18420 8607 18426 8659
rect 18478 8607 18484 8659
rect 18420 8601 18484 8607
rect 18575 8653 18639 8659
rect 18041 8531 18105 8537
rect 18575 8537 18581 8653
rect 18633 8537 18639 8653
rect 18954 8607 18960 8659
rect 19012 8607 19018 8659
rect 18954 8601 19018 8607
rect 19109 8653 19173 8659
rect 18575 8531 18639 8537
rect 19109 8537 19115 8653
rect 19167 8537 19173 8653
rect 19488 8607 19494 8659
rect 19546 8607 19552 8659
rect 19488 8601 19552 8607
rect 19643 8653 19707 8659
rect 19109 8531 19173 8537
rect 19643 8537 19649 8653
rect 19701 8537 19707 8653
rect 20022 8607 20028 8659
rect 20080 8607 20086 8659
rect 20022 8601 20086 8607
rect 20177 8653 20241 8659
rect 19643 8531 19707 8537
rect 20177 8537 20183 8653
rect 20235 8537 20241 8653
rect 20556 8607 20562 8659
rect 20614 8607 20620 8659
rect 20556 8601 20620 8607
rect 20711 8653 20775 8659
rect 20177 8531 20241 8537
rect 20711 8537 20717 8653
rect 20769 8537 20775 8653
rect 20711 8531 20775 8537
rect 11916 8023 11979 8075
rect 12105 8023 12116 8075
rect 11916 7675 12116 8023
rect 11462 7527 12116 7675
rect 11466 7358 11530 7364
rect 10856 7341 10984 7347
rect 10856 7289 10862 7341
rect 10978 7289 10984 7341
rect 10856 7283 10984 7289
rect 11466 7242 11472 7358
rect 11524 7242 11530 7358
rect 11466 7236 11530 7242
rect 10717 7208 10781 7214
rect 11663 7213 11727 7219
rect 10717 7092 10723 7208
rect 10775 7092 10781 7208
rect 10717 7086 10781 7092
rect 10984 7201 11058 7212
rect 10984 7075 10995 7201
rect 11047 7075 11058 7201
rect 10984 7064 11058 7075
rect 11114 7201 11188 7212
rect 11114 7075 11125 7201
rect 11177 7075 11188 7201
rect 11663 7161 11669 7213
rect 11721 7161 11727 7213
rect 11663 7155 11727 7161
rect 11114 7064 11188 7075
rect 11462 6878 11750 6963
rect 11462 6826 11613 6878
rect 11739 6826 11750 6878
rect 11462 6815 11750 6826
rect 11916 6741 12116 7527
rect 11916 6689 11979 6741
rect 12105 6689 12116 6741
rect 8626 6654 11800 6666
rect 8626 6620 8734 6654
rect 11692 6620 11800 6654
rect 8626 6608 11800 6620
rect 8626 6408 8684 6608
rect 11242 6533 11370 6539
rect 11242 6521 11248 6533
rect 8934 6481 11248 6521
rect 11364 6521 11370 6533
rect 11364 6481 11492 6521
rect 8934 6475 11492 6481
rect 11742 6408 11800 6608
rect 8618 6397 8692 6408
rect 8618 6271 8629 6397
rect 8681 6271 8692 6397
rect 8618 6260 8692 6271
rect 8752 6397 8826 6408
rect 8752 6271 8763 6397
rect 8815 6271 8826 6397
rect 8752 6260 8826 6271
rect 9108 6397 9182 6408
rect 9108 6271 9119 6397
rect 9171 6271 9182 6397
rect 9108 6260 9182 6271
rect 9464 6397 9538 6408
rect 9464 6271 9475 6397
rect 9527 6271 9538 6397
rect 9464 6260 9538 6271
rect 9820 6397 9894 6408
rect 9820 6271 9831 6397
rect 9883 6271 9894 6397
rect 9820 6260 9894 6271
rect 10176 6397 10250 6408
rect 10176 6271 10187 6397
rect 10239 6271 10250 6397
rect 10176 6260 10250 6271
rect 10532 6397 10606 6408
rect 10532 6271 10543 6397
rect 10595 6271 10606 6397
rect 10532 6260 10606 6271
rect 10888 6397 10962 6408
rect 10888 6271 10899 6397
rect 10951 6271 10962 6397
rect 10888 6260 10962 6271
rect 11244 6397 11318 6408
rect 11244 6271 11255 6397
rect 11307 6271 11318 6397
rect 11244 6260 11318 6271
rect 11600 6397 11674 6408
rect 11600 6271 11611 6397
rect 11663 6271 11674 6397
rect 11600 6260 11674 6271
rect 11734 6397 11808 6408
rect 11734 6271 11745 6397
rect 11797 6271 11808 6397
rect 11734 6260 11808 6271
rect 11916 6397 12116 6689
rect 11916 6271 11927 6397
rect 11979 6271 12116 6397
rect 8626 5332 8684 6260
rect 8930 6142 9004 6153
rect 8930 6016 8941 6142
rect 8993 6016 9004 6142
rect 8930 6005 9004 6016
rect 9286 6142 9360 6153
rect 9286 6016 9297 6142
rect 9349 6016 9360 6142
rect 9286 6005 9360 6016
rect 9642 6142 9716 6153
rect 9642 6016 9653 6142
rect 9705 6016 9716 6142
rect 9642 6005 9716 6016
rect 9998 6142 10072 6153
rect 9998 6016 10009 6142
rect 10061 6016 10072 6142
rect 9998 6005 10072 6016
rect 10354 6142 10428 6153
rect 10354 6016 10365 6142
rect 10417 6016 10428 6142
rect 10354 6005 10428 6016
rect 10710 6142 10784 6153
rect 10710 6016 10721 6142
rect 10773 6016 10784 6142
rect 10710 6005 10784 6016
rect 11066 6142 11140 6153
rect 11066 6016 11077 6142
rect 11129 6016 11140 6142
rect 11066 6005 11140 6016
rect 11422 6142 11496 6153
rect 11422 6016 11433 6142
rect 11485 6016 11496 6142
rect 11422 6005 11496 6016
rect 11742 5332 11800 6260
rect 8626 5320 11800 5332
rect 8626 5286 8734 5320
rect 11692 5286 11800 5320
rect 8626 5274 11800 5286
rect 11916 4888 12116 6271
rect 12172 8262 21338 8410
rect 12172 7133 12372 8262
rect 12421 8078 12495 8086
rect 21035 8078 21109 8086
rect 12421 8075 21109 8078
rect 12421 8023 12432 8075
rect 12484 8066 21046 8075
rect 12484 8032 12525 8066
rect 21001 8032 21046 8066
rect 12484 8023 21046 8032
rect 21098 8023 21109 8075
rect 12421 8020 21109 8023
rect 12421 8012 12495 8020
rect 12661 7945 12725 7951
rect 12661 7893 12667 7945
rect 12719 7933 12725 7945
rect 12969 7933 13017 8020
rect 13195 7945 13259 7951
rect 12719 7893 12791 7933
rect 12661 7887 12791 7893
rect 13195 7893 13201 7945
rect 13253 7933 13259 7945
rect 13503 7933 13551 8020
rect 13729 7945 13793 7951
rect 13253 7893 13325 7933
rect 13195 7887 13325 7893
rect 13729 7893 13735 7945
rect 13787 7933 13793 7945
rect 14037 7933 14085 8020
rect 14263 7945 14327 7951
rect 13787 7893 13859 7933
rect 13729 7887 13859 7893
rect 14263 7893 14269 7945
rect 14321 7933 14327 7945
rect 14571 7933 14619 8020
rect 14797 7945 14861 7951
rect 14321 7893 14393 7933
rect 14263 7887 14393 7893
rect 14797 7893 14803 7945
rect 14855 7933 14861 7945
rect 15105 7933 15153 8020
rect 15331 7945 15395 7951
rect 14855 7893 14927 7933
rect 14797 7887 14927 7893
rect 15331 7893 15337 7945
rect 15389 7933 15395 7945
rect 15639 7933 15687 8020
rect 15865 7945 15929 7951
rect 15389 7893 15461 7933
rect 15331 7887 15461 7893
rect 15865 7893 15871 7945
rect 15923 7933 15929 7945
rect 16173 7933 16221 8020
rect 16399 7945 16463 7951
rect 15923 7893 15995 7933
rect 15865 7887 15995 7893
rect 16399 7893 16405 7945
rect 16457 7933 16463 7945
rect 16707 7933 16755 8020
rect 16933 7945 16997 7951
rect 16457 7893 16529 7933
rect 16399 7887 16529 7893
rect 16933 7893 16939 7945
rect 16991 7933 16997 7945
rect 17241 7933 17289 8020
rect 17467 7945 17531 7951
rect 16991 7893 17063 7933
rect 16933 7887 17063 7893
rect 17467 7893 17473 7945
rect 17525 7933 17531 7945
rect 17775 7933 17823 8020
rect 18001 7945 18065 7951
rect 17525 7893 17597 7933
rect 17467 7887 17597 7893
rect 18001 7893 18007 7945
rect 18059 7933 18065 7945
rect 18309 7933 18357 8020
rect 18535 7945 18599 7951
rect 18059 7893 18131 7933
rect 18001 7887 18131 7893
rect 18535 7893 18541 7945
rect 18593 7933 18599 7945
rect 18843 7933 18891 8020
rect 19069 7945 19133 7951
rect 18593 7893 18665 7933
rect 18535 7887 18665 7893
rect 19069 7893 19075 7945
rect 19127 7933 19133 7945
rect 19377 7933 19425 8020
rect 19603 7945 19667 7951
rect 19127 7893 19199 7933
rect 19069 7887 19199 7893
rect 19603 7893 19609 7945
rect 19661 7933 19667 7945
rect 19911 7933 19959 8020
rect 20137 7945 20201 7951
rect 19661 7893 19733 7933
rect 19603 7887 19733 7893
rect 20137 7893 20143 7945
rect 20195 7933 20201 7945
rect 20445 7933 20493 8020
rect 21035 8012 21109 8020
rect 20671 7945 20735 7951
rect 20195 7893 20267 7933
rect 20137 7887 20267 7893
rect 20671 7893 20677 7945
rect 20729 7933 20735 7945
rect 20729 7893 20801 7933
rect 20671 7887 20801 7893
rect 12172 7007 12183 7133
rect 12235 7007 12372 7133
rect 12640 7098 12704 7102
rect 12602 7096 12704 7098
rect 12602 7044 12646 7096
rect 12698 7044 12704 7096
rect 12602 7042 12704 7044
rect 12640 7038 12704 7042
rect 12904 7096 12968 7102
rect 13174 7098 13238 7102
rect 12172 6515 12372 7007
rect 12904 6980 12910 7096
rect 12962 6980 12968 7096
rect 13136 7096 13238 7098
rect 13136 7044 13180 7096
rect 13232 7044 13238 7096
rect 13136 7042 13238 7044
rect 13174 7038 13238 7042
rect 13438 7096 13502 7102
rect 13708 7098 13772 7102
rect 12904 6974 12968 6980
rect 13438 6980 13444 7096
rect 13496 6980 13502 7096
rect 13670 7096 13772 7098
rect 13670 7044 13714 7096
rect 13766 7044 13772 7096
rect 13670 7042 13772 7044
rect 13708 7038 13772 7042
rect 13972 7096 14036 7102
rect 14242 7098 14306 7102
rect 13438 6974 13502 6980
rect 13972 6980 13978 7096
rect 14030 6980 14036 7096
rect 14204 7096 14306 7098
rect 14204 7044 14248 7096
rect 14300 7044 14306 7096
rect 14204 7042 14306 7044
rect 14242 7038 14306 7042
rect 14506 7096 14570 7102
rect 14776 7098 14840 7102
rect 13972 6974 14036 6980
rect 14506 6980 14512 7096
rect 14564 6980 14570 7096
rect 14738 7096 14840 7098
rect 14738 7044 14782 7096
rect 14834 7044 14840 7096
rect 14738 7042 14840 7044
rect 14776 7038 14840 7042
rect 15040 7096 15104 7102
rect 15310 7098 15374 7102
rect 14506 6974 14570 6980
rect 15040 6980 15046 7096
rect 15098 6980 15104 7096
rect 15272 7096 15374 7098
rect 15272 7044 15316 7096
rect 15368 7044 15374 7096
rect 15272 7042 15374 7044
rect 15310 7038 15374 7042
rect 15574 7096 15638 7102
rect 15844 7098 15908 7102
rect 15040 6974 15104 6980
rect 15574 6980 15580 7096
rect 15632 6980 15638 7096
rect 15806 7096 15908 7098
rect 15806 7044 15850 7096
rect 15902 7044 15908 7096
rect 15806 7042 15908 7044
rect 15844 7038 15908 7042
rect 16108 7096 16172 7102
rect 16378 7098 16442 7102
rect 15574 6974 15638 6980
rect 16108 6980 16114 7096
rect 16166 6980 16172 7096
rect 16340 7096 16442 7098
rect 16340 7044 16384 7096
rect 16436 7044 16442 7096
rect 16340 7042 16442 7044
rect 16378 7038 16442 7042
rect 16642 7096 16706 7102
rect 16912 7098 16976 7102
rect 16108 6974 16172 6980
rect 16642 6980 16648 7096
rect 16700 6980 16706 7096
rect 16874 7096 16976 7098
rect 16874 7044 16918 7096
rect 16970 7044 16976 7096
rect 16874 7042 16976 7044
rect 16912 7038 16976 7042
rect 17176 7096 17240 7102
rect 17446 7098 17510 7102
rect 16642 6974 16706 6980
rect 17176 6980 17182 7096
rect 17234 6980 17240 7096
rect 17408 7096 17510 7098
rect 17408 7044 17452 7096
rect 17504 7044 17510 7096
rect 17408 7042 17510 7044
rect 17446 7038 17510 7042
rect 17710 7096 17774 7102
rect 17980 7098 18044 7102
rect 17176 6974 17240 6980
rect 17710 6980 17716 7096
rect 17768 6980 17774 7096
rect 17942 7096 18044 7098
rect 17942 7044 17986 7096
rect 18038 7044 18044 7096
rect 17942 7042 18044 7044
rect 17980 7038 18044 7042
rect 18244 7096 18308 7102
rect 18514 7098 18578 7102
rect 17710 6974 17774 6980
rect 18244 6980 18250 7096
rect 18302 6980 18308 7096
rect 18476 7096 18578 7098
rect 18476 7044 18520 7096
rect 18572 7044 18578 7096
rect 18476 7042 18578 7044
rect 18514 7038 18578 7042
rect 18778 7096 18842 7102
rect 19048 7098 19112 7102
rect 18244 6974 18308 6980
rect 18778 6980 18784 7096
rect 18836 6980 18842 7096
rect 19010 7096 19112 7098
rect 19010 7044 19054 7096
rect 19106 7044 19112 7096
rect 19010 7042 19112 7044
rect 19048 7038 19112 7042
rect 19312 7096 19376 7102
rect 19582 7098 19646 7102
rect 18778 6974 18842 6980
rect 19312 6980 19318 7096
rect 19370 6980 19376 7096
rect 19544 7096 19646 7098
rect 19544 7044 19588 7096
rect 19640 7044 19646 7096
rect 19544 7042 19646 7044
rect 19582 7038 19646 7042
rect 19846 7096 19910 7102
rect 20116 7098 20180 7102
rect 19312 6974 19376 6980
rect 19846 6980 19852 7096
rect 19904 6980 19910 7096
rect 20078 7096 20180 7098
rect 20078 7044 20122 7096
rect 20174 7044 20180 7096
rect 20078 7042 20180 7044
rect 20116 7038 20180 7042
rect 20380 7096 20444 7102
rect 20650 7098 20714 7102
rect 19846 6974 19910 6980
rect 20380 6980 20386 7096
rect 20438 6980 20444 7096
rect 20612 7096 20714 7098
rect 20612 7044 20656 7096
rect 20708 7044 20714 7096
rect 20612 7042 20714 7044
rect 20650 7038 20714 7042
rect 20914 7096 20978 7102
rect 20380 6974 20444 6980
rect 20914 6980 20920 7096
rect 20972 6980 20978 7096
rect 20914 6974 20978 6980
rect 12726 6965 12790 6971
rect 12726 6849 12732 6965
rect 12784 6849 12790 6965
rect 12726 6843 12790 6849
rect 13260 6968 13324 6974
rect 13260 6852 13266 6968
rect 13318 6852 13324 6968
rect 13260 6846 13324 6852
rect 13794 6968 13858 6974
rect 13794 6852 13800 6968
rect 13852 6852 13858 6968
rect 13794 6846 13858 6852
rect 14328 6968 14392 6974
rect 14328 6852 14334 6968
rect 14386 6852 14392 6968
rect 14328 6846 14392 6852
rect 14862 6968 14926 6974
rect 14862 6852 14868 6968
rect 14920 6852 14926 6968
rect 14862 6846 14926 6852
rect 15396 6968 15460 6974
rect 15396 6852 15402 6968
rect 15454 6852 15460 6968
rect 15396 6846 15460 6852
rect 15930 6968 15994 6974
rect 15930 6852 15936 6968
rect 15988 6852 15994 6968
rect 15930 6846 15994 6852
rect 16464 6968 16528 6974
rect 16464 6852 16470 6968
rect 16522 6852 16528 6968
rect 16464 6846 16528 6852
rect 16998 6968 17062 6974
rect 16998 6852 17004 6968
rect 17056 6852 17062 6968
rect 16998 6846 17062 6852
rect 17532 6968 17596 6974
rect 17532 6852 17538 6968
rect 17590 6852 17596 6968
rect 17532 6846 17596 6852
rect 18066 6968 18130 6974
rect 18066 6852 18072 6968
rect 18124 6852 18130 6968
rect 18066 6846 18130 6852
rect 18600 6968 18664 6974
rect 18600 6852 18606 6968
rect 18658 6852 18664 6968
rect 18600 6846 18664 6852
rect 19134 6968 19198 6974
rect 19134 6852 19140 6968
rect 19192 6852 19198 6968
rect 19134 6846 19198 6852
rect 19668 6968 19732 6974
rect 19668 6852 19674 6968
rect 19726 6852 19732 6968
rect 19668 6846 19732 6852
rect 20202 6968 20266 6974
rect 20202 6852 20208 6968
rect 20260 6852 20266 6968
rect 20202 6846 20266 6852
rect 20736 6968 20800 6974
rect 20736 6852 20742 6968
rect 20794 6852 20800 6968
rect 20736 6846 20800 6852
rect 12417 6744 12491 6752
rect 21035 6744 21109 6752
rect 12417 6741 21109 6744
rect 12417 6689 12428 6741
rect 12480 6732 21046 6741
rect 12480 6698 12525 6732
rect 21001 6698 21046 6732
rect 12480 6689 21046 6698
rect 21098 6689 21109 6741
rect 12417 6686 21109 6689
rect 12417 6678 12491 6686
rect 21035 6678 21109 6686
rect 12417 6515 12475 6517
rect 15657 6515 15715 6517
rect 17446 6515 17504 6517
rect 19402 6515 19460 6517
rect 21051 6515 21109 6517
rect 21138 6515 21338 8262
rect 12172 6505 21338 6515
rect 12172 6471 12429 6505
rect 20905 6471 21063 6505
rect 21097 6471 21338 6505
rect 12172 6460 21338 6471
rect 12172 5144 12372 6460
rect 12417 6459 12475 6460
rect 12613 6385 12677 6391
rect 12613 6333 12619 6385
rect 12671 6333 12677 6385
rect 12613 6327 12677 6333
rect 12725 6327 12791 6373
rect 12965 6367 13021 6460
rect 13147 6385 13211 6391
rect 13147 6333 13153 6385
rect 13205 6333 13211 6385
rect 13147 6327 13211 6333
rect 13259 6327 13325 6373
rect 13499 6367 13555 6460
rect 13681 6385 13745 6391
rect 13681 6333 13687 6385
rect 13739 6333 13745 6385
rect 13681 6327 13745 6333
rect 13793 6327 13859 6373
rect 14033 6367 14089 6460
rect 14215 6385 14279 6391
rect 14215 6333 14221 6385
rect 14273 6333 14279 6385
rect 14215 6327 14279 6333
rect 14327 6327 14393 6373
rect 14567 6367 14623 6460
rect 14749 6385 14813 6391
rect 14749 6333 14755 6385
rect 14807 6333 14813 6385
rect 14749 6327 14813 6333
rect 14861 6327 14927 6373
rect 15101 6367 15157 6460
rect 15635 6459 15715 6460
rect 15283 6385 15347 6391
rect 15283 6333 15289 6385
rect 15341 6333 15347 6385
rect 15283 6327 15347 6333
rect 15395 6327 15461 6373
rect 15635 6367 15691 6459
rect 15817 6385 15881 6391
rect 15817 6333 15823 6385
rect 15875 6333 15881 6385
rect 15817 6327 15881 6333
rect 15929 6327 15995 6373
rect 16169 6367 16225 6460
rect 16351 6385 16415 6391
rect 16351 6333 16357 6385
rect 16409 6333 16415 6385
rect 16351 6327 16415 6333
rect 16463 6327 16529 6373
rect 16703 6367 16759 6460
rect 16885 6385 16949 6391
rect 16885 6333 16891 6385
rect 16943 6333 16949 6385
rect 16885 6327 16949 6333
rect 16997 6327 17063 6373
rect 17237 6367 17293 6460
rect 17446 6459 17504 6460
rect 17419 6385 17483 6391
rect 17419 6333 17425 6385
rect 17477 6333 17483 6385
rect 17419 6327 17483 6333
rect 17531 6327 17597 6373
rect 17771 6367 17827 6460
rect 17953 6385 18017 6391
rect 17953 6333 17959 6385
rect 18011 6333 18017 6385
rect 17953 6327 18017 6333
rect 18065 6327 18131 6373
rect 18305 6367 18361 6460
rect 18487 6385 18551 6391
rect 18487 6333 18493 6385
rect 18545 6333 18551 6385
rect 18487 6327 18551 6333
rect 18599 6327 18665 6373
rect 18839 6367 18895 6460
rect 19373 6459 19460 6460
rect 19021 6385 19085 6391
rect 19021 6333 19027 6385
rect 19079 6333 19085 6385
rect 19021 6327 19085 6333
rect 19133 6327 19199 6373
rect 19373 6367 19429 6459
rect 19555 6385 19619 6391
rect 19555 6333 19561 6385
rect 19613 6333 19619 6385
rect 19555 6327 19619 6333
rect 19667 6327 19733 6373
rect 19907 6367 19963 6460
rect 20089 6385 20153 6391
rect 20089 6333 20095 6385
rect 20147 6333 20153 6385
rect 20089 6327 20153 6333
rect 20201 6327 20267 6373
rect 20441 6367 20497 6460
rect 21051 6459 21109 6460
rect 20623 6385 20687 6391
rect 20623 6333 20629 6385
rect 20681 6333 20687 6385
rect 20623 6327 20687 6333
rect 20735 6327 20801 6373
rect 12726 6286 12790 6292
rect 12548 6182 12612 6188
rect 12548 6066 12554 6182
rect 12606 6066 12612 6182
rect 12726 6170 12732 6286
rect 12784 6170 12790 6286
rect 13260 6289 13324 6295
rect 12726 6164 12790 6170
rect 12904 6182 12968 6188
rect 12548 6060 12612 6066
rect 12904 6066 12910 6182
rect 12962 6066 12968 6182
rect 12904 6060 12968 6066
rect 13082 6182 13146 6188
rect 13082 6066 13088 6182
rect 13140 6066 13146 6182
rect 13260 6173 13266 6289
rect 13318 6173 13324 6289
rect 13794 6289 13858 6295
rect 13260 6167 13324 6173
rect 13438 6182 13502 6188
rect 13082 6060 13146 6066
rect 13438 6066 13444 6182
rect 13496 6066 13502 6182
rect 13438 6060 13502 6066
rect 13616 6182 13680 6188
rect 13616 6066 13622 6182
rect 13674 6066 13680 6182
rect 13794 6173 13800 6289
rect 13852 6173 13858 6289
rect 14328 6289 14392 6295
rect 13794 6167 13858 6173
rect 13972 6182 14036 6188
rect 13616 6060 13680 6066
rect 13972 6066 13978 6182
rect 14030 6066 14036 6182
rect 13972 6060 14036 6066
rect 14150 6182 14214 6188
rect 14150 6066 14156 6182
rect 14208 6066 14214 6182
rect 14328 6173 14334 6289
rect 14386 6173 14392 6289
rect 14862 6289 14926 6295
rect 14328 6167 14392 6173
rect 14506 6182 14570 6188
rect 14150 6060 14214 6066
rect 14506 6066 14512 6182
rect 14564 6066 14570 6182
rect 14506 6060 14570 6066
rect 14684 6182 14748 6188
rect 14684 6066 14690 6182
rect 14742 6066 14748 6182
rect 14862 6173 14868 6289
rect 14920 6173 14926 6289
rect 15396 6289 15460 6295
rect 14862 6167 14926 6173
rect 15040 6182 15104 6188
rect 14684 6060 14748 6066
rect 15040 6066 15046 6182
rect 15098 6066 15104 6182
rect 15040 6060 15104 6066
rect 15218 6182 15282 6188
rect 15218 6066 15224 6182
rect 15276 6066 15282 6182
rect 15396 6173 15402 6289
rect 15454 6173 15460 6289
rect 15930 6289 15994 6295
rect 15396 6167 15460 6173
rect 15574 6182 15638 6188
rect 15218 6060 15282 6066
rect 15574 6066 15580 6182
rect 15632 6066 15638 6182
rect 15574 6060 15638 6066
rect 15752 6182 15816 6188
rect 15752 6066 15758 6182
rect 15810 6066 15816 6182
rect 15930 6173 15936 6289
rect 15988 6173 15994 6289
rect 16464 6289 16528 6295
rect 15930 6167 15994 6173
rect 16108 6182 16172 6188
rect 15752 6060 15816 6066
rect 16108 6066 16114 6182
rect 16166 6066 16172 6182
rect 16108 6060 16172 6066
rect 16286 6182 16350 6188
rect 16286 6066 16292 6182
rect 16344 6066 16350 6182
rect 16464 6173 16470 6289
rect 16522 6173 16528 6289
rect 16998 6289 17062 6295
rect 16464 6167 16528 6173
rect 16642 6182 16706 6188
rect 16286 6060 16350 6066
rect 16642 6066 16648 6182
rect 16700 6066 16706 6182
rect 16642 6060 16706 6066
rect 16820 6182 16884 6188
rect 16820 6066 16826 6182
rect 16878 6066 16884 6182
rect 16998 6173 17004 6289
rect 17056 6173 17062 6289
rect 17532 6289 17596 6295
rect 16998 6167 17062 6173
rect 17176 6182 17240 6188
rect 16820 6060 16884 6066
rect 17176 6066 17182 6182
rect 17234 6066 17240 6182
rect 17176 6060 17240 6066
rect 17354 6182 17418 6188
rect 17354 6066 17360 6182
rect 17412 6066 17418 6182
rect 17532 6173 17538 6289
rect 17590 6173 17596 6289
rect 18066 6289 18130 6295
rect 17532 6167 17596 6173
rect 17710 6182 17774 6188
rect 17354 6060 17418 6066
rect 17710 6066 17716 6182
rect 17768 6066 17774 6182
rect 17710 6060 17774 6066
rect 17888 6182 17952 6188
rect 17888 6066 17894 6182
rect 17946 6066 17952 6182
rect 18066 6173 18072 6289
rect 18124 6173 18130 6289
rect 18600 6289 18664 6295
rect 18066 6167 18130 6173
rect 18244 6182 18308 6188
rect 17888 6060 17952 6066
rect 18244 6066 18250 6182
rect 18302 6066 18308 6182
rect 18244 6060 18308 6066
rect 18422 6182 18486 6188
rect 18422 6066 18428 6182
rect 18480 6066 18486 6182
rect 18600 6173 18606 6289
rect 18658 6173 18664 6289
rect 19134 6289 19198 6295
rect 18600 6167 18664 6173
rect 18778 6182 18842 6188
rect 18422 6060 18486 6066
rect 18778 6066 18784 6182
rect 18836 6066 18842 6182
rect 18778 6060 18842 6066
rect 18956 6182 19020 6188
rect 18956 6066 18962 6182
rect 19014 6066 19020 6182
rect 19134 6173 19140 6289
rect 19192 6173 19198 6289
rect 19668 6289 19732 6295
rect 19134 6167 19198 6173
rect 19312 6182 19376 6188
rect 18956 6060 19020 6066
rect 19312 6066 19318 6182
rect 19370 6066 19376 6182
rect 19312 6060 19376 6066
rect 19490 6182 19554 6188
rect 19490 6066 19496 6182
rect 19548 6066 19554 6182
rect 19668 6173 19674 6289
rect 19726 6173 19732 6289
rect 20202 6289 20266 6295
rect 19668 6167 19732 6173
rect 19846 6182 19910 6188
rect 19490 6060 19554 6066
rect 19846 6066 19852 6182
rect 19904 6066 19910 6182
rect 19846 6060 19910 6066
rect 20024 6182 20088 6188
rect 20024 6066 20030 6182
rect 20082 6066 20088 6182
rect 20202 6173 20208 6289
rect 20260 6173 20266 6289
rect 20736 6289 20800 6295
rect 20202 6167 20266 6173
rect 20380 6182 20444 6188
rect 20024 6060 20088 6066
rect 20380 6066 20386 6182
rect 20438 6066 20444 6182
rect 20380 6060 20444 6066
rect 20558 6182 20622 6188
rect 20558 6066 20564 6182
rect 20616 6066 20622 6182
rect 20736 6173 20742 6289
rect 20794 6173 20800 6289
rect 20736 6167 20800 6173
rect 20914 6182 20978 6188
rect 20558 6060 20622 6066
rect 20914 6066 20920 6182
rect 20972 6066 20978 6182
rect 20914 6060 20978 6066
rect 12726 5432 12790 5438
rect 12726 5316 12732 5432
rect 12784 5316 12790 5432
rect 12726 5310 12790 5316
rect 13260 5435 13324 5441
rect 13260 5319 13266 5435
rect 13318 5319 13324 5435
rect 13260 5313 13324 5319
rect 13794 5435 13858 5441
rect 13794 5319 13800 5435
rect 13852 5319 13858 5435
rect 13794 5313 13858 5319
rect 14328 5435 14392 5441
rect 14328 5319 14334 5435
rect 14386 5319 14392 5435
rect 14328 5313 14392 5319
rect 14862 5435 14926 5441
rect 14862 5319 14868 5435
rect 14920 5319 14926 5435
rect 14862 5313 14926 5319
rect 15396 5435 15460 5441
rect 15396 5319 15402 5435
rect 15454 5319 15460 5435
rect 15396 5313 15460 5319
rect 15930 5435 15994 5441
rect 15930 5319 15936 5435
rect 15988 5319 15994 5435
rect 15930 5313 15994 5319
rect 16464 5435 16528 5441
rect 16464 5319 16470 5435
rect 16522 5319 16528 5435
rect 16464 5313 16528 5319
rect 16998 5435 17062 5441
rect 16998 5319 17004 5435
rect 17056 5319 17062 5435
rect 16998 5313 17062 5319
rect 17532 5435 17596 5441
rect 17532 5319 17538 5435
rect 17590 5319 17596 5435
rect 17532 5313 17596 5319
rect 18066 5435 18130 5441
rect 18066 5319 18072 5435
rect 18124 5319 18130 5435
rect 18066 5313 18130 5319
rect 18600 5435 18664 5441
rect 18600 5319 18606 5435
rect 18658 5319 18664 5435
rect 18600 5313 18664 5319
rect 19134 5435 19198 5441
rect 19134 5319 19140 5435
rect 19192 5319 19198 5435
rect 19134 5313 19198 5319
rect 19668 5435 19732 5441
rect 19668 5319 19674 5435
rect 19726 5319 19732 5435
rect 19668 5313 19732 5319
rect 20202 5435 20266 5441
rect 20202 5319 20208 5435
rect 20260 5319 20266 5435
rect 20202 5313 20266 5319
rect 20736 5435 20800 5441
rect 20736 5319 20742 5435
rect 20794 5319 20800 5435
rect 20736 5313 20800 5319
rect 12512 5179 12570 5191
rect 12512 5145 12524 5179
rect 12558 5145 12570 5179
rect 12512 5144 12570 5145
rect 14554 5179 14612 5191
rect 14554 5145 14566 5179
rect 14600 5145 14612 5179
rect 14554 5144 14612 5145
rect 16169 5188 16227 5200
rect 16169 5154 16181 5188
rect 16215 5154 16227 5188
rect 16169 5144 16227 5154
rect 18825 5185 18883 5197
rect 18825 5151 18837 5185
rect 18871 5151 18883 5185
rect 18825 5144 18883 5151
rect 20965 5183 21023 5195
rect 20965 5149 20977 5183
rect 21011 5149 21023 5183
rect 20965 5144 21023 5149
rect 21138 5144 21338 6460
rect 12172 5084 21338 5144
rect 12172 5002 21198 5084
rect 12172 4950 12476 5002
rect 12592 4952 21198 5002
rect 21330 4952 21338 5084
rect 12592 4950 21338 4952
rect 12172 4944 21338 4950
rect 21394 8075 21594 8974
rect 21394 8023 21405 8075
rect 21531 8023 21594 8075
rect 21394 6741 21594 8023
rect 21394 6689 21405 6741
rect 21531 6689 21594 6741
rect 21394 4888 21594 6689
rect 11916 4688 21594 4888
rect 12470 4628 12598 4632
rect 489 4626 27136 4628
rect 489 4616 12476 4626
rect 12592 4616 27136 4626
rect 489 4582 596 4616
rect 27028 4582 27136 4616
rect 489 4574 12476 4582
rect 12592 4574 27136 4582
rect 489 4572 27136 4574
rect 489 4520 545 4572
rect 12470 4568 12598 4572
rect 489 -3380 500 4520
rect 534 -3380 545 4520
rect 27080 4520 27136 4572
rect 27080 4480 27090 4520
rect 691 4312 697 4460
rect 845 4312 851 4460
rect 1280 4059 1396 4480
rect 2036 4059 2152 4480
rect 2792 4059 2908 4480
rect 3548 4059 3664 4480
rect 4304 4059 4420 4480
rect 5060 4059 5176 4480
rect 5816 4059 5932 4480
rect 6572 4059 6688 4480
rect 7328 4059 7444 4480
rect 8084 4059 8200 4480
rect 8840 4059 8956 4480
rect 9596 4059 9712 4480
rect 10352 4059 10468 4480
rect 11108 4059 11224 4480
rect 11864 4059 11980 4480
rect 12620 4059 12736 4480
rect 13376 4059 13492 4480
rect 14132 4474 14248 4480
rect 14132 4358 14164 4474
rect 14216 4358 14248 4474
rect 14132 4059 14248 4358
rect 14888 4474 15004 4480
rect 14888 4358 14920 4474
rect 14972 4358 15004 4474
rect 14888 4059 15004 4358
rect 15644 4474 15760 4480
rect 15644 4358 15676 4474
rect 15728 4358 15760 4474
rect 15644 4059 15760 4358
rect 16400 4474 16516 4480
rect 16400 4358 16432 4474
rect 16484 4358 16516 4474
rect 16400 4059 16516 4358
rect 17156 4059 17272 4480
rect 17912 4059 18028 4480
rect 18668 4059 18784 4480
rect 19424 4059 19540 4480
rect 20180 4059 20296 4480
rect 20936 4059 21052 4480
rect 21692 4059 21808 4480
rect 22448 4059 22564 4480
rect 23204 4059 23320 4480
rect 23960 4059 24076 4480
rect 24716 4059 24832 4480
rect 25472 4059 25588 4480
rect 26228 4059 26344 4480
rect 26773 4313 26779 4461
rect 26927 4313 26933 4461
rect 27079 4059 27090 4480
rect 902 -3340 1018 -2919
rect 1658 -3340 1774 -2919
rect 2414 -3340 2530 -2919
rect 3170 -3340 3286 -2919
rect 3926 -3340 4042 -2919
rect 4682 -3340 4798 -2919
rect 5438 -3340 5554 -2919
rect 6194 -3340 6310 -2919
rect 6950 -3340 7066 -2919
rect 7706 -3340 7822 -2919
rect 8462 -3340 8578 -2919
rect 9218 -3340 9334 -2919
rect 9974 -3340 10090 -2919
rect 10730 -3340 10846 -2919
rect 11486 -3340 11602 -2919
rect 12242 -3340 12358 -2919
rect 12998 -3340 13114 -2919
rect 13754 -2990 13870 -2919
rect 13754 -3046 13785 -2990
rect 13841 -3046 13870 -2990
rect 13754 -3340 13870 -3046
rect 14510 -2976 14626 -2919
rect 14510 -3032 14541 -2976
rect 14597 -3032 14626 -2976
rect 14510 -3340 14626 -3032
rect 15266 -2990 15382 -2919
rect 15266 -3046 15297 -2990
rect 15353 -3046 15382 -2990
rect 15266 -3340 15382 -3046
rect 16022 -2990 16138 -2919
rect 16022 -3046 16053 -2990
rect 16109 -3046 16138 -2990
rect 16022 -3340 16138 -3046
rect 16778 -3340 16894 -2919
rect 17534 -3340 17650 -2919
rect 18290 -3340 18406 -2919
rect 19046 -3340 19162 -2919
rect 19802 -3340 19918 -2919
rect 20558 -3340 20674 -2919
rect 21314 -3340 21430 -2919
rect 22070 -3340 22186 -2919
rect 22826 -3340 22942 -2919
rect 23582 -3340 23698 -2919
rect 24338 -3340 24454 -2919
rect 25094 -3340 25210 -2919
rect 25850 -3340 25966 -2919
rect 26606 -3340 26722 -2919
rect 489 -3431 545 -3380
rect 27080 -3380 27090 4059
rect 27124 -3380 27136 4520
rect 27080 -3431 27136 -3380
rect 489 -3442 27136 -3431
rect 489 -3476 596 -3442
rect 27028 -3476 27136 -3442
rect 489 -3487 27136 -3476
<< via1 >>
rect 12552 8650 12604 8659
rect 12552 8616 12561 8650
rect 12561 8616 12595 8650
rect 12595 8616 12604 8650
rect 12552 8607 12604 8616
rect 12707 8644 12759 8653
rect 12707 8546 12716 8644
rect 12716 8546 12750 8644
rect 12750 8546 12759 8644
rect 12707 8537 12759 8546
rect 13086 8650 13138 8659
rect 13086 8616 13095 8650
rect 13095 8616 13129 8650
rect 13129 8616 13138 8650
rect 13086 8607 13138 8616
rect 13241 8644 13293 8653
rect 13241 8546 13250 8644
rect 13250 8546 13284 8644
rect 13284 8546 13293 8644
rect 13241 8537 13293 8546
rect 13620 8650 13672 8659
rect 13620 8616 13629 8650
rect 13629 8616 13663 8650
rect 13663 8616 13672 8650
rect 13620 8607 13672 8616
rect 13775 8644 13827 8653
rect 13775 8546 13784 8644
rect 13784 8546 13818 8644
rect 13818 8546 13827 8644
rect 13775 8537 13827 8546
rect 14154 8650 14206 8659
rect 14154 8616 14163 8650
rect 14163 8616 14197 8650
rect 14197 8616 14206 8650
rect 14154 8607 14206 8616
rect 14309 8644 14361 8653
rect 14309 8546 14318 8644
rect 14318 8546 14352 8644
rect 14352 8546 14361 8644
rect 14309 8537 14361 8546
rect 14688 8650 14740 8659
rect 14688 8616 14697 8650
rect 14697 8616 14731 8650
rect 14731 8616 14740 8650
rect 14688 8607 14740 8616
rect 14843 8644 14895 8653
rect 14843 8546 14852 8644
rect 14852 8546 14886 8644
rect 14886 8546 14895 8644
rect 14843 8537 14895 8546
rect 15222 8650 15274 8659
rect 15222 8616 15231 8650
rect 15231 8616 15265 8650
rect 15265 8616 15274 8650
rect 15222 8607 15274 8616
rect 15377 8644 15429 8653
rect 15377 8546 15386 8644
rect 15386 8546 15420 8644
rect 15420 8546 15429 8644
rect 15377 8537 15429 8546
rect 15756 8650 15808 8659
rect 15756 8616 15765 8650
rect 15765 8616 15799 8650
rect 15799 8616 15808 8650
rect 15756 8607 15808 8616
rect 15911 8644 15963 8653
rect 15911 8546 15920 8644
rect 15920 8546 15954 8644
rect 15954 8546 15963 8644
rect 15911 8537 15963 8546
rect 16290 8650 16342 8659
rect 16290 8616 16299 8650
rect 16299 8616 16333 8650
rect 16333 8616 16342 8650
rect 16290 8607 16342 8616
rect 16445 8644 16497 8653
rect 16445 8546 16454 8644
rect 16454 8546 16488 8644
rect 16488 8546 16497 8644
rect 16445 8537 16497 8546
rect 16824 8650 16876 8659
rect 16824 8616 16833 8650
rect 16833 8616 16867 8650
rect 16867 8616 16876 8650
rect 16824 8607 16876 8616
rect 16979 8644 17031 8653
rect 16979 8546 16988 8644
rect 16988 8546 17022 8644
rect 17022 8546 17031 8644
rect 16979 8537 17031 8546
rect 17358 8650 17410 8659
rect 17358 8616 17367 8650
rect 17367 8616 17401 8650
rect 17401 8616 17410 8650
rect 17358 8607 17410 8616
rect 17513 8644 17565 8653
rect 17513 8546 17522 8644
rect 17522 8546 17556 8644
rect 17556 8546 17565 8644
rect 17513 8537 17565 8546
rect 17892 8650 17944 8659
rect 17892 8616 17901 8650
rect 17901 8616 17935 8650
rect 17935 8616 17944 8650
rect 17892 8607 17944 8616
rect 18047 8644 18099 8653
rect 18047 8546 18056 8644
rect 18056 8546 18090 8644
rect 18090 8546 18099 8644
rect 18047 8537 18099 8546
rect 18426 8650 18478 8659
rect 18426 8616 18435 8650
rect 18435 8616 18469 8650
rect 18469 8616 18478 8650
rect 18426 8607 18478 8616
rect 18581 8644 18633 8653
rect 18581 8546 18590 8644
rect 18590 8546 18624 8644
rect 18624 8546 18633 8644
rect 18581 8537 18633 8546
rect 18960 8650 19012 8659
rect 18960 8616 18969 8650
rect 18969 8616 19003 8650
rect 19003 8616 19012 8650
rect 18960 8607 19012 8616
rect 19115 8644 19167 8653
rect 19115 8546 19124 8644
rect 19124 8546 19158 8644
rect 19158 8546 19167 8644
rect 19115 8537 19167 8546
rect 19494 8650 19546 8659
rect 19494 8616 19503 8650
rect 19503 8616 19537 8650
rect 19537 8616 19546 8650
rect 19494 8607 19546 8616
rect 19649 8644 19701 8653
rect 19649 8546 19658 8644
rect 19658 8546 19692 8644
rect 19692 8546 19701 8644
rect 19649 8537 19701 8546
rect 20028 8650 20080 8659
rect 20028 8616 20037 8650
rect 20037 8616 20071 8650
rect 20071 8616 20080 8650
rect 20028 8607 20080 8616
rect 20183 8644 20235 8653
rect 20183 8546 20192 8644
rect 20192 8546 20226 8644
rect 20226 8546 20235 8644
rect 20183 8537 20235 8546
rect 20562 8650 20614 8659
rect 20562 8616 20571 8650
rect 20571 8616 20605 8650
rect 20605 8616 20614 8650
rect 20562 8607 20614 8616
rect 20717 8644 20769 8653
rect 20717 8546 20726 8644
rect 20726 8546 20760 8644
rect 20760 8546 20769 8644
rect 20717 8537 20769 8546
rect 11979 8023 12105 8075
rect 10862 7289 10978 7341
rect 11472 7349 11524 7358
rect 11472 7251 11481 7349
rect 11481 7251 11515 7349
rect 11515 7251 11524 7349
rect 11472 7242 11524 7251
rect 10723 7092 10775 7208
rect 10995 7075 11047 7201
rect 11125 7187 11177 7201
rect 11125 7089 11134 7187
rect 11134 7089 11168 7187
rect 11168 7089 11177 7187
rect 11125 7075 11177 7089
rect 11669 7204 11721 7213
rect 11669 7168 11675 7204
rect 11675 7168 11714 7204
rect 11714 7168 11721 7204
rect 11669 7161 11721 7168
rect 11613 6826 11739 6878
rect 11979 6689 12105 6741
rect 11248 6481 11364 6533
rect 8629 6383 8681 6397
rect 8629 6285 8638 6383
rect 8638 6285 8672 6383
rect 8672 6285 8681 6383
rect 8629 6271 8681 6285
rect 8763 6271 8815 6397
rect 9119 6271 9171 6397
rect 9475 6271 9527 6397
rect 9831 6271 9883 6397
rect 10187 6271 10239 6397
rect 10543 6271 10595 6397
rect 10899 6271 10951 6397
rect 11255 6271 11307 6397
rect 11611 6271 11663 6397
rect 11745 6383 11797 6397
rect 11745 6285 11754 6383
rect 11754 6285 11788 6383
rect 11788 6285 11797 6383
rect 11745 6271 11797 6285
rect 11927 6271 11979 6397
rect 8941 6016 8993 6142
rect 9297 6016 9349 6142
rect 9653 6016 9705 6142
rect 10009 6016 10061 6142
rect 10365 6016 10417 6142
rect 10721 6016 10773 6142
rect 11077 6016 11129 6142
rect 11433 6016 11485 6142
rect 12432 8066 12484 8075
rect 21046 8066 21098 8075
rect 12432 8032 12441 8066
rect 12441 8032 12475 8066
rect 12475 8032 12484 8066
rect 21046 8032 21055 8066
rect 21055 8032 21089 8066
rect 21089 8032 21098 8066
rect 12432 8023 12484 8032
rect 21046 8023 21098 8032
rect 12667 7893 12719 7945
rect 13201 7893 13253 7945
rect 13735 7893 13787 7945
rect 14269 7893 14321 7945
rect 14803 7893 14855 7945
rect 15337 7893 15389 7945
rect 15871 7893 15923 7945
rect 16405 7893 16457 7945
rect 16939 7893 16991 7945
rect 17473 7893 17525 7945
rect 18007 7893 18059 7945
rect 18541 7893 18593 7945
rect 19075 7893 19127 7945
rect 19609 7893 19661 7945
rect 20143 7893 20195 7945
rect 20677 7893 20729 7945
rect 12183 7007 12235 7133
rect 12646 7044 12698 7096
rect 12910 6980 12962 7096
rect 13180 7044 13232 7096
rect 13444 6980 13496 7096
rect 13714 7044 13766 7096
rect 13978 6980 14030 7096
rect 14248 7044 14300 7096
rect 14512 6980 14564 7096
rect 14782 7044 14834 7096
rect 15046 6980 15098 7096
rect 15316 7044 15368 7096
rect 15580 6980 15632 7096
rect 15850 7044 15902 7096
rect 16114 6980 16166 7096
rect 16384 7044 16436 7096
rect 16648 6980 16700 7096
rect 16918 7044 16970 7096
rect 17182 6980 17234 7096
rect 17452 7044 17504 7096
rect 17716 6980 17768 7096
rect 17986 7044 18038 7096
rect 18250 6980 18302 7096
rect 18520 7044 18572 7096
rect 18784 6980 18836 7096
rect 19054 7044 19106 7096
rect 19318 6980 19370 7096
rect 19588 7044 19640 7096
rect 19852 6980 19904 7096
rect 20122 7044 20174 7096
rect 20386 6980 20438 7096
rect 20656 7044 20708 7096
rect 20920 6980 20972 7096
rect 12732 6849 12784 6965
rect 13266 6852 13318 6968
rect 13800 6852 13852 6968
rect 14334 6852 14386 6968
rect 14868 6852 14920 6968
rect 15402 6852 15454 6968
rect 15936 6852 15988 6968
rect 16470 6852 16522 6968
rect 17004 6852 17056 6968
rect 17538 6852 17590 6968
rect 18072 6852 18124 6968
rect 18606 6852 18658 6968
rect 19140 6852 19192 6968
rect 19674 6852 19726 6968
rect 20208 6852 20260 6968
rect 20742 6852 20794 6968
rect 12428 6732 12480 6741
rect 21046 6732 21098 6741
rect 12428 6698 12437 6732
rect 12437 6698 12471 6732
rect 12471 6698 12480 6732
rect 21046 6698 21055 6732
rect 21055 6698 21089 6732
rect 21089 6698 21098 6732
rect 12428 6689 12480 6698
rect 21046 6689 21098 6698
rect 12619 6333 12671 6385
rect 13153 6333 13205 6385
rect 13687 6333 13739 6385
rect 14221 6333 14273 6385
rect 14755 6333 14807 6385
rect 15289 6333 15341 6385
rect 15823 6333 15875 6385
rect 16357 6333 16409 6385
rect 16891 6333 16943 6385
rect 17425 6333 17477 6385
rect 17959 6333 18011 6385
rect 18493 6333 18545 6385
rect 19027 6333 19079 6385
rect 19561 6333 19613 6385
rect 20095 6333 20147 6385
rect 20629 6333 20681 6385
rect 12554 6066 12606 6182
rect 12732 6170 12784 6286
rect 12910 6066 12962 6182
rect 13088 6066 13140 6182
rect 13266 6173 13318 6289
rect 13444 6066 13496 6182
rect 13622 6066 13674 6182
rect 13800 6173 13852 6289
rect 13978 6066 14030 6182
rect 14156 6066 14208 6182
rect 14334 6173 14386 6289
rect 14512 6066 14564 6182
rect 14690 6066 14742 6182
rect 14868 6173 14920 6289
rect 15046 6066 15098 6182
rect 15224 6066 15276 6182
rect 15402 6173 15454 6289
rect 15580 6066 15632 6182
rect 15758 6066 15810 6182
rect 15936 6173 15988 6289
rect 16114 6066 16166 6182
rect 16292 6066 16344 6182
rect 16470 6173 16522 6289
rect 16648 6066 16700 6182
rect 16826 6066 16878 6182
rect 17004 6173 17056 6289
rect 17182 6066 17234 6182
rect 17360 6066 17412 6182
rect 17538 6173 17590 6289
rect 17716 6066 17768 6182
rect 17894 6066 17946 6182
rect 18072 6173 18124 6289
rect 18250 6066 18302 6182
rect 18428 6066 18480 6182
rect 18606 6173 18658 6289
rect 18784 6066 18836 6182
rect 18962 6066 19014 6182
rect 19140 6173 19192 6289
rect 19318 6066 19370 6182
rect 19496 6066 19548 6182
rect 19674 6173 19726 6289
rect 19852 6066 19904 6182
rect 20030 6066 20082 6182
rect 20208 6173 20260 6289
rect 20386 6066 20438 6182
rect 20564 6066 20616 6182
rect 20742 6173 20794 6289
rect 20920 6066 20972 6182
rect 12732 5316 12784 5432
rect 13266 5319 13318 5435
rect 13800 5319 13852 5435
rect 14334 5319 14386 5435
rect 14868 5319 14920 5435
rect 15402 5319 15454 5435
rect 15936 5319 15988 5435
rect 16470 5319 16522 5435
rect 17004 5319 17056 5435
rect 17538 5319 17590 5435
rect 18072 5319 18124 5435
rect 18606 5319 18658 5435
rect 19140 5319 19192 5435
rect 19674 5319 19726 5435
rect 20208 5319 20260 5435
rect 20742 5319 20794 5435
rect 12476 4950 12592 5002
rect 21198 4952 21330 5084
rect 21405 8023 21531 8075
rect 21405 6689 21531 6741
rect 12476 4616 12592 4626
rect 12476 4582 12592 4616
rect 12476 4574 12592 4582
rect 697 4312 845 4460
rect 14164 4358 14216 4474
rect 14920 4358 14972 4474
rect 15676 4358 15728 4474
rect 16432 4358 16484 4474
rect 26779 4313 26927 4461
rect 13785 -3046 13841 -2990
rect 14541 -3032 14597 -2976
rect 15297 -3046 15353 -2990
rect 16053 -3046 16109 -2990
<< metal2 >>
rect 12546 8659 12610 8665
rect 13080 8659 13144 8665
rect 13614 8659 13678 8665
rect 14148 8659 14212 8665
rect 14682 8659 14746 8665
rect 15216 8659 15280 8665
rect 15750 8659 15814 8665
rect 16284 8659 16348 8665
rect 16818 8659 16882 8665
rect 17352 8659 17416 8665
rect 17886 8659 17950 8665
rect 18420 8659 18484 8665
rect 18954 8659 19018 8665
rect 19488 8659 19552 8665
rect 20022 8659 20086 8665
rect 20556 8659 20620 8665
rect 12546 8607 12552 8659
rect 12604 8607 12610 8659
rect 12546 8601 12610 8607
rect 12701 8653 12765 8659
rect 11968 8077 12116 8086
rect 11968 8021 11977 8077
rect 12107 8021 12116 8077
rect 11968 8012 12116 8021
rect 12421 8077 12495 8086
rect 12421 8021 12430 8077
rect 12486 8021 12495 8077
rect 12421 8012 12495 8021
rect 11466 7358 11530 7364
rect 11466 7347 11472 7358
rect 10856 7341 11472 7347
rect 10856 7289 10862 7341
rect 10978 7289 11472 7341
rect 10856 7283 11472 7289
rect 10717 7208 10781 7214
rect 10717 7092 10723 7208
rect 10775 7092 10781 7208
rect 10717 7086 10781 7092
rect 10984 7203 11058 7212
rect 8618 6399 8692 6408
rect 8618 6269 8627 6399
rect 8683 6269 8692 6399
rect 8618 6260 8692 6269
rect 8752 6399 8826 6408
rect 8752 6269 8761 6399
rect 8817 6269 8826 6399
rect 8752 6260 8826 6269
rect 9108 6399 9182 6408
rect 9108 6269 9117 6399
rect 9173 6269 9182 6399
rect 9108 6260 9182 6269
rect 9464 6399 9538 6408
rect 9464 6269 9473 6399
rect 9529 6269 9538 6399
rect 9464 6260 9538 6269
rect 9820 6399 9894 6408
rect 9820 6269 9829 6399
rect 9885 6269 9894 6399
rect 9820 6260 9894 6269
rect 10176 6399 10250 6408
rect 10176 6269 10185 6399
rect 10241 6269 10250 6399
rect 10176 6260 10250 6269
rect 10532 6399 10606 6408
rect 10532 6269 10541 6399
rect 10597 6269 10606 6399
rect 10532 6260 10606 6269
rect 10718 6153 10776 7086
rect 10984 7073 10993 7203
rect 11049 7117 11058 7203
rect 11114 7201 11188 7212
rect 11114 7117 11125 7201
rect 11049 7075 11125 7117
rect 11177 7075 11188 7201
rect 11049 7073 11188 7075
rect 10984 7064 11188 7073
rect 11275 6539 11331 7283
rect 11466 7242 11472 7283
rect 11524 7242 11530 7358
rect 11466 7236 11530 7242
rect 11663 7213 11727 7219
rect 11663 7161 11669 7213
rect 11721 7161 11727 7213
rect 11663 7155 11727 7161
rect 12172 7135 12246 7144
rect 12172 7005 12181 7135
rect 12237 7005 12246 7135
rect 12172 6996 12246 7005
rect 11602 6880 11750 6889
rect 11602 6824 11611 6880
rect 11741 6824 11750 6880
rect 11602 6815 11750 6824
rect 11968 6743 12116 6752
rect 11968 6687 11977 6743
rect 12107 6687 12116 6743
rect 11968 6678 12116 6687
rect 12417 6743 12491 6752
rect 12417 6687 12426 6743
rect 12482 6687 12491 6743
rect 12417 6678 12491 6687
rect 11242 6533 11370 6539
rect 11242 6481 11248 6533
rect 11364 6481 11370 6533
rect 11242 6475 11370 6481
rect 10888 6399 10962 6408
rect 10888 6269 10897 6399
rect 10953 6269 10962 6399
rect 10888 6260 10962 6269
rect 11244 6399 11318 6408
rect 11244 6269 11253 6399
rect 11309 6269 11318 6399
rect 11244 6260 11318 6269
rect 11600 6399 11674 6408
rect 11600 6269 11609 6399
rect 11665 6269 11674 6399
rect 11600 6260 11674 6269
rect 11734 6399 11808 6408
rect 11734 6269 11743 6399
rect 11799 6269 11808 6399
rect 11734 6260 11808 6269
rect 11916 6399 11990 6408
rect 11916 6269 11925 6399
rect 11981 6269 11990 6399
rect 12552 6391 12608 8601
rect 12701 8581 12707 8653
rect 12664 8537 12707 8581
rect 12759 8537 12765 8653
rect 13080 8607 13086 8659
rect 13138 8607 13144 8659
rect 13080 8601 13144 8607
rect 13235 8653 13299 8659
rect 12664 8531 12765 8537
rect 12664 7951 12720 8531
rect 12661 7945 12725 7951
rect 12661 7893 12667 7945
rect 12719 7893 12725 7945
rect 12661 7887 12725 7893
rect 12899 7104 12973 7113
rect 12640 7098 12704 7102
rect 12899 7098 12908 7104
rect 12640 7096 12908 7098
rect 12640 7044 12646 7096
rect 12698 7044 12908 7096
rect 12640 7042 12908 7044
rect 12640 7038 12704 7042
rect 12899 6974 12908 7042
rect 12964 6974 12973 7104
rect 12726 6965 12790 6971
rect 12899 6965 12973 6974
rect 12726 6849 12732 6965
rect 12784 6849 12790 6965
rect 12726 6843 12790 6849
rect 12552 6385 12677 6391
rect 12552 6333 12619 6385
rect 12671 6333 12677 6385
rect 12552 6327 12677 6333
rect 12730 6292 12786 6843
rect 11916 6260 11990 6269
rect 12726 6286 12790 6292
rect 12548 6182 12612 6188
rect 8930 6144 9078 6153
rect 8930 6014 8939 6144
rect 9069 6014 9078 6144
rect 697 4813 845 4818
rect 693 4675 702 4813
rect 840 4675 849 4813
rect 8930 4809 9078 6014
rect 9286 6144 9360 6153
rect 9286 6014 9295 6144
rect 9351 6014 9360 6144
rect 9286 6005 9360 6014
rect 9642 6144 9716 6153
rect 9642 6014 9651 6144
rect 9707 6014 9716 6144
rect 9642 6005 9716 6014
rect 9998 6144 10072 6153
rect 9998 6014 10007 6144
rect 10063 6014 10072 6144
rect 9998 6005 10072 6014
rect 10354 6144 10428 6153
rect 10354 6014 10363 6144
rect 10419 6014 10428 6144
rect 10354 6005 10428 6014
rect 10710 6144 10784 6153
rect 10710 6014 10719 6144
rect 10775 6014 10784 6144
rect 10710 6005 10784 6014
rect 11066 6144 11140 6153
rect 11066 6014 11075 6144
rect 11131 6014 11140 6144
rect 11066 6005 11140 6014
rect 11422 6144 11496 6153
rect 11422 6014 11431 6144
rect 11487 6014 11496 6144
rect 12548 6066 12554 6182
rect 12606 6116 12612 6182
rect 12726 6170 12732 6286
rect 12784 6170 12790 6286
rect 12908 6188 12964 6965
rect 13086 6391 13142 8601
rect 13235 8581 13241 8653
rect 13198 8537 13241 8581
rect 13293 8537 13299 8653
rect 13614 8607 13620 8659
rect 13672 8607 13678 8659
rect 13614 8601 13678 8607
rect 13769 8653 13833 8659
rect 13198 8531 13299 8537
rect 13198 7951 13254 8531
rect 13195 7945 13259 7951
rect 13195 7893 13201 7945
rect 13253 7893 13259 7945
rect 13195 7887 13259 7893
rect 13433 7104 13507 7113
rect 13174 7098 13238 7102
rect 13433 7098 13442 7104
rect 13174 7096 13442 7098
rect 13174 7044 13180 7096
rect 13232 7044 13442 7096
rect 13174 7042 13442 7044
rect 13174 7038 13238 7042
rect 13433 6974 13442 7042
rect 13498 6974 13507 7104
rect 13260 6968 13324 6974
rect 13260 6852 13266 6968
rect 13318 6852 13324 6968
rect 13433 6965 13507 6974
rect 13260 6846 13324 6852
rect 13086 6385 13211 6391
rect 13086 6333 13153 6385
rect 13205 6333 13211 6385
rect 13086 6327 13211 6333
rect 13264 6295 13320 6846
rect 13260 6289 13324 6295
rect 12726 6164 12790 6170
rect 12904 6182 12968 6188
rect 12904 6116 12910 6182
rect 12606 6066 12910 6116
rect 12962 6066 12968 6182
rect 12548 6060 12968 6066
rect 13082 6182 13146 6188
rect 13082 6066 13088 6182
rect 13140 6116 13146 6182
rect 13260 6173 13266 6289
rect 13318 6173 13324 6289
rect 13442 6188 13498 6965
rect 13620 6391 13676 8601
rect 13769 8581 13775 8653
rect 13732 8537 13775 8581
rect 13827 8537 13833 8653
rect 14148 8607 14154 8659
rect 14206 8607 14212 8659
rect 14148 8601 14212 8607
rect 14303 8653 14367 8659
rect 13732 8531 13833 8537
rect 13732 7951 13788 8531
rect 13729 7945 13793 7951
rect 13729 7893 13735 7945
rect 13787 7893 13793 7945
rect 13729 7887 13793 7893
rect 13967 7104 14041 7113
rect 13708 7098 13772 7102
rect 13967 7098 13976 7104
rect 13708 7096 13976 7098
rect 13708 7044 13714 7096
rect 13766 7044 13976 7096
rect 13708 7042 13976 7044
rect 13708 7038 13772 7042
rect 13967 6974 13976 7042
rect 14032 6974 14041 7104
rect 13794 6968 13858 6974
rect 13794 6852 13800 6968
rect 13852 6852 13858 6968
rect 13967 6965 14041 6974
rect 13794 6846 13858 6852
rect 13620 6385 13745 6391
rect 13620 6333 13687 6385
rect 13739 6333 13745 6385
rect 13620 6327 13745 6333
rect 13798 6295 13854 6846
rect 13794 6289 13858 6295
rect 13260 6167 13324 6173
rect 13438 6182 13502 6188
rect 13438 6116 13444 6182
rect 13140 6066 13444 6116
rect 13496 6066 13502 6182
rect 13082 6060 13502 6066
rect 13616 6182 13680 6188
rect 13616 6066 13622 6182
rect 13674 6116 13680 6182
rect 13794 6173 13800 6289
rect 13852 6173 13858 6289
rect 13976 6188 14032 6965
rect 14154 6391 14210 8601
rect 14303 8581 14309 8653
rect 14266 8537 14309 8581
rect 14361 8537 14367 8653
rect 14682 8607 14688 8659
rect 14740 8607 14746 8659
rect 14682 8601 14746 8607
rect 14837 8653 14901 8659
rect 14266 8531 14367 8537
rect 14266 7951 14322 8531
rect 14263 7945 14327 7951
rect 14263 7893 14269 7945
rect 14321 7893 14327 7945
rect 14263 7887 14327 7893
rect 14501 7104 14575 7113
rect 14242 7098 14306 7102
rect 14501 7098 14510 7104
rect 14242 7096 14510 7098
rect 14242 7044 14248 7096
rect 14300 7044 14510 7096
rect 14242 7042 14510 7044
rect 14242 7038 14306 7042
rect 14501 6974 14510 7042
rect 14566 6974 14575 7104
rect 14328 6968 14392 6974
rect 14328 6852 14334 6968
rect 14386 6852 14392 6968
rect 14501 6965 14575 6974
rect 14328 6846 14392 6852
rect 14154 6385 14279 6391
rect 14154 6333 14221 6385
rect 14273 6333 14279 6385
rect 14154 6327 14279 6333
rect 14332 6295 14388 6846
rect 14328 6289 14392 6295
rect 13794 6167 13858 6173
rect 13972 6182 14036 6188
rect 13972 6116 13978 6182
rect 13674 6066 13978 6116
rect 14030 6066 14036 6182
rect 13616 6060 14036 6066
rect 14150 6182 14214 6188
rect 14150 6066 14156 6182
rect 14208 6116 14214 6182
rect 14328 6173 14334 6289
rect 14386 6173 14392 6289
rect 14510 6188 14566 6965
rect 14688 6391 14744 8601
rect 14837 8581 14843 8653
rect 14800 8537 14843 8581
rect 14895 8537 14901 8653
rect 15216 8607 15222 8659
rect 15274 8607 15280 8659
rect 15216 8601 15280 8607
rect 15371 8653 15435 8659
rect 14800 8531 14901 8537
rect 14800 7951 14856 8531
rect 14797 7945 14861 7951
rect 14797 7893 14803 7945
rect 14855 7893 14861 7945
rect 14797 7887 14861 7893
rect 15035 7104 15109 7113
rect 14776 7098 14840 7102
rect 15035 7098 15044 7104
rect 14776 7096 15044 7098
rect 14776 7044 14782 7096
rect 14834 7044 15044 7096
rect 14776 7042 15044 7044
rect 14776 7038 14840 7042
rect 15035 6974 15044 7042
rect 15100 6974 15109 7104
rect 14862 6968 14926 6974
rect 14862 6852 14868 6968
rect 14920 6852 14926 6968
rect 15035 6965 15109 6974
rect 14862 6846 14926 6852
rect 14688 6385 14813 6391
rect 14688 6333 14755 6385
rect 14807 6333 14813 6385
rect 14688 6327 14813 6333
rect 14866 6295 14922 6846
rect 14862 6289 14926 6295
rect 14328 6167 14392 6173
rect 14506 6182 14570 6188
rect 14506 6116 14512 6182
rect 14208 6066 14512 6116
rect 14564 6066 14570 6182
rect 14150 6060 14570 6066
rect 14684 6182 14748 6188
rect 14684 6066 14690 6182
rect 14742 6116 14748 6182
rect 14862 6173 14868 6289
rect 14920 6173 14926 6289
rect 15044 6188 15100 6965
rect 15222 6391 15278 8601
rect 15371 8581 15377 8653
rect 15334 8537 15377 8581
rect 15429 8537 15435 8653
rect 15750 8607 15756 8659
rect 15808 8607 15814 8659
rect 15750 8601 15814 8607
rect 15905 8653 15969 8659
rect 15334 8531 15435 8537
rect 15334 7951 15390 8531
rect 15331 7945 15395 7951
rect 15331 7893 15337 7945
rect 15389 7893 15395 7945
rect 15331 7887 15395 7893
rect 15569 7104 15643 7113
rect 15310 7098 15374 7102
rect 15569 7098 15578 7104
rect 15310 7096 15578 7098
rect 15310 7044 15316 7096
rect 15368 7044 15578 7096
rect 15310 7042 15578 7044
rect 15310 7038 15374 7042
rect 15569 6974 15578 7042
rect 15634 6974 15643 7104
rect 15396 6968 15460 6974
rect 15396 6852 15402 6968
rect 15454 6852 15460 6968
rect 15569 6965 15643 6974
rect 15396 6846 15460 6852
rect 15222 6385 15347 6391
rect 15222 6333 15289 6385
rect 15341 6333 15347 6385
rect 15222 6327 15347 6333
rect 15400 6295 15456 6846
rect 15396 6289 15460 6295
rect 14862 6167 14926 6173
rect 15040 6182 15104 6188
rect 15040 6116 15046 6182
rect 14742 6066 15046 6116
rect 15098 6066 15104 6182
rect 14684 6060 15104 6066
rect 15218 6182 15282 6188
rect 15218 6066 15224 6182
rect 15276 6116 15282 6182
rect 15396 6173 15402 6289
rect 15454 6173 15460 6289
rect 15578 6188 15634 6965
rect 15756 6391 15812 8601
rect 15905 8581 15911 8653
rect 15868 8537 15911 8581
rect 15963 8537 15969 8653
rect 16284 8607 16290 8659
rect 16342 8607 16348 8659
rect 16284 8601 16348 8607
rect 16439 8653 16503 8659
rect 15868 8531 15969 8537
rect 15868 7951 15924 8531
rect 15865 7945 15929 7951
rect 15865 7893 15871 7945
rect 15923 7893 15929 7945
rect 15865 7887 15929 7893
rect 16103 7104 16177 7113
rect 15844 7098 15908 7102
rect 16103 7098 16112 7104
rect 15844 7096 16112 7098
rect 15844 7044 15850 7096
rect 15902 7044 16112 7096
rect 15844 7042 16112 7044
rect 15844 7038 15908 7042
rect 16103 6974 16112 7042
rect 16168 6974 16177 7104
rect 15930 6968 15994 6974
rect 15930 6852 15936 6968
rect 15988 6852 15994 6968
rect 16103 6965 16177 6974
rect 15930 6846 15994 6852
rect 15756 6385 15881 6391
rect 15756 6333 15823 6385
rect 15875 6333 15881 6385
rect 15756 6327 15881 6333
rect 15934 6295 15990 6846
rect 15930 6289 15994 6295
rect 15396 6167 15460 6173
rect 15574 6182 15638 6188
rect 15574 6116 15580 6182
rect 15276 6066 15580 6116
rect 15632 6066 15638 6182
rect 15218 6060 15638 6066
rect 15752 6182 15816 6188
rect 15752 6066 15758 6182
rect 15810 6116 15816 6182
rect 15930 6173 15936 6289
rect 15988 6173 15994 6289
rect 16112 6188 16168 6965
rect 16290 6391 16346 8601
rect 16439 8581 16445 8653
rect 16402 8537 16445 8581
rect 16497 8537 16503 8653
rect 16818 8607 16824 8659
rect 16876 8607 16882 8659
rect 16818 8601 16882 8607
rect 16973 8653 17037 8659
rect 16402 8531 16503 8537
rect 16402 7951 16458 8531
rect 16399 7945 16463 7951
rect 16399 7893 16405 7945
rect 16457 7893 16463 7945
rect 16399 7887 16463 7893
rect 16637 7104 16711 7113
rect 16378 7098 16442 7102
rect 16637 7098 16646 7104
rect 16378 7096 16646 7098
rect 16378 7044 16384 7096
rect 16436 7044 16646 7096
rect 16378 7042 16646 7044
rect 16378 7038 16442 7042
rect 16637 6974 16646 7042
rect 16702 6974 16711 7104
rect 16464 6968 16528 6974
rect 16464 6852 16470 6968
rect 16522 6852 16528 6968
rect 16637 6965 16711 6974
rect 16464 6846 16528 6852
rect 16290 6385 16415 6391
rect 16290 6333 16357 6385
rect 16409 6333 16415 6385
rect 16290 6327 16415 6333
rect 16468 6295 16524 6846
rect 16464 6289 16528 6295
rect 15930 6167 15994 6173
rect 16108 6182 16172 6188
rect 16108 6116 16114 6182
rect 15810 6066 16114 6116
rect 16166 6066 16172 6182
rect 15752 6060 16172 6066
rect 16286 6182 16350 6188
rect 16286 6066 16292 6182
rect 16344 6116 16350 6182
rect 16464 6173 16470 6289
rect 16522 6173 16528 6289
rect 16646 6188 16702 6965
rect 16824 6391 16880 8601
rect 16973 8581 16979 8653
rect 16936 8537 16979 8581
rect 17031 8537 17037 8653
rect 17352 8607 17358 8659
rect 17410 8607 17416 8659
rect 17352 8601 17416 8607
rect 17507 8653 17571 8659
rect 16936 8531 17037 8537
rect 16936 7951 16992 8531
rect 16933 7945 16997 7951
rect 16933 7893 16939 7945
rect 16991 7893 16997 7945
rect 16933 7887 16997 7893
rect 17171 7104 17245 7113
rect 16912 7098 16976 7102
rect 17171 7098 17180 7104
rect 16912 7096 17180 7098
rect 16912 7044 16918 7096
rect 16970 7044 17180 7096
rect 16912 7042 17180 7044
rect 16912 7038 16976 7042
rect 17171 6974 17180 7042
rect 17236 6974 17245 7104
rect 16998 6968 17062 6974
rect 16998 6852 17004 6968
rect 17056 6852 17062 6968
rect 17171 6965 17245 6974
rect 16998 6846 17062 6852
rect 16824 6385 16949 6391
rect 16824 6333 16891 6385
rect 16943 6333 16949 6385
rect 16824 6327 16949 6333
rect 17002 6295 17058 6846
rect 16998 6289 17062 6295
rect 16464 6167 16528 6173
rect 16642 6182 16706 6188
rect 16642 6116 16648 6182
rect 16344 6066 16648 6116
rect 16700 6066 16706 6182
rect 16286 6060 16706 6066
rect 16820 6182 16884 6188
rect 16820 6066 16826 6182
rect 16878 6116 16884 6182
rect 16998 6173 17004 6289
rect 17056 6173 17062 6289
rect 17180 6188 17236 6965
rect 17358 6391 17414 8601
rect 17507 8581 17513 8653
rect 17470 8537 17513 8581
rect 17565 8537 17571 8653
rect 17886 8607 17892 8659
rect 17944 8607 17950 8659
rect 17886 8601 17950 8607
rect 18041 8653 18105 8659
rect 17470 8531 17571 8537
rect 17470 7951 17526 8531
rect 17467 7945 17531 7951
rect 17467 7893 17473 7945
rect 17525 7893 17531 7945
rect 17467 7887 17531 7893
rect 17705 7104 17779 7113
rect 17446 7098 17510 7102
rect 17705 7098 17714 7104
rect 17446 7096 17714 7098
rect 17446 7044 17452 7096
rect 17504 7044 17714 7096
rect 17446 7042 17714 7044
rect 17446 7038 17510 7042
rect 17705 6974 17714 7042
rect 17770 6974 17779 7104
rect 17532 6968 17596 6974
rect 17532 6852 17538 6968
rect 17590 6852 17596 6968
rect 17705 6965 17779 6974
rect 17532 6846 17596 6852
rect 17358 6385 17483 6391
rect 17358 6333 17425 6385
rect 17477 6333 17483 6385
rect 17358 6327 17483 6333
rect 17536 6295 17592 6846
rect 17532 6289 17596 6295
rect 16998 6167 17062 6173
rect 17176 6182 17240 6188
rect 17176 6116 17182 6182
rect 16878 6066 17182 6116
rect 17234 6066 17240 6182
rect 16820 6060 17240 6066
rect 17354 6182 17418 6188
rect 17354 6066 17360 6182
rect 17412 6116 17418 6182
rect 17532 6173 17538 6289
rect 17590 6173 17596 6289
rect 17714 6188 17770 6965
rect 17892 6391 17948 8601
rect 18041 8581 18047 8653
rect 18004 8537 18047 8581
rect 18099 8537 18105 8653
rect 18420 8607 18426 8659
rect 18478 8607 18484 8659
rect 18420 8601 18484 8607
rect 18575 8653 18639 8659
rect 18004 8531 18105 8537
rect 18004 7951 18060 8531
rect 18001 7945 18065 7951
rect 18001 7893 18007 7945
rect 18059 7893 18065 7945
rect 18001 7887 18065 7893
rect 18239 7104 18313 7113
rect 17980 7098 18044 7102
rect 18239 7098 18248 7104
rect 17980 7096 18248 7098
rect 17980 7044 17986 7096
rect 18038 7044 18248 7096
rect 17980 7042 18248 7044
rect 17980 7038 18044 7042
rect 18239 6974 18248 7042
rect 18304 6974 18313 7104
rect 18066 6968 18130 6974
rect 18066 6852 18072 6968
rect 18124 6852 18130 6968
rect 18239 6965 18313 6974
rect 18066 6846 18130 6852
rect 17892 6385 18017 6391
rect 17892 6333 17959 6385
rect 18011 6333 18017 6385
rect 17892 6327 18017 6333
rect 18070 6295 18126 6846
rect 18066 6289 18130 6295
rect 17532 6167 17596 6173
rect 17710 6182 17774 6188
rect 17710 6116 17716 6182
rect 17412 6066 17716 6116
rect 17768 6066 17774 6182
rect 17354 6060 17774 6066
rect 17888 6182 17952 6188
rect 17888 6066 17894 6182
rect 17946 6116 17952 6182
rect 18066 6173 18072 6289
rect 18124 6173 18130 6289
rect 18248 6188 18304 6965
rect 18426 6391 18482 8601
rect 18575 8581 18581 8653
rect 18538 8537 18581 8581
rect 18633 8537 18639 8653
rect 18954 8607 18960 8659
rect 19012 8607 19018 8659
rect 18954 8601 19018 8607
rect 19109 8653 19173 8659
rect 18538 8531 18639 8537
rect 18538 7951 18594 8531
rect 18535 7945 18599 7951
rect 18535 7893 18541 7945
rect 18593 7893 18599 7945
rect 18535 7887 18599 7893
rect 18773 7104 18847 7113
rect 18514 7098 18578 7102
rect 18773 7098 18782 7104
rect 18514 7096 18782 7098
rect 18514 7044 18520 7096
rect 18572 7044 18782 7096
rect 18514 7042 18782 7044
rect 18514 7038 18578 7042
rect 18773 6974 18782 7042
rect 18838 6974 18847 7104
rect 18600 6968 18664 6974
rect 18600 6852 18606 6968
rect 18658 6852 18664 6968
rect 18773 6965 18847 6974
rect 18600 6846 18664 6852
rect 18426 6385 18551 6391
rect 18426 6333 18493 6385
rect 18545 6333 18551 6385
rect 18426 6327 18551 6333
rect 18604 6295 18660 6846
rect 18600 6289 18664 6295
rect 18066 6167 18130 6173
rect 18244 6182 18308 6188
rect 18244 6116 18250 6182
rect 17946 6066 18250 6116
rect 18302 6066 18308 6182
rect 17888 6060 18308 6066
rect 18422 6182 18486 6188
rect 18422 6066 18428 6182
rect 18480 6116 18486 6182
rect 18600 6173 18606 6289
rect 18658 6173 18664 6289
rect 18782 6188 18838 6965
rect 18960 6391 19016 8601
rect 19109 8581 19115 8653
rect 19072 8537 19115 8581
rect 19167 8537 19173 8653
rect 19488 8607 19494 8659
rect 19546 8607 19552 8659
rect 19488 8601 19552 8607
rect 19643 8653 19707 8659
rect 19072 8531 19173 8537
rect 19072 7951 19128 8531
rect 19069 7945 19133 7951
rect 19069 7893 19075 7945
rect 19127 7893 19133 7945
rect 19069 7887 19133 7893
rect 19307 7104 19381 7113
rect 19048 7098 19112 7102
rect 19307 7098 19316 7104
rect 19048 7096 19316 7098
rect 19048 7044 19054 7096
rect 19106 7044 19316 7096
rect 19048 7042 19316 7044
rect 19048 7038 19112 7042
rect 19307 6974 19316 7042
rect 19372 6974 19381 7104
rect 19134 6968 19198 6974
rect 19134 6852 19140 6968
rect 19192 6852 19198 6968
rect 19307 6965 19381 6974
rect 19134 6846 19198 6852
rect 18960 6385 19085 6391
rect 18960 6333 19027 6385
rect 19079 6333 19085 6385
rect 18960 6327 19085 6333
rect 19138 6295 19194 6846
rect 19134 6289 19198 6295
rect 18600 6167 18664 6173
rect 18778 6182 18842 6188
rect 18778 6116 18784 6182
rect 18480 6066 18784 6116
rect 18836 6066 18842 6182
rect 18422 6060 18842 6066
rect 18956 6182 19020 6188
rect 18956 6066 18962 6182
rect 19014 6116 19020 6182
rect 19134 6173 19140 6289
rect 19192 6173 19198 6289
rect 19316 6188 19372 6965
rect 19494 6391 19550 8601
rect 19643 8581 19649 8653
rect 19606 8537 19649 8581
rect 19701 8537 19707 8653
rect 20022 8607 20028 8659
rect 20080 8607 20086 8659
rect 20022 8601 20086 8607
rect 20177 8653 20241 8659
rect 19606 8531 19707 8537
rect 19606 7951 19662 8531
rect 19603 7945 19667 7951
rect 19603 7893 19609 7945
rect 19661 7893 19667 7945
rect 19603 7887 19667 7893
rect 19841 7104 19915 7113
rect 19582 7098 19646 7102
rect 19841 7098 19850 7104
rect 19582 7096 19850 7098
rect 19582 7044 19588 7096
rect 19640 7044 19850 7096
rect 19582 7042 19850 7044
rect 19582 7038 19646 7042
rect 19841 6974 19850 7042
rect 19906 6974 19915 7104
rect 19668 6968 19732 6974
rect 19668 6852 19674 6968
rect 19726 6852 19732 6968
rect 19841 6965 19915 6974
rect 19668 6846 19732 6852
rect 19494 6385 19619 6391
rect 19494 6333 19561 6385
rect 19613 6333 19619 6385
rect 19494 6327 19619 6333
rect 19672 6295 19728 6846
rect 19668 6289 19732 6295
rect 19134 6167 19198 6173
rect 19312 6182 19376 6188
rect 19312 6116 19318 6182
rect 19014 6066 19318 6116
rect 19370 6066 19376 6182
rect 18956 6060 19376 6066
rect 19490 6182 19554 6188
rect 19490 6066 19496 6182
rect 19548 6116 19554 6182
rect 19668 6173 19674 6289
rect 19726 6173 19732 6289
rect 19850 6188 19906 6965
rect 20028 6391 20084 8601
rect 20177 8581 20183 8653
rect 20140 8537 20183 8581
rect 20235 8537 20241 8653
rect 20556 8607 20562 8659
rect 20614 8607 20620 8659
rect 20556 8601 20620 8607
rect 20711 8653 20775 8659
rect 20140 8531 20241 8537
rect 20140 7951 20196 8531
rect 20137 7945 20201 7951
rect 20137 7893 20143 7945
rect 20195 7893 20201 7945
rect 20137 7887 20201 7893
rect 20375 7104 20449 7113
rect 20116 7098 20180 7102
rect 20375 7098 20384 7104
rect 20116 7096 20384 7098
rect 20116 7044 20122 7096
rect 20174 7044 20384 7096
rect 20116 7042 20384 7044
rect 20116 7038 20180 7042
rect 20375 6974 20384 7042
rect 20440 6974 20449 7104
rect 20202 6968 20266 6974
rect 20202 6852 20208 6968
rect 20260 6852 20266 6968
rect 20375 6965 20449 6974
rect 20202 6846 20266 6852
rect 20028 6385 20153 6391
rect 20028 6333 20095 6385
rect 20147 6333 20153 6385
rect 20028 6327 20153 6333
rect 20206 6295 20262 6846
rect 20202 6289 20266 6295
rect 19668 6167 19732 6173
rect 19846 6182 19910 6188
rect 19846 6116 19852 6182
rect 19548 6066 19852 6116
rect 19904 6066 19910 6182
rect 19490 6060 19910 6066
rect 20024 6182 20088 6188
rect 20024 6066 20030 6182
rect 20082 6116 20088 6182
rect 20202 6173 20208 6289
rect 20260 6173 20266 6289
rect 20384 6188 20440 6965
rect 20562 6391 20618 8601
rect 20711 8581 20717 8653
rect 20674 8537 20717 8581
rect 20769 8537 20775 8653
rect 20674 8531 20775 8537
rect 20674 7951 20730 8531
rect 21035 8077 21109 8086
rect 21035 8021 21044 8077
rect 21100 8021 21109 8077
rect 21035 8012 21109 8021
rect 21394 8077 21542 8086
rect 21394 8021 21403 8077
rect 21533 8021 21542 8077
rect 21394 8012 21542 8021
rect 20671 7945 20735 7951
rect 20671 7893 20677 7945
rect 20729 7893 20735 7945
rect 20671 7887 20735 7893
rect 20909 7104 20983 7113
rect 20650 7098 20714 7102
rect 20909 7098 20918 7104
rect 20650 7096 20918 7098
rect 20650 7044 20656 7096
rect 20708 7044 20918 7096
rect 20650 7042 20918 7044
rect 20650 7038 20714 7042
rect 20909 6974 20918 7042
rect 20974 6974 20983 7104
rect 20736 6968 20800 6974
rect 20736 6852 20742 6968
rect 20794 6852 20800 6968
rect 20909 6965 20983 6974
rect 20736 6846 20800 6852
rect 20562 6385 20687 6391
rect 20562 6333 20629 6385
rect 20681 6333 20687 6385
rect 20562 6327 20687 6333
rect 20740 6295 20796 6846
rect 20736 6289 20800 6295
rect 20202 6167 20266 6173
rect 20380 6182 20444 6188
rect 20380 6116 20386 6182
rect 20082 6066 20386 6116
rect 20438 6066 20444 6182
rect 20024 6060 20444 6066
rect 20558 6182 20622 6188
rect 20558 6066 20564 6182
rect 20616 6116 20622 6182
rect 20736 6173 20742 6289
rect 20794 6173 20800 6289
rect 20918 6188 20974 6965
rect 21035 6743 21109 6752
rect 21035 6687 21044 6743
rect 21100 6687 21109 6743
rect 21035 6678 21109 6687
rect 21394 6743 21542 6752
rect 21394 6687 21403 6743
rect 21533 6687 21542 6743
rect 21394 6678 21542 6687
rect 20736 6167 20800 6173
rect 20914 6182 20978 6188
rect 20914 6116 20920 6182
rect 20616 6066 20920 6116
rect 20972 6066 20978 6182
rect 20558 6060 20978 6066
rect 11422 6005 11496 6014
rect 15401 5695 15457 5702
rect 19669 5695 19729 5704
rect 15399 5693 15459 5695
rect 15399 5637 15401 5693
rect 15457 5637 15459 5693
rect 14866 5544 14922 5551
rect 14864 5542 14924 5544
rect 14864 5486 14866 5542
rect 14922 5486 14924 5542
rect 14864 5441 14924 5486
rect 15399 5441 15459 5637
rect 19669 5626 19729 5635
rect 19138 5544 19198 5553
rect 19138 5475 19198 5484
rect 19140 5441 19196 5475
rect 19671 5441 19727 5626
rect 12726 5432 12790 5438
rect 12726 5316 12732 5432
rect 12784 5316 12790 5432
rect 12726 5310 12790 5316
rect 13260 5435 13324 5441
rect 13260 5319 13266 5435
rect 13318 5319 13324 5435
rect 13260 5313 13324 5319
rect 13794 5435 13858 5441
rect 13794 5319 13800 5435
rect 13852 5319 13858 5435
rect 13794 5313 13858 5319
rect 14328 5435 14392 5441
rect 14328 5319 14334 5435
rect 14386 5319 14392 5435
rect 14328 5313 14392 5319
rect 14862 5435 14926 5441
rect 14862 5319 14868 5435
rect 14920 5319 14926 5435
rect 14862 5313 14926 5319
rect 15396 5435 15460 5441
rect 15396 5319 15402 5435
rect 15454 5319 15460 5435
rect 15396 5313 15460 5319
rect 15930 5435 15994 5441
rect 15930 5319 15936 5435
rect 15988 5319 15994 5435
rect 15930 5313 15994 5319
rect 16464 5435 16528 5441
rect 16464 5319 16470 5435
rect 16522 5319 16528 5435
rect 16464 5313 16528 5319
rect 16998 5435 17062 5441
rect 16998 5319 17004 5435
rect 17056 5319 17062 5435
rect 16998 5313 17062 5319
rect 17532 5435 17596 5441
rect 17532 5319 17538 5435
rect 17590 5319 17596 5435
rect 17532 5313 17596 5319
rect 18066 5435 18130 5441
rect 18066 5319 18072 5435
rect 18124 5319 18130 5435
rect 18066 5313 18130 5319
rect 18600 5435 18664 5441
rect 18600 5319 18606 5435
rect 18658 5319 18664 5435
rect 18600 5313 18664 5319
rect 19134 5435 19198 5441
rect 19134 5319 19140 5435
rect 19192 5319 19198 5435
rect 19134 5313 19198 5319
rect 19668 5435 19732 5441
rect 19668 5319 19674 5435
rect 19726 5319 19732 5435
rect 19668 5313 19732 5319
rect 20202 5435 20266 5441
rect 20202 5319 20208 5435
rect 20260 5319 20266 5435
rect 20202 5313 20266 5319
rect 20736 5435 20800 5441
rect 20736 5319 20742 5435
rect 20794 5319 20800 5435
rect 20736 5313 20800 5319
rect 12727 5276 12786 5310
rect 12783 5220 12786 5276
rect 12727 5211 12786 5220
rect 8930 4679 8939 4809
rect 9069 4679 9078 4809
rect 697 4460 845 4675
rect 8930 4670 9078 4679
rect 12470 5002 12598 5008
rect 12470 4950 12476 5002
rect 12592 4950 12598 5002
rect 12470 4626 12598 4950
rect 12470 4574 12476 4626
rect 12592 4574 12598 4626
rect 12470 4568 12598 4574
rect 12730 4519 12786 5211
rect 13264 5145 13320 5313
rect 13263 5136 13320 5145
rect 13319 5080 13320 5136
rect 13263 5071 13320 5080
rect 13264 4653 13320 5071
rect 13798 5010 13854 5313
rect 13798 5001 13855 5010
rect 13798 4945 13799 5001
rect 13798 4936 13855 4945
rect 13798 4784 13854 4936
rect 14332 4920 14388 5313
rect 14866 5036 14922 5313
rect 15400 5268 15456 5313
rect 15404 5179 15455 5268
rect 15935 5229 15991 5313
rect 16466 5251 16522 5313
rect 17003 5278 17059 5313
rect 15404 5128 15726 5179
rect 15935 5173 16109 5229
rect 14866 4980 15355 5036
rect 14332 4864 14977 4920
rect 14976 4808 14977 4864
rect 14920 4799 14977 4808
rect 13798 4728 14597 4784
rect 13264 4597 14219 4653
rect 12730 4463 13841 4519
rect 697 4306 845 4312
rect 13785 -2990 13841 4463
rect 14158 4480 14219 4597
rect 14158 4474 14222 4480
rect 14158 4358 14164 4474
rect 14216 4358 14222 4474
rect 14158 4352 14222 4358
rect 14541 -2976 14597 4728
rect 14921 4480 14977 4799
rect 15299 4481 15355 4980
rect 14914 4474 14978 4480
rect 14914 4358 14920 4474
rect 14972 4358 14978 4474
rect 14914 4352 14978 4358
rect 15297 4402 15355 4481
rect 15675 4480 15726 5128
rect 16053 4714 16109 5173
rect 16052 4705 16109 4714
rect 16108 4649 16109 4705
rect 16052 4640 16109 4649
rect 15670 4474 15734 4480
rect 14541 -3038 14597 -3032
rect 15297 -2990 15353 4402
rect 15670 4358 15676 4474
rect 15728 4358 15734 4474
rect 15670 4352 15734 4358
rect 13785 -3052 13841 -3046
rect 15297 -3052 15353 -3046
rect 16053 -2990 16109 4640
rect 16431 5199 16522 5251
rect 16992 5218 17001 5278
rect 17061 5218 17070 5278
rect 16431 4567 16483 5199
rect 17538 5147 17594 5313
rect 17536 5138 17596 5147
rect 17536 5069 17596 5078
rect 18067 5012 18123 5313
rect 18065 5003 18125 5012
rect 18065 4934 18125 4943
rect 18604 4875 18660 5313
rect 19140 5220 19196 5313
rect 19671 5220 19727 5313
rect 18602 4866 18662 4875
rect 18602 4797 18662 4806
rect 20206 4716 20262 5313
rect 20204 4707 20264 4716
rect 20204 4638 20264 4647
rect 20740 4569 20796 5313
rect 21190 5084 21338 5092
rect 21190 4952 21198 5084
rect 21330 4952 21338 5084
rect 21190 4827 21338 4952
rect 26784 4836 26922 4840
rect 21190 4697 21199 4827
rect 21329 4697 21338 4827
rect 21190 4688 21338 4697
rect 26779 4831 26927 4836
rect 26779 4693 26784 4831
rect 26922 4693 26927 4831
rect 16431 4558 16487 4567
rect 16431 4480 16487 4502
rect 20738 4560 20798 4569
rect 20738 4491 20798 4500
rect 16426 4474 16490 4480
rect 16426 4358 16432 4474
rect 16484 4358 16490 4474
rect 16426 4352 16490 4358
rect 26779 4461 26927 4693
rect 26779 4307 26927 4313
rect 16053 -3052 16109 -3046
<< via2 >>
rect 11977 8075 12107 8077
rect 11977 8023 11979 8075
rect 11979 8023 12105 8075
rect 12105 8023 12107 8075
rect 11977 8021 12107 8023
rect 12430 8075 12486 8077
rect 12430 8023 12432 8075
rect 12432 8023 12484 8075
rect 12484 8023 12486 8075
rect 12430 8021 12486 8023
rect 8627 6397 8683 6399
rect 8627 6271 8629 6397
rect 8629 6271 8681 6397
rect 8681 6271 8683 6397
rect 8627 6269 8683 6271
rect 8761 6397 8817 6399
rect 8761 6271 8763 6397
rect 8763 6271 8815 6397
rect 8815 6271 8817 6397
rect 8761 6269 8817 6271
rect 9117 6397 9173 6399
rect 9117 6271 9119 6397
rect 9119 6271 9171 6397
rect 9171 6271 9173 6397
rect 9117 6269 9173 6271
rect 9473 6397 9529 6399
rect 9473 6271 9475 6397
rect 9475 6271 9527 6397
rect 9527 6271 9529 6397
rect 9473 6269 9529 6271
rect 9829 6397 9885 6399
rect 9829 6271 9831 6397
rect 9831 6271 9883 6397
rect 9883 6271 9885 6397
rect 9829 6269 9885 6271
rect 10185 6397 10241 6399
rect 10185 6271 10187 6397
rect 10187 6271 10239 6397
rect 10239 6271 10241 6397
rect 10185 6269 10241 6271
rect 10541 6397 10597 6399
rect 10541 6271 10543 6397
rect 10543 6271 10595 6397
rect 10595 6271 10597 6397
rect 10541 6269 10597 6271
rect 10993 7201 11049 7203
rect 10993 7075 10995 7201
rect 10995 7075 11047 7201
rect 11047 7075 11049 7201
rect 10993 7073 11049 7075
rect 12181 7133 12237 7135
rect 12181 7007 12183 7133
rect 12183 7007 12235 7133
rect 12235 7007 12237 7133
rect 12181 7005 12237 7007
rect 11611 6878 11741 6880
rect 11611 6826 11613 6878
rect 11613 6826 11739 6878
rect 11739 6826 11741 6878
rect 11611 6824 11741 6826
rect 11977 6741 12107 6743
rect 11977 6689 11979 6741
rect 11979 6689 12105 6741
rect 12105 6689 12107 6741
rect 11977 6687 12107 6689
rect 12426 6741 12482 6743
rect 12426 6689 12428 6741
rect 12428 6689 12480 6741
rect 12480 6689 12482 6741
rect 12426 6687 12482 6689
rect 10897 6397 10953 6399
rect 10897 6271 10899 6397
rect 10899 6271 10951 6397
rect 10951 6271 10953 6397
rect 10897 6269 10953 6271
rect 11253 6397 11309 6399
rect 11253 6271 11255 6397
rect 11255 6271 11307 6397
rect 11307 6271 11309 6397
rect 11253 6269 11309 6271
rect 11609 6397 11665 6399
rect 11609 6271 11611 6397
rect 11611 6271 11663 6397
rect 11663 6271 11665 6397
rect 11609 6269 11665 6271
rect 11743 6397 11799 6399
rect 11743 6271 11745 6397
rect 11745 6271 11797 6397
rect 11797 6271 11799 6397
rect 11743 6269 11799 6271
rect 11925 6397 11981 6399
rect 11925 6271 11927 6397
rect 11927 6271 11979 6397
rect 11979 6271 11981 6397
rect 11925 6269 11981 6271
rect 12908 7096 12964 7104
rect 12908 6980 12910 7096
rect 12910 6980 12962 7096
rect 12962 6980 12964 7096
rect 12908 6974 12964 6980
rect 8939 6142 9069 6144
rect 8939 6016 8941 6142
rect 8941 6016 8993 6142
rect 8993 6016 9069 6142
rect 8939 6014 9069 6016
rect 702 4675 840 4813
rect 9295 6142 9351 6144
rect 9295 6016 9297 6142
rect 9297 6016 9349 6142
rect 9349 6016 9351 6142
rect 9295 6014 9351 6016
rect 9651 6142 9707 6144
rect 9651 6016 9653 6142
rect 9653 6016 9705 6142
rect 9705 6016 9707 6142
rect 9651 6014 9707 6016
rect 10007 6142 10063 6144
rect 10007 6016 10009 6142
rect 10009 6016 10061 6142
rect 10061 6016 10063 6142
rect 10007 6014 10063 6016
rect 10363 6142 10419 6144
rect 10363 6016 10365 6142
rect 10365 6016 10417 6142
rect 10417 6016 10419 6142
rect 10363 6014 10419 6016
rect 10719 6142 10775 6144
rect 10719 6016 10721 6142
rect 10721 6016 10773 6142
rect 10773 6016 10775 6142
rect 10719 6014 10775 6016
rect 11075 6142 11131 6144
rect 11075 6016 11077 6142
rect 11077 6016 11129 6142
rect 11129 6016 11131 6142
rect 11075 6014 11131 6016
rect 11431 6142 11487 6144
rect 11431 6016 11433 6142
rect 11433 6016 11485 6142
rect 11485 6016 11487 6142
rect 11431 6014 11487 6016
rect 13442 7096 13498 7104
rect 13442 6980 13444 7096
rect 13444 6980 13496 7096
rect 13496 6980 13498 7096
rect 13442 6974 13498 6980
rect 13976 7096 14032 7104
rect 13976 6980 13978 7096
rect 13978 6980 14030 7096
rect 14030 6980 14032 7096
rect 13976 6974 14032 6980
rect 14510 7096 14566 7104
rect 14510 6980 14512 7096
rect 14512 6980 14564 7096
rect 14564 6980 14566 7096
rect 14510 6974 14566 6980
rect 15044 7096 15100 7104
rect 15044 6980 15046 7096
rect 15046 6980 15098 7096
rect 15098 6980 15100 7096
rect 15044 6974 15100 6980
rect 15578 7096 15634 7104
rect 15578 6980 15580 7096
rect 15580 6980 15632 7096
rect 15632 6980 15634 7096
rect 15578 6974 15634 6980
rect 16112 7096 16168 7104
rect 16112 6980 16114 7096
rect 16114 6980 16166 7096
rect 16166 6980 16168 7096
rect 16112 6974 16168 6980
rect 16646 7096 16702 7104
rect 16646 6980 16648 7096
rect 16648 6980 16700 7096
rect 16700 6980 16702 7096
rect 16646 6974 16702 6980
rect 17180 7096 17236 7104
rect 17180 6980 17182 7096
rect 17182 6980 17234 7096
rect 17234 6980 17236 7096
rect 17180 6974 17236 6980
rect 17714 7096 17770 7104
rect 17714 6980 17716 7096
rect 17716 6980 17768 7096
rect 17768 6980 17770 7096
rect 17714 6974 17770 6980
rect 18248 7096 18304 7104
rect 18248 6980 18250 7096
rect 18250 6980 18302 7096
rect 18302 6980 18304 7096
rect 18248 6974 18304 6980
rect 18782 7096 18838 7104
rect 18782 6980 18784 7096
rect 18784 6980 18836 7096
rect 18836 6980 18838 7096
rect 18782 6974 18838 6980
rect 19316 7096 19372 7104
rect 19316 6980 19318 7096
rect 19318 6980 19370 7096
rect 19370 6980 19372 7096
rect 19316 6974 19372 6980
rect 19850 7096 19906 7104
rect 19850 6980 19852 7096
rect 19852 6980 19904 7096
rect 19904 6980 19906 7096
rect 19850 6974 19906 6980
rect 20384 7096 20440 7104
rect 20384 6980 20386 7096
rect 20386 6980 20438 7096
rect 20438 6980 20440 7096
rect 20384 6974 20440 6980
rect 21044 8075 21100 8077
rect 21044 8023 21046 8075
rect 21046 8023 21098 8075
rect 21098 8023 21100 8075
rect 21044 8021 21100 8023
rect 21403 8075 21533 8077
rect 21403 8023 21405 8075
rect 21405 8023 21531 8075
rect 21531 8023 21533 8075
rect 21403 8021 21533 8023
rect 20918 7096 20974 7104
rect 20918 6980 20920 7096
rect 20920 6980 20972 7096
rect 20972 6980 20974 7096
rect 20918 6974 20974 6980
rect 21044 6741 21100 6743
rect 21044 6689 21046 6741
rect 21046 6689 21098 6741
rect 21098 6689 21100 6741
rect 21044 6687 21100 6689
rect 21403 6741 21533 6743
rect 21403 6689 21405 6741
rect 21405 6689 21531 6741
rect 21531 6689 21533 6741
rect 21403 6687 21533 6689
rect 15401 5637 15457 5693
rect 14866 5486 14922 5542
rect 19669 5635 19729 5695
rect 19138 5484 19198 5544
rect 12727 5220 12783 5276
rect 8939 4679 9069 4809
rect 13263 5080 13319 5136
rect 13799 4945 13855 5001
rect 14920 4808 14976 4864
rect 16052 4649 16108 4705
rect 17001 5218 17061 5278
rect 17536 5078 17596 5138
rect 18065 4943 18125 5003
rect 18602 4806 18662 4866
rect 20204 4647 20264 4707
rect 21199 4697 21329 4827
rect 26784 4693 26922 4831
rect 16431 4502 16487 4558
rect 20738 4500 20798 4560
<< metal3 >>
rect 11968 8077 12495 8086
rect 11968 8021 11977 8077
rect 12107 8021 12430 8077
rect 12486 8021 12495 8077
rect 11968 8012 12495 8021
rect 21035 8077 21542 8086
rect 21035 8021 21044 8077
rect 21100 8021 21403 8077
rect 21533 8021 21542 8077
rect 21035 8012 21542 8021
rect 10984 7203 11058 7212
rect 10984 7073 10993 7203
rect 11049 7093 11058 7203
rect 12172 7135 12246 7144
rect 12172 7093 12181 7135
rect 11049 7073 12181 7093
rect 10984 7033 12181 7073
rect 11650 6889 11710 7033
rect 12172 7005 12181 7033
rect 12237 7005 12246 7135
rect 12172 6996 12246 7005
rect 12899 7104 12973 7113
rect 12899 6974 12908 7104
rect 12964 7066 12973 7104
rect 13433 7104 13507 7113
rect 13433 7066 13442 7104
rect 12964 7006 13442 7066
rect 12964 6974 12973 7006
rect 12899 6965 12973 6974
rect 13433 6974 13442 7006
rect 13498 7066 13507 7104
rect 13967 7104 14041 7113
rect 13967 7066 13976 7104
rect 13498 7006 13976 7066
rect 13498 6974 13507 7006
rect 13433 6965 13507 6974
rect 13967 6974 13976 7006
rect 14032 7066 14041 7104
rect 14501 7104 14575 7113
rect 14501 7066 14510 7104
rect 14032 7006 14510 7066
rect 14032 6974 14041 7006
rect 13967 6965 14041 6974
rect 14501 6974 14510 7006
rect 14566 7066 14575 7104
rect 15035 7104 15109 7113
rect 15035 7066 15044 7104
rect 14566 7006 15044 7066
rect 14566 6974 14575 7006
rect 14501 6965 14575 6974
rect 15035 6974 15044 7006
rect 15100 7066 15109 7104
rect 15569 7104 15643 7113
rect 15569 7066 15578 7104
rect 15100 7006 15578 7066
rect 15100 6974 15109 7006
rect 15035 6965 15109 6974
rect 15569 6974 15578 7006
rect 15634 7066 15643 7104
rect 16103 7104 16177 7113
rect 16103 7066 16112 7104
rect 15634 7006 16112 7066
rect 15634 6974 15643 7006
rect 15569 6965 15643 6974
rect 16103 6974 16112 7006
rect 16168 7066 16177 7104
rect 16637 7104 16711 7113
rect 16637 7066 16646 7104
rect 16168 7006 16646 7066
rect 16168 6974 16177 7006
rect 16103 6965 16177 6974
rect 16637 6974 16646 7006
rect 16702 6974 16711 7104
rect 16637 6965 16711 6974
rect 17171 7104 17245 7113
rect 17171 6974 17180 7104
rect 17236 7066 17245 7104
rect 17705 7104 17779 7113
rect 17705 7066 17714 7104
rect 17236 7006 17714 7066
rect 17236 6974 17245 7006
rect 17171 6965 17245 6974
rect 17705 6974 17714 7006
rect 17770 7066 17779 7104
rect 18239 7104 18313 7113
rect 18239 7066 18248 7104
rect 17770 7006 18248 7066
rect 17770 6974 17779 7006
rect 17705 6965 17779 6974
rect 18239 6974 18248 7006
rect 18304 7066 18313 7104
rect 18773 7104 18847 7113
rect 18773 7066 18782 7104
rect 18304 7006 18782 7066
rect 18304 6974 18313 7006
rect 18239 6965 18313 6974
rect 18773 6974 18782 7006
rect 18838 7066 18847 7104
rect 19307 7104 19381 7113
rect 19307 7066 19316 7104
rect 18838 7006 19316 7066
rect 18838 6974 18847 7006
rect 18773 6965 18847 6974
rect 19307 6974 19316 7006
rect 19372 7066 19381 7104
rect 19841 7104 19915 7113
rect 19841 7066 19850 7104
rect 19372 7006 19850 7066
rect 19372 6974 19381 7006
rect 19307 6965 19381 6974
rect 19841 6974 19850 7006
rect 19906 7066 19915 7104
rect 20375 7104 20449 7113
rect 20375 7066 20384 7104
rect 19906 7006 20384 7066
rect 19906 6974 19915 7006
rect 19841 6965 19915 6974
rect 20375 6974 20384 7006
rect 20440 7066 20449 7104
rect 20909 7104 20983 7113
rect 20909 7066 20918 7104
rect 20440 7006 20918 7066
rect 20440 6974 20449 7006
rect 20375 6965 20449 6974
rect 20909 6974 20918 7006
rect 20974 6974 20983 7104
rect 20909 6965 20983 6974
rect 11602 6880 11750 6889
rect 11602 6824 11611 6880
rect 11741 6824 11750 6880
rect 11602 6815 11750 6824
rect 11968 6743 12491 6752
rect 11968 6687 11977 6743
rect 12107 6687 12426 6743
rect 12482 6687 12491 6743
rect 11968 6678 12491 6687
rect 21035 6743 21542 6752
rect 21035 6687 21044 6743
rect 21100 6687 21403 6743
rect 21533 6687 21542 6743
rect 21035 6678 21542 6687
rect 8618 6399 11990 6408
rect 8618 6269 8627 6399
rect 8683 6269 8761 6399
rect 8817 6269 9117 6399
rect 9173 6269 9473 6399
rect 9529 6269 9829 6399
rect 9885 6269 10185 6399
rect 10241 6269 10541 6399
rect 10597 6269 10897 6399
rect 10953 6269 11253 6399
rect 11309 6269 11609 6399
rect 11665 6269 11743 6399
rect 11799 6269 11925 6399
rect 11981 6269 11990 6399
rect 8618 6260 11990 6269
rect 8930 6144 11496 6153
rect 8930 6014 8939 6144
rect 9069 6014 9295 6144
rect 9351 6014 9651 6144
rect 9707 6014 10007 6144
rect 10063 6014 10363 6144
rect 10419 6014 10719 6144
rect 10775 6014 11075 6144
rect 11131 6014 11431 6144
rect 11487 6014 11496 6144
rect 8930 6005 11496 6014
rect 15396 5695 15462 5698
rect 19664 5695 19734 5700
rect 15396 5693 19669 5695
rect 15396 5637 15401 5693
rect 15457 5637 19669 5693
rect 15396 5635 19669 5637
rect 19729 5635 19734 5695
rect 15396 5632 15462 5635
rect 19664 5630 19734 5635
rect 14861 5544 14927 5547
rect 19133 5544 19203 5549
rect 14861 5542 19138 5544
rect 14861 5486 14866 5542
rect 14922 5486 19138 5542
rect 14861 5484 19138 5486
rect 19198 5484 19203 5544
rect 14861 5481 14927 5484
rect 19133 5479 19203 5484
rect 12722 5278 12788 5281
rect 16996 5278 17066 5283
rect 12722 5276 17001 5278
rect 12722 5220 12727 5276
rect 12783 5220 17001 5276
rect 12722 5218 17001 5220
rect 17061 5218 17066 5278
rect 12722 5215 12788 5218
rect 16996 5213 17066 5218
rect 13258 5138 13324 5141
rect 17531 5138 17601 5143
rect 13258 5136 17536 5138
rect 13258 5080 13263 5136
rect 13319 5080 17536 5136
rect 13258 5078 17536 5080
rect 17596 5078 17601 5138
rect 13258 5075 13324 5078
rect 17531 5073 17601 5078
rect 13794 5003 13860 5006
rect 18060 5003 18130 5008
rect 13794 5001 18065 5003
rect 13794 4945 13799 5001
rect 13855 4945 18065 5001
rect 13794 4943 18065 4945
rect 18125 4943 18130 5003
rect 13794 4940 13860 4943
rect 18060 4938 18130 4943
rect 14915 4866 14981 4869
rect 18597 4866 18667 4871
rect 14915 4864 18602 4866
rect 697 4813 9078 4818
rect 697 4675 702 4813
rect 840 4809 9078 4813
rect 840 4679 8939 4809
rect 9069 4679 9078 4809
rect 14915 4808 14920 4864
rect 14976 4808 18602 4864
rect 14915 4806 18602 4808
rect 18662 4806 18667 4866
rect 14915 4803 14981 4806
rect 18597 4801 18667 4806
rect 21190 4831 26927 4836
rect 21190 4827 26784 4831
rect 840 4675 9078 4679
rect 697 4670 9078 4675
rect 16047 4707 16113 4710
rect 20199 4707 20269 4712
rect 16047 4705 20204 4707
rect 16047 4649 16052 4705
rect 16108 4649 20204 4705
rect 16047 4647 20204 4649
rect 20264 4647 20269 4707
rect 21190 4697 21199 4827
rect 21329 4697 26784 4827
rect 21190 4693 26784 4697
rect 26922 4693 26927 4831
rect 21190 4688 26927 4693
rect 16047 4644 16113 4647
rect 20199 4642 20269 4647
rect 16426 4560 16492 4563
rect 20733 4560 20803 4565
rect 16426 4558 20738 4560
rect 16426 4502 16431 4558
rect 16487 4502 20738 4558
rect 16426 4500 20738 4502
rect 20798 4500 20803 4560
rect 16426 4497 16492 4500
rect 20733 4495 20803 4500
use sky130_fd_pr__nfet_g5v0d10v5_CD9S2Z  sky130_fd_pr__nfet_g5v0d10v5_CD9S2Z_0
timestamp 1712467038
transform 1 0 10888 0 1 7151
box -328 -358 328 358
use sky130_fd_pr__nfet_g5v0d10v5_K8JYEQ  sky130_fd_pr__nfet_g5v0d10v5_K8JYEQ_0
timestamp 1712467038
transform 1 0 16763 0 1 5826
box -4382 -727 4382 727
use sky130_fd_pr__pfet_g5v0d10v5_4Z8MHY  sky130_fd_pr__pfet_g5v0d10v5_4Z8MHY_0
timestamp 1712467038
transform 1 0 16763 0 1 7382
box -4412 -762 4412 762
use sky130_fd_pr__pfet_g5v0d10v5_WY4TLZ  sky130_fd_pr__pfet_g5v0d10v5_WY4TLZ_0
timestamp 1712467038
transform 1 0 10213 0 1 5970
box -1653 -762 1653 762
use sky130_fd_pr__res_xhigh_po_1p41_9VZRJ2  sky130_fd_pr__res_xhigh_po_1p41_9VZRJ2_0
timestamp 1712594819
transform 1 0 13812 0 1 570
box -13348 -4082 13348 4082
use sky130_fd_sc_hvl__inv_1  sky130_fd_sc_hvl__inv_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
array 0 15 534 0 0 0
timestamp 1707688321
transform 1 0 12499 0 1 8285
box -66 -43 354 897
use sky130_fd_sc_hvl__inv_1  sky130_fd_sc_hvl__inv_1_1
timestamp 1707688321
transform -1 0 11750 0 1 6838
box -66 -43 354 897
<< labels >>
flabel metal2 s 12546 8665 12546 8665 0 FreeSans 240 0 0 0 otrip_decoded_avdd[0]
port 11 nsew
flabel metal2 s 13080 8665 13080 8665 0 FreeSans 240 0 0 0 otrip_decoded_avdd[1]
port 10 nsew
flabel metal2 s 13614 8665 13614 8665 0 FreeSans 240 0 0 0 otrip_decoded_avdd[2]
port 9 nsew
flabel metal2 s 14148 8665 14148 8665 0 FreeSans 240 0 0 0 otrip_decoded_avdd[3]
port 8 nsew
flabel metal2 s 14682 8665 14682 8665 0 FreeSans 240 0 0 0 otrip_decoded_avdd[4]
port 7 nsew
flabel metal2 s 15216 8665 15216 8665 0 FreeSans 240 0 0 0 otrip_decoded_avdd[5]
port 6 nsew
flabel metal2 s 15750 8665 15750 8665 0 FreeSans 240 0 0 0 otrip_decoded_avdd[6]
port 5 nsew
flabel metal2 s 12765 8531 12765 8531 0 FreeSans 160 0 0 0 otrip_decoded_b_avdd[0]
flabel metal2 s 13299 8531 13299 8531 0 FreeSans 160 0 0 0 otrip_decoded_b_avdd[1]
flabel metal2 s 13833 8531 13833 8531 0 FreeSans 160 0 0 0 otrip_decoded_b_avdd[2]
flabel metal2 s 14367 8531 14367 8531 0 FreeSans 160 0 0 0 otrip_decoded_b_avdd[3]
flabel metal2 s 14901 8531 14901 8531 0 FreeSans 160 0 0 0 otrip_decoded_b_avdd[4]
flabel metal2 s 15435 8531 15435 8531 0 FreeSans 160 0 0 0 otrip_decoded_b_avdd[5]
flabel metal2 s 15969 8531 15969 8531 0 FreeSans 160 0 0 0 otrip_decoded_b_avdd[6]
flabel metal1 s 14142 4480 14142 4480 0 FreeSans 800 0 0 0 vtrip1
flabel metal1 s 14898 4480 14898 4480 0 FreeSans 800 0 0 0 vtrip3
flabel metal1 s 15654 4480 15654 4480 0 FreeSans 800 0 0 0 vtrip5
flabel metal1 s 16410 4480 16410 4480 0 FreeSans 800 0 0 0 vtrip7
flabel metal1 s 12172 8410 12172 8410 0 FreeSans 1200 0 0 0 avss
port 21 nsew
flabel metal1 s 11916 9122 11916 9122 0 FreeSans 1200 0 0 0 avdd
port 1 nsew
flabel metal2 s 11727 7219 11727 7219 0 FreeSans 1200 0 0 0 ena
port 3 nsew
flabel metal2 s 11274 7347 11274 7347 0 FreeSans 800 0 0 0 ena_b
flabel metal2 s 16284 8665 16284 8665 0 FreeSans 240 0 0 0 otrip_decoded_avdd[7]
port 4 nsew
flabel metal2 s 16503 8531 16503 8531 0 FreeSans 160 0 0 0 otrip_decoded_b_avdd[7]
flabel metal1 s 14001 -3130 14001 -3130 0 FreeSans 800 0 0 0 vtrip0
flabel metal1 s 14757 -3130 14757 -3130 0 FreeSans 800 0 0 0 vtrip2
flabel metal1 s 15513 -3130 15513 -3130 0 FreeSans 800 0 0 0 vtrip4
flabel metal1 s 16269 -3130 16269 -3130 0 FreeSans 800 0 0 0 vtrip6
flabel metal2 16818 8665 16818 8665 0 FreeSans 240 0 0 0 vtrip_decoded_avdd[0]
port 19 nsew
flabel metal2 17352 8665 17352 8665 0 FreeSans 240 0 0 0 vtrip_decoded_avdd[1]
port 18 nsew
flabel metal2 17886 8665 17886 8665 0 FreeSans 240 0 0 0 vtrip_decoded_avdd[2]
port 17 nsew
flabel metal2 18420 8665 18420 8665 0 FreeSans 240 0 0 0 vtrip_decoded_avdd[3]
port 16 nsew
flabel metal2 18954 8665 18954 8665 0 FreeSans 240 0 0 0 vtrip_decoded_avdd[4]
port 15 nsew
flabel metal2 19488 8665 19488 8665 0 FreeSans 240 0 0 0 vtrip_decoded_avdd[5]
port 14 nsew
flabel metal2 20022 8665 20022 8665 0 FreeSans 240 0 0 0 vtrip_decoded_avdd[6]
port 13 nsew
flabel metal2 20556 8665 20556 8665 0 FreeSans 240 0 0 0 vtrip_decoded_avdd[7]
port 12 nsew
flabel metal2 17037 8531 17037 8531 0 FreeSans 160 0 0 0 vtrip_decoded_b_avdd[0]
flabel metal2 17571 8531 17571 8531 0 FreeSans 160 0 0 0 vtrip_decoded_b_avdd[1]
flabel metal2 18105 8531 18105 8531 0 FreeSans 160 0 0 0 vtrip_decoded_b_avdd[2]
flabel metal2 18639 8531 18639 8531 0 FreeSans 160 0 0 0 vtrip_decoded_b_avdd[3]
flabel metal2 19173 8531 19173 8531 0 FreeSans 160 0 0 0 vtrip_decoded_b_avdd[4]
flabel metal2 19707 8531 19707 8531 0 FreeSans 160 0 0 0 vtrip_decoded_b_avdd[5]
flabel metal2 20241 8531 20241 8531 0 FreeSans 160 0 0 0 vtrip_decoded_b_avdd[6]
flabel metal2 20775 8531 20775 8531 0 FreeSans 160 0 0 0 vtrip_decoded_b_avdd[7]
flabel metal3 s 20983 7113 20983 7113 0 FreeSans 1200 0 0 0 vout_vunder
port 20 nsew
flabel metal3 s 16711 7113 16711 7113 0 FreeSans 1200 0 0 0 vout_brout
port 2 nsew
flabel metal2 s 8930 5097 8930 5097 0 FreeSans 800 0 0 0 vtop
<< end >>
